magic
tech gf180mcuD
magscale 1 10
timestamp 1764342644
<< nwell >>
rect 15280 46078 15875 46628
<< nmos >>
rect 15581 45872 15637 45992
<< pmos >>
rect 15581 46164 15637 46404
<< ndiff >>
rect 15492 45979 15581 45992
rect 15492 45887 15506 45979
rect 15552 45887 15581 45979
rect 15492 45872 15581 45887
rect 15637 45978 15725 45992
rect 15637 45886 15666 45978
rect 15712 45886 15725 45978
rect 15637 45872 15725 45886
<< pdiff >>
rect 15493 46390 15581 46404
rect 15493 46177 15506 46390
rect 15552 46177 15581 46390
rect 15493 46164 15581 46177
rect 15637 46390 15725 46404
rect 15637 46177 15666 46390
rect 15712 46177 15725 46390
rect 15637 46164 15725 46177
<< ndiffc >>
rect 15506 45887 15552 45979
rect 15666 45886 15712 45978
<< pdiffc >>
rect 15506 46177 15552 46390
rect 15666 46177 15712 46390
<< psubdiff >>
rect 15366 45791 15789 45806
rect 15366 45745 15379 45791
rect 15425 45745 15730 45791
rect 15776 45745 15789 45791
rect 15366 45730 15789 45745
<< nsubdiff >>
rect 15366 46531 15789 46546
rect 15366 46485 15379 46531
rect 15425 46485 15730 46531
rect 15776 46485 15789 46531
rect 15366 46470 15789 46485
<< psubdiffcont >>
rect 15379 45745 15425 45791
rect 15730 45745 15776 45791
<< nsubdiffcont >>
rect 15379 46485 15425 46531
rect 15730 46485 15776 46531
<< polysilicon >>
rect 15581 46404 15637 46450
rect 15396 46241 15468 46254
rect 15396 46121 15409 46241
rect 15455 46144 15468 46241
rect 15581 46144 15637 46164
rect 15455 46121 15637 46144
rect 15396 46108 15637 46121
rect 15397 46045 15637 46058
rect 15397 45925 15410 46045
rect 15456 46022 15637 46045
rect 15456 45925 15469 46022
rect 15581 45992 15637 46022
rect 15397 45912 15469 45925
rect 15581 45828 15637 45872
<< polycontact >>
rect 15409 46121 15455 46241
rect 15410 45925 15456 46045
<< metal1 >>
rect 15366 46531 15789 46542
rect 15366 46485 15379 46531
rect 15425 46485 15730 46531
rect 15776 46485 15789 46531
rect 15366 46467 15789 46485
rect 15506 46390 15552 46401
rect 15409 46241 15455 46252
rect 15409 46110 15455 46121
rect 15410 46045 15456 46056
rect 15410 45914 15456 45925
rect 15506 45979 15552 46177
rect 15506 45876 15552 45887
rect 15666 46390 15712 46401
rect 15666 45978 15712 46177
rect 15666 45875 15712 45886
rect 15366 45791 15789 45810
rect 15366 45745 15379 45791
rect 15425 45745 15730 45791
rect 15776 45745 15789 45791
rect 15366 45734 15789 45745
<< end >>
