magic
tech gf180mcuD
magscale 1 10
timestamp 1764775243
<< metal2 >>
rect -400 12949 13200 13065
rect -400 12893 -254 12949
rect -198 12893 -130 12949
rect -74 12893 -6 12949
rect 50 12893 118 12949
rect 174 12893 242 12949
rect 298 12893 366 12949
rect 422 12893 490 12949
rect 546 12893 614 12949
rect 670 12893 738 12949
rect 794 12893 862 12949
rect 918 12893 986 12949
rect 1042 12893 1110 12949
rect 1166 12893 1234 12949
rect 1290 12893 1358 12949
rect 1414 12893 1482 12949
rect 1538 12893 1606 12949
rect 1662 12893 1730 12949
rect 1786 12893 1854 12949
rect 1910 12893 1978 12949
rect 2034 12893 2102 12949
rect 2158 12893 2226 12949
rect 2282 12893 2350 12949
rect 2406 12893 2474 12949
rect 2530 12893 2598 12949
rect 2654 12893 2722 12949
rect 2778 12893 2846 12949
rect 2902 12893 2970 12949
rect 3026 12893 3094 12949
rect 3150 12893 3218 12949
rect 3274 12893 3342 12949
rect 3398 12893 3466 12949
rect 3522 12893 3590 12949
rect 3646 12893 3714 12949
rect 3770 12893 3838 12949
rect 3894 12893 3962 12949
rect 4018 12893 4086 12949
rect 4142 12893 4210 12949
rect 4266 12893 4334 12949
rect 4390 12893 4458 12949
rect 4514 12893 4582 12949
rect 4638 12893 4706 12949
rect 4762 12893 4830 12949
rect 4886 12893 4954 12949
rect 5010 12893 5078 12949
rect 5134 12893 5202 12949
rect 5258 12893 5326 12949
rect 5382 12893 5450 12949
rect 5506 12893 5574 12949
rect 5630 12893 5698 12949
rect 5754 12893 5822 12949
rect 5878 12893 5946 12949
rect 6002 12893 6070 12949
rect 6126 12893 6194 12949
rect 6250 12893 6318 12949
rect 6374 12893 6442 12949
rect 6498 12893 6566 12949
rect 6622 12893 6690 12949
rect 6746 12893 6814 12949
rect 6870 12893 6938 12949
rect 6994 12893 7062 12949
rect 7118 12893 7186 12949
rect 7242 12893 7310 12949
rect 7366 12893 7434 12949
rect 7490 12893 7558 12949
rect 7614 12893 7682 12949
rect 7738 12893 7806 12949
rect 7862 12893 7930 12949
rect 7986 12893 8054 12949
rect 8110 12893 8178 12949
rect 8234 12893 8302 12949
rect 8358 12893 8426 12949
rect 8482 12893 8550 12949
rect 8606 12893 8674 12949
rect 8730 12893 8798 12949
rect 8854 12893 8922 12949
rect 8978 12893 9046 12949
rect 9102 12893 9170 12949
rect 9226 12893 9294 12949
rect 9350 12893 9418 12949
rect 9474 12893 9542 12949
rect 9598 12893 9666 12949
rect 9722 12893 9790 12949
rect 9846 12893 9914 12949
rect 9970 12893 10038 12949
rect 10094 12893 10162 12949
rect 10218 12893 10286 12949
rect 10342 12893 10410 12949
rect 10466 12893 10534 12949
rect 10590 12893 10658 12949
rect 10714 12893 10782 12949
rect 10838 12893 10906 12949
rect 10962 12893 11030 12949
rect 11086 12893 11154 12949
rect 11210 12893 11278 12949
rect 11334 12893 11402 12949
rect 11458 12893 11526 12949
rect 11582 12893 11650 12949
rect 11706 12893 11774 12949
rect 11830 12893 11898 12949
rect 11954 12893 12022 12949
rect 12078 12893 12146 12949
rect 12202 12893 12270 12949
rect 12326 12893 12394 12949
rect 12450 12893 12518 12949
rect 12574 12893 12642 12949
rect 12698 12893 12766 12949
rect 12822 12893 12890 12949
rect 12946 12893 13014 12949
rect 13070 12893 13200 12949
rect -400 12825 13200 12893
rect -400 12769 -254 12825
rect -198 12769 -130 12825
rect -74 12769 -6 12825
rect 50 12769 118 12825
rect 174 12769 242 12825
rect 298 12769 366 12825
rect 422 12769 490 12825
rect 546 12769 614 12825
rect 670 12769 738 12825
rect 794 12769 862 12825
rect 918 12769 986 12825
rect 1042 12769 1110 12825
rect 1166 12769 1234 12825
rect 1290 12769 1358 12825
rect 1414 12769 1482 12825
rect 1538 12769 1606 12825
rect 1662 12769 1730 12825
rect 1786 12769 1854 12825
rect 1910 12769 1978 12825
rect 2034 12769 2102 12825
rect 2158 12769 2226 12825
rect 2282 12769 2350 12825
rect 2406 12769 2474 12825
rect 2530 12769 2598 12825
rect 2654 12769 2722 12825
rect 2778 12769 2846 12825
rect 2902 12769 2970 12825
rect 3026 12769 3094 12825
rect 3150 12769 3218 12825
rect 3274 12769 3342 12825
rect 3398 12769 3466 12825
rect 3522 12769 3590 12825
rect 3646 12769 3714 12825
rect 3770 12769 3838 12825
rect 3894 12769 3962 12825
rect 4018 12769 4086 12825
rect 4142 12769 4210 12825
rect 4266 12769 4334 12825
rect 4390 12769 4458 12825
rect 4514 12769 4582 12825
rect 4638 12769 4706 12825
rect 4762 12769 4830 12825
rect 4886 12769 4954 12825
rect 5010 12769 5078 12825
rect 5134 12769 5202 12825
rect 5258 12769 5326 12825
rect 5382 12769 5450 12825
rect 5506 12769 5574 12825
rect 5630 12769 5698 12825
rect 5754 12769 5822 12825
rect 5878 12769 5946 12825
rect 6002 12769 6070 12825
rect 6126 12769 6194 12825
rect 6250 12769 6318 12825
rect 6374 12769 6442 12825
rect 6498 12769 6566 12825
rect 6622 12769 6690 12825
rect 6746 12769 6814 12825
rect 6870 12769 6938 12825
rect 6994 12769 7062 12825
rect 7118 12769 7186 12825
rect 7242 12769 7310 12825
rect 7366 12769 7434 12825
rect 7490 12769 7558 12825
rect 7614 12769 7682 12825
rect 7738 12769 7806 12825
rect 7862 12769 7930 12825
rect 7986 12769 8054 12825
rect 8110 12769 8178 12825
rect 8234 12769 8302 12825
rect 8358 12769 8426 12825
rect 8482 12769 8550 12825
rect 8606 12769 8674 12825
rect 8730 12769 8798 12825
rect 8854 12769 8922 12825
rect 8978 12769 9046 12825
rect 9102 12769 9170 12825
rect 9226 12769 9294 12825
rect 9350 12769 9418 12825
rect 9474 12769 9542 12825
rect 9598 12769 9666 12825
rect 9722 12769 9790 12825
rect 9846 12769 9914 12825
rect 9970 12769 10038 12825
rect 10094 12769 10162 12825
rect 10218 12769 10286 12825
rect 10342 12769 10410 12825
rect 10466 12769 10534 12825
rect 10590 12769 10658 12825
rect 10714 12769 10782 12825
rect 10838 12769 10906 12825
rect 10962 12769 11030 12825
rect 11086 12769 11154 12825
rect 11210 12769 11278 12825
rect 11334 12769 11402 12825
rect 11458 12769 11526 12825
rect 11582 12769 11650 12825
rect 11706 12769 11774 12825
rect 11830 12769 11898 12825
rect 11954 12769 12022 12825
rect 12078 12769 12146 12825
rect 12202 12769 12270 12825
rect 12326 12769 12394 12825
rect 12450 12769 12518 12825
rect 12574 12769 12642 12825
rect 12698 12769 12766 12825
rect 12822 12769 12890 12825
rect 12946 12769 13014 12825
rect 13070 12769 13200 12825
rect -400 12701 13200 12769
rect -400 12645 -254 12701
rect -198 12645 -130 12701
rect -74 12645 -6 12701
rect 50 12645 118 12701
rect 174 12645 242 12701
rect 298 12645 366 12701
rect 422 12645 490 12701
rect 546 12645 614 12701
rect 670 12645 738 12701
rect 794 12645 862 12701
rect 918 12645 986 12701
rect 1042 12645 1110 12701
rect 1166 12645 1234 12701
rect 1290 12645 1358 12701
rect 1414 12645 1482 12701
rect 1538 12645 1606 12701
rect 1662 12645 1730 12701
rect 1786 12645 1854 12701
rect 1910 12645 1978 12701
rect 2034 12645 2102 12701
rect 2158 12645 2226 12701
rect 2282 12645 2350 12701
rect 2406 12645 2474 12701
rect 2530 12645 2598 12701
rect 2654 12645 2722 12701
rect 2778 12645 2846 12701
rect 2902 12645 2970 12701
rect 3026 12645 3094 12701
rect 3150 12645 3218 12701
rect 3274 12645 3342 12701
rect 3398 12645 3466 12701
rect 3522 12645 3590 12701
rect 3646 12645 3714 12701
rect 3770 12645 3838 12701
rect 3894 12645 3962 12701
rect 4018 12645 4086 12701
rect 4142 12645 4210 12701
rect 4266 12645 4334 12701
rect 4390 12645 4458 12701
rect 4514 12645 4582 12701
rect 4638 12645 4706 12701
rect 4762 12645 4830 12701
rect 4886 12645 4954 12701
rect 5010 12645 5078 12701
rect 5134 12645 5202 12701
rect 5258 12645 5326 12701
rect 5382 12645 5450 12701
rect 5506 12645 5574 12701
rect 5630 12645 5698 12701
rect 5754 12645 5822 12701
rect 5878 12645 5946 12701
rect 6002 12645 6070 12701
rect 6126 12645 6194 12701
rect 6250 12645 6318 12701
rect 6374 12645 6442 12701
rect 6498 12645 6566 12701
rect 6622 12645 6690 12701
rect 6746 12645 6814 12701
rect 6870 12645 6938 12701
rect 6994 12645 7062 12701
rect 7118 12645 7186 12701
rect 7242 12645 7310 12701
rect 7366 12645 7434 12701
rect 7490 12645 7558 12701
rect 7614 12645 7682 12701
rect 7738 12645 7806 12701
rect 7862 12645 7930 12701
rect 7986 12645 8054 12701
rect 8110 12645 8178 12701
rect 8234 12645 8302 12701
rect 8358 12645 8426 12701
rect 8482 12645 8550 12701
rect 8606 12645 8674 12701
rect 8730 12645 8798 12701
rect 8854 12645 8922 12701
rect 8978 12645 9046 12701
rect 9102 12645 9170 12701
rect 9226 12645 9294 12701
rect 9350 12645 9418 12701
rect 9474 12645 9542 12701
rect 9598 12645 9666 12701
rect 9722 12645 9790 12701
rect 9846 12645 9914 12701
rect 9970 12645 10038 12701
rect 10094 12645 10162 12701
rect 10218 12645 10286 12701
rect 10342 12645 10410 12701
rect 10466 12645 10534 12701
rect 10590 12645 10658 12701
rect 10714 12645 10782 12701
rect 10838 12645 10906 12701
rect 10962 12645 11030 12701
rect 11086 12645 11154 12701
rect 11210 12645 11278 12701
rect 11334 12645 11402 12701
rect 11458 12645 11526 12701
rect 11582 12645 11650 12701
rect 11706 12645 11774 12701
rect 11830 12645 11898 12701
rect 11954 12645 12022 12701
rect 12078 12645 12146 12701
rect 12202 12645 12270 12701
rect 12326 12645 12394 12701
rect 12450 12645 12518 12701
rect 12574 12645 12642 12701
rect 12698 12645 12766 12701
rect 12822 12645 12890 12701
rect 12946 12645 13014 12701
rect 13070 12645 13200 12701
rect -400 12577 13200 12645
rect -400 12521 -254 12577
rect -198 12521 -130 12577
rect -74 12521 -6 12577
rect 50 12521 118 12577
rect 174 12521 242 12577
rect 298 12521 366 12577
rect 422 12521 490 12577
rect 546 12521 614 12577
rect 670 12521 738 12577
rect 794 12521 862 12577
rect 918 12521 986 12577
rect 1042 12521 1110 12577
rect 1166 12521 1234 12577
rect 1290 12521 1358 12577
rect 1414 12521 1482 12577
rect 1538 12521 1606 12577
rect 1662 12521 1730 12577
rect 1786 12521 1854 12577
rect 1910 12521 1978 12577
rect 2034 12521 2102 12577
rect 2158 12521 2226 12577
rect 2282 12521 2350 12577
rect 2406 12521 2474 12577
rect 2530 12521 2598 12577
rect 2654 12521 2722 12577
rect 2778 12521 2846 12577
rect 2902 12521 2970 12577
rect 3026 12521 3094 12577
rect 3150 12521 3218 12577
rect 3274 12521 3342 12577
rect 3398 12521 3466 12577
rect 3522 12521 3590 12577
rect 3646 12521 3714 12577
rect 3770 12521 3838 12577
rect 3894 12521 3962 12577
rect 4018 12521 4086 12577
rect 4142 12521 4210 12577
rect 4266 12521 4334 12577
rect 4390 12521 4458 12577
rect 4514 12521 4582 12577
rect 4638 12521 4706 12577
rect 4762 12521 4830 12577
rect 4886 12521 4954 12577
rect 5010 12521 5078 12577
rect 5134 12521 5202 12577
rect 5258 12521 5326 12577
rect 5382 12521 5450 12577
rect 5506 12521 5574 12577
rect 5630 12521 5698 12577
rect 5754 12521 5822 12577
rect 5878 12521 5946 12577
rect 6002 12521 6070 12577
rect 6126 12521 6194 12577
rect 6250 12521 6318 12577
rect 6374 12521 6442 12577
rect 6498 12521 6566 12577
rect 6622 12521 6690 12577
rect 6746 12521 6814 12577
rect 6870 12521 6938 12577
rect 6994 12521 7062 12577
rect 7118 12521 7186 12577
rect 7242 12521 7310 12577
rect 7366 12521 7434 12577
rect 7490 12521 7558 12577
rect 7614 12521 7682 12577
rect 7738 12521 7806 12577
rect 7862 12521 7930 12577
rect 7986 12521 8054 12577
rect 8110 12521 8178 12577
rect 8234 12521 8302 12577
rect 8358 12521 8426 12577
rect 8482 12521 8550 12577
rect 8606 12521 8674 12577
rect 8730 12521 8798 12577
rect 8854 12521 8922 12577
rect 8978 12521 9046 12577
rect 9102 12521 9170 12577
rect 9226 12521 9294 12577
rect 9350 12521 9418 12577
rect 9474 12521 9542 12577
rect 9598 12521 9666 12577
rect 9722 12521 9790 12577
rect 9846 12521 9914 12577
rect 9970 12521 10038 12577
rect 10094 12521 10162 12577
rect 10218 12521 10286 12577
rect 10342 12521 10410 12577
rect 10466 12521 10534 12577
rect 10590 12521 10658 12577
rect 10714 12521 10782 12577
rect 10838 12521 10906 12577
rect 10962 12521 11030 12577
rect 11086 12521 11154 12577
rect 11210 12521 11278 12577
rect 11334 12521 11402 12577
rect 11458 12521 11526 12577
rect 11582 12521 11650 12577
rect 11706 12521 11774 12577
rect 11830 12521 11898 12577
rect 11954 12521 12022 12577
rect 12078 12521 12146 12577
rect 12202 12521 12270 12577
rect 12326 12521 12394 12577
rect 12450 12521 12518 12577
rect 12574 12521 12642 12577
rect 12698 12521 12766 12577
rect 12822 12521 12890 12577
rect 12946 12521 13014 12577
rect 13070 12521 13200 12577
rect -400 12400 13200 12521
rect -400 12358 400 12400
rect -400 12302 -286 12358
rect -230 12302 -162 12358
rect -106 12302 -38 12358
rect 18 12302 86 12358
rect 142 12302 210 12358
rect 266 12302 400 12358
rect -400 12234 400 12302
rect -400 12178 -286 12234
rect -230 12178 -162 12234
rect -106 12178 -38 12234
rect 18 12178 86 12234
rect 142 12178 210 12234
rect 266 12178 400 12234
rect -400 12110 400 12178
rect -400 12054 -286 12110
rect -230 12054 -162 12110
rect -106 12054 -38 12110
rect 18 12054 86 12110
rect 142 12054 210 12110
rect 266 12054 400 12110
rect -400 11986 400 12054
rect -400 11930 -286 11986
rect -230 11930 -162 11986
rect -106 11930 -38 11986
rect 18 11930 86 11986
rect 142 11930 210 11986
rect 266 11930 400 11986
rect -400 11862 400 11930
rect -400 11806 -286 11862
rect -230 11806 -162 11862
rect -106 11806 -38 11862
rect 18 11806 86 11862
rect 142 11806 210 11862
rect 266 11806 400 11862
rect -400 11738 400 11806
rect -400 11682 -286 11738
rect -230 11682 -162 11738
rect -106 11682 -38 11738
rect 18 11682 86 11738
rect 142 11682 210 11738
rect 266 11682 400 11738
rect -400 11614 400 11682
rect -400 11558 -286 11614
rect -230 11558 -162 11614
rect -106 11558 -38 11614
rect 18 11558 86 11614
rect 142 11558 210 11614
rect 266 11558 400 11614
rect -400 11490 400 11558
rect -400 11434 -286 11490
rect -230 11434 -162 11490
rect -106 11434 -38 11490
rect 18 11434 86 11490
rect 142 11434 210 11490
rect 266 11434 400 11490
rect -400 11366 400 11434
rect -400 11310 -286 11366
rect -230 11310 -162 11366
rect -106 11310 -38 11366
rect 18 11310 86 11366
rect 142 11310 210 11366
rect 266 11310 400 11366
rect -400 11242 400 11310
rect -400 11186 -286 11242
rect -230 11186 -162 11242
rect -106 11186 -38 11242
rect 18 11186 86 11242
rect 142 11186 210 11242
rect 266 11186 400 11242
rect -400 11118 400 11186
rect -400 11062 -286 11118
rect -230 11062 -162 11118
rect -106 11062 -38 11118
rect 18 11062 86 11118
rect 142 11062 210 11118
rect 266 11062 400 11118
rect -400 10994 400 11062
rect -400 10938 -286 10994
rect -230 10938 -162 10994
rect -106 10938 -38 10994
rect 18 10938 86 10994
rect 142 10938 210 10994
rect 266 10938 400 10994
rect -400 10870 400 10938
rect -400 10814 -286 10870
rect -230 10814 -162 10870
rect -106 10814 -38 10870
rect 18 10814 86 10870
rect 142 10814 210 10870
rect 266 10814 400 10870
rect -400 10746 400 10814
rect -400 10690 -286 10746
rect -230 10690 -162 10746
rect -106 10690 -38 10746
rect 18 10690 86 10746
rect 142 10690 210 10746
rect 266 10690 400 10746
rect -400 10622 400 10690
rect -400 10566 -286 10622
rect -230 10566 -162 10622
rect -106 10566 -38 10622
rect 18 10566 86 10622
rect 142 10566 210 10622
rect 266 10566 400 10622
rect -400 10498 400 10566
rect -400 10442 -286 10498
rect -230 10442 -162 10498
rect -106 10442 -38 10498
rect 18 10442 86 10498
rect 142 10442 210 10498
rect 266 10442 400 10498
rect -400 10374 400 10442
rect -400 10318 -286 10374
rect -230 10318 -162 10374
rect -106 10318 -38 10374
rect 18 10318 86 10374
rect 142 10318 210 10374
rect 266 10318 400 10374
rect -400 10250 400 10318
rect -400 10194 -286 10250
rect -230 10194 -162 10250
rect -106 10194 -38 10250
rect 18 10194 86 10250
rect 142 10194 210 10250
rect 266 10194 400 10250
rect -400 10126 400 10194
rect -400 10070 -286 10126
rect -230 10070 -162 10126
rect -106 10070 -38 10126
rect 18 10070 86 10126
rect 142 10070 210 10126
rect 266 10070 400 10126
rect -400 10002 400 10070
rect -400 9946 -286 10002
rect -230 9946 -162 10002
rect -106 9946 -38 10002
rect 18 9946 86 10002
rect 142 9946 210 10002
rect 266 9946 400 10002
rect -400 9878 400 9946
rect -400 9822 -286 9878
rect -230 9822 -162 9878
rect -106 9822 -38 9878
rect 18 9822 86 9878
rect 142 9822 210 9878
rect 266 9822 400 9878
rect -400 9754 400 9822
rect -400 9698 -286 9754
rect -230 9698 -162 9754
rect -106 9698 -38 9754
rect 18 9698 86 9754
rect 142 9698 210 9754
rect 266 9698 400 9754
rect -400 9630 400 9698
rect -400 9574 -286 9630
rect -230 9574 -162 9630
rect -106 9574 -38 9630
rect 18 9574 86 9630
rect 142 9574 210 9630
rect 266 9574 400 9630
rect -400 9506 400 9574
rect -400 9450 -286 9506
rect -230 9450 -162 9506
rect -106 9450 -38 9506
rect 18 9450 86 9506
rect 142 9450 210 9506
rect 266 9450 400 9506
rect -400 9382 400 9450
rect -400 9326 -286 9382
rect -230 9326 -162 9382
rect -106 9326 -38 9382
rect 18 9326 86 9382
rect 142 9326 210 9382
rect 266 9326 400 9382
rect -400 9258 400 9326
rect -400 9202 -286 9258
rect -230 9202 -162 9258
rect -106 9202 -38 9258
rect 18 9202 86 9258
rect 142 9202 210 9258
rect 266 9202 400 9258
rect -400 9134 400 9202
rect -400 9078 -286 9134
rect -230 9078 -162 9134
rect -106 9078 -38 9134
rect 18 9078 86 9134
rect 142 9078 210 9134
rect 266 9078 400 9134
rect -400 9010 400 9078
rect -400 8954 -286 9010
rect -230 8954 -162 9010
rect -106 8954 -38 9010
rect 18 8954 86 9010
rect 142 8954 210 9010
rect 266 8954 400 9010
rect -400 8886 400 8954
rect -400 8830 -286 8886
rect -230 8830 -162 8886
rect -106 8830 -38 8886
rect 18 8830 86 8886
rect 142 8830 210 8886
rect 266 8830 400 8886
rect -400 8762 400 8830
rect -400 8706 -286 8762
rect -230 8706 -162 8762
rect -106 8706 -38 8762
rect 18 8706 86 8762
rect 142 8706 210 8762
rect 266 8706 400 8762
rect -400 8638 400 8706
rect -400 8582 -286 8638
rect -230 8582 -162 8638
rect -106 8582 -38 8638
rect 18 8582 86 8638
rect 142 8582 210 8638
rect 266 8582 400 8638
rect -400 8514 400 8582
rect -400 8458 -286 8514
rect -230 8458 -162 8514
rect -106 8458 -38 8514
rect 18 8458 86 8514
rect 142 8458 210 8514
rect 266 8458 400 8514
rect -400 8390 400 8458
rect -400 8334 -286 8390
rect -230 8334 -162 8390
rect -106 8334 -38 8390
rect 18 8334 86 8390
rect 142 8334 210 8390
rect 266 8334 400 8390
rect -400 8266 400 8334
rect -400 8210 -286 8266
rect -230 8210 -162 8266
rect -106 8210 -38 8266
rect 18 8210 86 8266
rect 142 8210 210 8266
rect 266 8210 400 8266
rect -400 8142 400 8210
rect -400 8086 -286 8142
rect -230 8086 -162 8142
rect -106 8086 -38 8142
rect 18 8086 86 8142
rect 142 8086 210 8142
rect 266 8086 400 8142
rect -400 8018 400 8086
rect -400 7962 -286 8018
rect -230 7962 -162 8018
rect -106 7962 -38 8018
rect 18 7962 86 8018
rect 142 7962 210 8018
rect 266 7962 400 8018
rect -400 7894 400 7962
rect -400 7838 -286 7894
rect -230 7838 -162 7894
rect -106 7838 -38 7894
rect 18 7838 86 7894
rect 142 7838 210 7894
rect 266 7838 400 7894
rect -400 7770 400 7838
rect -400 7714 -286 7770
rect -230 7714 -162 7770
rect -106 7714 -38 7770
rect 18 7714 86 7770
rect 142 7714 210 7770
rect 266 7714 400 7770
rect -400 7646 400 7714
rect -400 7590 -286 7646
rect -230 7590 -162 7646
rect -106 7590 -38 7646
rect 18 7590 86 7646
rect 142 7590 210 7646
rect 266 7590 400 7646
rect -400 7522 400 7590
rect -400 7466 -286 7522
rect -230 7466 -162 7522
rect -106 7466 -38 7522
rect 18 7466 86 7522
rect 142 7466 210 7522
rect 266 7466 400 7522
rect -400 7398 400 7466
rect -400 7342 -286 7398
rect -230 7342 -162 7398
rect -106 7342 -38 7398
rect 18 7342 86 7398
rect 142 7342 210 7398
rect 266 7342 400 7398
rect -400 7274 400 7342
rect -400 7218 -286 7274
rect -230 7218 -162 7274
rect -106 7218 -38 7274
rect 18 7218 86 7274
rect 142 7218 210 7274
rect 266 7218 400 7274
rect -400 7150 400 7218
rect -400 7094 -286 7150
rect -230 7094 -162 7150
rect -106 7094 -38 7150
rect 18 7094 86 7150
rect 142 7094 210 7150
rect 266 7094 400 7150
rect -400 7026 400 7094
rect -400 6970 -286 7026
rect -230 6970 -162 7026
rect -106 6970 -38 7026
rect 18 6970 86 7026
rect 142 6970 210 7026
rect 266 6970 400 7026
rect -400 6902 400 6970
rect -400 6846 -286 6902
rect -230 6846 -162 6902
rect -106 6846 -38 6902
rect 18 6846 86 6902
rect 142 6846 210 6902
rect 266 6846 400 6902
rect -400 6778 400 6846
rect -400 6722 -286 6778
rect -230 6722 -162 6778
rect -106 6722 -38 6778
rect 18 6722 86 6778
rect 142 6722 210 6778
rect 266 6722 400 6778
rect -400 6654 400 6722
rect -400 6598 -286 6654
rect -230 6598 -162 6654
rect -106 6598 -38 6654
rect 18 6598 86 6654
rect 142 6598 210 6654
rect 266 6598 400 6654
rect -400 6530 400 6598
rect -400 6474 -286 6530
rect -230 6474 -162 6530
rect -106 6474 -38 6530
rect 18 6474 86 6530
rect 142 6474 210 6530
rect 266 6474 400 6530
rect -400 6406 400 6474
rect -400 6350 -286 6406
rect -230 6350 -162 6406
rect -106 6350 -38 6406
rect 18 6350 86 6406
rect 142 6350 210 6406
rect 266 6350 400 6406
rect -400 6282 400 6350
rect -400 6226 -286 6282
rect -230 6226 -162 6282
rect -106 6226 -38 6282
rect 18 6226 86 6282
rect 142 6226 210 6282
rect 266 6226 400 6282
rect -400 6158 400 6226
rect -400 6102 -286 6158
rect -230 6102 -162 6158
rect -106 6102 -38 6158
rect 18 6102 86 6158
rect 142 6102 210 6158
rect 266 6102 400 6158
rect -400 6034 400 6102
rect -400 5978 -286 6034
rect -230 5978 -162 6034
rect -106 5978 -38 6034
rect 18 5978 86 6034
rect 142 5978 210 6034
rect 266 5978 400 6034
rect -400 5910 400 5978
rect -400 5854 -286 5910
rect -230 5854 -162 5910
rect -106 5854 -38 5910
rect 18 5854 86 5910
rect 142 5854 210 5910
rect 266 5854 400 5910
rect -400 5786 400 5854
rect -400 5730 -286 5786
rect -230 5730 -162 5786
rect -106 5730 -38 5786
rect 18 5730 86 5786
rect 142 5730 210 5786
rect 266 5730 400 5786
rect -400 5662 400 5730
rect -400 5606 -286 5662
rect -230 5606 -162 5662
rect -106 5606 -38 5662
rect 18 5606 86 5662
rect 142 5606 210 5662
rect 266 5606 400 5662
rect -400 5538 400 5606
rect -400 5482 -286 5538
rect -230 5482 -162 5538
rect -106 5482 -38 5538
rect 18 5482 86 5538
rect 142 5482 210 5538
rect 266 5482 400 5538
rect -400 5414 400 5482
rect -400 5358 -286 5414
rect -230 5358 -162 5414
rect -106 5358 -38 5414
rect 18 5358 86 5414
rect 142 5358 210 5414
rect 266 5358 400 5414
rect -400 5290 400 5358
rect -400 5234 -286 5290
rect -230 5234 -162 5290
rect -106 5234 -38 5290
rect 18 5234 86 5290
rect 142 5234 210 5290
rect 266 5234 400 5290
rect -400 5166 400 5234
rect -400 5110 -286 5166
rect -230 5110 -162 5166
rect -106 5110 -38 5166
rect 18 5110 86 5166
rect 142 5110 210 5166
rect 266 5110 400 5166
rect -400 5042 400 5110
rect -400 4986 -286 5042
rect -230 4986 -162 5042
rect -106 4986 -38 5042
rect 18 4986 86 5042
rect 142 4986 210 5042
rect 266 4986 400 5042
rect -400 4918 400 4986
rect -400 4862 -286 4918
rect -230 4862 -162 4918
rect -106 4862 -38 4918
rect 18 4862 86 4918
rect 142 4862 210 4918
rect 266 4862 400 4918
rect -400 4794 400 4862
rect -400 4738 -286 4794
rect -230 4738 -162 4794
rect -106 4738 -38 4794
rect 18 4738 86 4794
rect 142 4738 210 4794
rect 266 4738 400 4794
rect -400 4670 400 4738
rect -400 4614 -286 4670
rect -230 4614 -162 4670
rect -106 4614 -38 4670
rect 18 4614 86 4670
rect 142 4614 210 4670
rect 266 4614 400 4670
rect -400 4546 400 4614
rect -400 4490 -286 4546
rect -230 4490 -162 4546
rect -106 4490 -38 4546
rect 18 4490 86 4546
rect 142 4490 210 4546
rect 266 4490 400 4546
rect -400 4422 400 4490
rect -400 4366 -286 4422
rect -230 4366 -162 4422
rect -106 4366 -38 4422
rect 18 4366 86 4422
rect 142 4366 210 4422
rect 266 4366 400 4422
rect -400 4298 400 4366
rect -400 4242 -286 4298
rect -230 4242 -162 4298
rect -106 4242 -38 4298
rect 18 4242 86 4298
rect 142 4242 210 4298
rect 266 4242 400 4298
rect -400 4174 400 4242
rect -400 4118 -286 4174
rect -230 4118 -162 4174
rect -106 4118 -38 4174
rect 18 4118 86 4174
rect 142 4118 210 4174
rect 266 4118 400 4174
rect -400 4050 400 4118
rect -400 3994 -286 4050
rect -230 3994 -162 4050
rect -106 3994 -38 4050
rect 18 3994 86 4050
rect 142 3994 210 4050
rect 266 3994 400 4050
rect -400 3926 400 3994
rect -400 3870 -286 3926
rect -230 3870 -162 3926
rect -106 3870 -38 3926
rect 18 3870 86 3926
rect 142 3870 210 3926
rect 266 3870 400 3926
rect -400 3802 400 3870
rect -400 3746 -286 3802
rect -230 3746 -162 3802
rect -106 3746 -38 3802
rect 18 3746 86 3802
rect 142 3746 210 3802
rect 266 3746 400 3802
rect -400 3678 400 3746
rect -400 3622 -286 3678
rect -230 3622 -162 3678
rect -106 3622 -38 3678
rect 18 3622 86 3678
rect 142 3622 210 3678
rect 266 3622 400 3678
rect -400 3554 400 3622
rect -400 3498 -286 3554
rect -230 3498 -162 3554
rect -106 3498 -38 3554
rect 18 3498 86 3554
rect 142 3498 210 3554
rect 266 3498 400 3554
rect -400 3430 400 3498
rect -400 3374 -286 3430
rect -230 3374 -162 3430
rect -106 3374 -38 3430
rect 18 3374 86 3430
rect 142 3374 210 3430
rect 266 3374 400 3430
rect -400 3306 400 3374
rect -400 3250 -286 3306
rect -230 3250 -162 3306
rect -106 3250 -38 3306
rect 18 3250 86 3306
rect 142 3250 210 3306
rect 266 3250 400 3306
rect -400 3182 400 3250
rect -400 3126 -286 3182
rect -230 3126 -162 3182
rect -106 3126 -38 3182
rect 18 3126 86 3182
rect 142 3126 210 3182
rect 266 3126 400 3182
rect -400 3058 400 3126
rect -400 3002 -286 3058
rect -230 3002 -162 3058
rect -106 3002 -38 3058
rect 18 3002 86 3058
rect 142 3002 210 3058
rect 266 3002 400 3058
rect -400 2934 400 3002
rect -400 2878 -286 2934
rect -230 2878 -162 2934
rect -106 2878 -38 2934
rect 18 2878 86 2934
rect 142 2878 210 2934
rect 266 2878 400 2934
rect -400 2810 400 2878
rect -400 2754 -286 2810
rect -230 2754 -162 2810
rect -106 2754 -38 2810
rect 18 2754 86 2810
rect 142 2754 210 2810
rect 266 2754 400 2810
rect -400 2686 400 2754
rect -400 2630 -286 2686
rect -230 2630 -162 2686
rect -106 2630 -38 2686
rect 18 2630 86 2686
rect 142 2630 210 2686
rect 266 2630 400 2686
rect -400 2562 400 2630
rect -400 2506 -286 2562
rect -230 2506 -162 2562
rect -106 2506 -38 2562
rect 18 2506 86 2562
rect 142 2506 210 2562
rect 266 2506 400 2562
rect -400 2438 400 2506
rect -400 2382 -286 2438
rect -230 2382 -162 2438
rect -106 2382 -38 2438
rect 18 2382 86 2438
rect 142 2382 210 2438
rect 266 2382 400 2438
rect -400 2314 400 2382
rect -400 2258 -286 2314
rect -230 2258 -162 2314
rect -106 2258 -38 2314
rect 18 2258 86 2314
rect 142 2258 210 2314
rect 266 2258 400 2314
rect -400 2190 400 2258
rect -400 2134 -286 2190
rect -230 2134 -162 2190
rect -106 2134 -38 2190
rect 18 2134 86 2190
rect 142 2134 210 2190
rect 266 2134 400 2190
rect -400 2066 400 2134
rect -400 2010 -286 2066
rect -230 2010 -162 2066
rect -106 2010 -38 2066
rect 18 2010 86 2066
rect 142 2010 210 2066
rect 266 2010 400 2066
rect -400 1942 400 2010
rect -400 1886 -286 1942
rect -230 1886 -162 1942
rect -106 1886 -38 1942
rect 18 1886 86 1942
rect 142 1886 210 1942
rect 266 1886 400 1942
rect -400 1818 400 1886
rect -400 1762 -286 1818
rect -230 1762 -162 1818
rect -106 1762 -38 1818
rect 18 1762 86 1818
rect 142 1762 210 1818
rect 266 1762 400 1818
rect -400 1694 400 1762
rect -400 1638 -286 1694
rect -230 1638 -162 1694
rect -106 1638 -38 1694
rect 18 1638 86 1694
rect 142 1638 210 1694
rect 266 1638 400 1694
rect -400 1570 400 1638
rect -400 1514 -286 1570
rect -230 1514 -162 1570
rect -106 1514 -38 1570
rect 18 1514 86 1570
rect 142 1514 210 1570
rect 266 1514 400 1570
rect -400 1446 400 1514
rect -400 1390 -286 1446
rect -230 1390 -162 1446
rect -106 1390 -38 1446
rect 18 1390 86 1446
rect 142 1390 210 1446
rect 266 1390 400 1446
rect -400 1322 400 1390
rect -400 1266 -286 1322
rect -230 1266 -162 1322
rect -106 1266 -38 1322
rect 18 1266 86 1322
rect 142 1266 210 1322
rect 266 1266 400 1322
rect -400 1198 400 1266
rect -400 1142 -286 1198
rect -230 1142 -162 1198
rect -106 1142 -38 1198
rect 18 1142 86 1198
rect 142 1142 210 1198
rect 266 1142 400 1198
rect -400 1074 400 1142
rect -400 1018 -286 1074
rect -230 1018 -162 1074
rect -106 1018 -38 1074
rect 18 1018 86 1074
rect 142 1018 210 1074
rect 266 1018 400 1074
rect -400 950 400 1018
rect -400 894 -286 950
rect -230 894 -162 950
rect -106 894 -38 950
rect 18 894 86 950
rect 142 894 210 950
rect 266 894 400 950
rect -400 826 400 894
rect -400 770 -286 826
rect -230 770 -162 826
rect -106 770 -38 826
rect 18 770 86 826
rect 142 770 210 826
rect 266 770 400 826
rect -400 702 400 770
rect -400 646 -286 702
rect -230 646 -162 702
rect -106 646 -38 702
rect 18 646 86 702
rect 142 646 210 702
rect 266 646 400 702
rect -400 578 400 646
rect -400 522 -286 578
rect -230 522 -162 578
rect -106 522 -38 578
rect 18 522 86 578
rect 142 522 210 578
rect 266 522 400 578
rect -400 454 400 522
rect -400 398 -286 454
rect -230 398 -162 454
rect -106 398 -38 454
rect 18 398 86 454
rect 142 398 210 454
rect 266 400 400 454
rect 830 12310 1170 12400
rect 830 12254 903 12310
rect 959 12254 1045 12310
rect 1101 12254 1170 12310
rect 830 12168 1170 12254
rect 830 12112 903 12168
rect 959 12112 1045 12168
rect 1101 12112 1170 12168
rect 830 12026 1170 12112
rect 830 11970 903 12026
rect 959 11970 1045 12026
rect 1101 11970 1170 12026
rect 830 11884 1170 11970
rect 830 11828 903 11884
rect 959 11828 1045 11884
rect 1101 11828 1170 11884
rect 830 11742 1170 11828
rect 830 11686 903 11742
rect 959 11686 1045 11742
rect 1101 11686 1170 11742
rect 830 11600 1170 11686
rect 830 11544 903 11600
rect 959 11544 1045 11600
rect 1101 11544 1170 11600
rect 830 11458 1170 11544
rect 830 11402 903 11458
rect 959 11402 1045 11458
rect 1101 11402 1170 11458
rect 830 11316 1170 11402
rect 830 11260 903 11316
rect 959 11260 1045 11316
rect 1101 11260 1170 11316
rect 830 11174 1170 11260
rect 830 11118 903 11174
rect 959 11118 1045 11174
rect 1101 11118 1170 11174
rect 830 11032 1170 11118
rect 830 10976 903 11032
rect 959 10976 1045 11032
rect 1101 10976 1170 11032
rect 830 10890 1170 10976
rect 830 10834 903 10890
rect 959 10834 1045 10890
rect 1101 10834 1170 10890
rect 830 10748 1170 10834
rect 830 10692 903 10748
rect 959 10692 1045 10748
rect 1101 10692 1170 10748
rect 830 10606 1170 10692
rect 830 10550 903 10606
rect 959 10550 1045 10606
rect 1101 10550 1170 10606
rect 830 10464 1170 10550
rect 830 10408 903 10464
rect 959 10408 1045 10464
rect 1101 10408 1170 10464
rect 830 10322 1170 10408
rect 830 10266 903 10322
rect 959 10266 1045 10322
rect 1101 10266 1170 10322
rect 830 10180 1170 10266
rect 830 10124 903 10180
rect 959 10124 1045 10180
rect 1101 10124 1170 10180
rect 830 10038 1170 10124
rect 830 9982 903 10038
rect 959 9982 1045 10038
rect 1101 9982 1170 10038
rect 830 9896 1170 9982
rect 830 9840 903 9896
rect 959 9840 1045 9896
rect 1101 9840 1170 9896
rect 830 9754 1170 9840
rect 830 9698 903 9754
rect 959 9698 1045 9754
rect 1101 9698 1170 9754
rect 830 9612 1170 9698
rect 830 9556 903 9612
rect 959 9556 1045 9612
rect 1101 9556 1170 9612
rect 830 9470 1170 9556
rect 830 9414 903 9470
rect 959 9414 1045 9470
rect 1101 9414 1170 9470
rect 830 9328 1170 9414
rect 830 9272 903 9328
rect 959 9272 1045 9328
rect 1101 9272 1170 9328
rect 830 9186 1170 9272
rect 830 9130 903 9186
rect 959 9130 1045 9186
rect 1101 9130 1170 9186
rect 830 9044 1170 9130
rect 830 8988 903 9044
rect 959 8988 1045 9044
rect 1101 8988 1170 9044
rect 830 8902 1170 8988
rect 830 8846 903 8902
rect 959 8846 1045 8902
rect 1101 8846 1170 8902
rect 830 8760 1170 8846
rect 830 8704 903 8760
rect 959 8704 1045 8760
rect 1101 8704 1170 8760
rect 830 8618 1170 8704
rect 830 8562 903 8618
rect 959 8562 1045 8618
rect 1101 8562 1170 8618
rect 830 8476 1170 8562
rect 830 8420 903 8476
rect 959 8420 1045 8476
rect 1101 8420 1170 8476
rect 830 8334 1170 8420
rect 830 8278 903 8334
rect 959 8278 1045 8334
rect 1101 8278 1170 8334
rect 830 8192 1170 8278
rect 830 8136 903 8192
rect 959 8136 1045 8192
rect 1101 8136 1170 8192
rect 830 8050 1170 8136
rect 830 7994 903 8050
rect 959 7994 1045 8050
rect 1101 7994 1170 8050
rect 830 7908 1170 7994
rect 830 7852 903 7908
rect 959 7852 1045 7908
rect 1101 7852 1170 7908
rect 830 7766 1170 7852
rect 830 7710 903 7766
rect 959 7710 1045 7766
rect 1101 7710 1170 7766
rect 830 7624 1170 7710
rect 830 7568 903 7624
rect 959 7568 1045 7624
rect 1101 7568 1170 7624
rect 830 7482 1170 7568
rect 830 7426 903 7482
rect 959 7426 1045 7482
rect 1101 7426 1170 7482
rect 830 7340 1170 7426
rect 830 7284 903 7340
rect 959 7284 1045 7340
rect 1101 7284 1170 7340
rect 830 7198 1170 7284
rect 830 7142 903 7198
rect 959 7142 1045 7198
rect 1101 7142 1170 7198
rect 830 7056 1170 7142
rect 830 7000 903 7056
rect 959 7000 1045 7056
rect 1101 7000 1170 7056
rect 830 6914 1170 7000
rect 830 6858 903 6914
rect 959 6858 1045 6914
rect 1101 6858 1170 6914
rect 830 6772 1170 6858
rect 830 6716 903 6772
rect 959 6716 1045 6772
rect 1101 6716 1170 6772
rect 830 6630 1170 6716
rect 830 6574 903 6630
rect 959 6574 1045 6630
rect 1101 6574 1170 6630
rect 830 6488 1170 6574
rect 830 6432 903 6488
rect 959 6432 1045 6488
rect 1101 6432 1170 6488
rect 830 6346 1170 6432
rect 830 6290 903 6346
rect 959 6290 1045 6346
rect 1101 6290 1170 6346
rect 830 6204 1170 6290
rect 830 6148 903 6204
rect 959 6148 1045 6204
rect 1101 6148 1170 6204
rect 830 6062 1170 6148
rect 830 6006 903 6062
rect 959 6006 1045 6062
rect 1101 6006 1170 6062
rect 830 5920 1170 6006
rect 830 5864 903 5920
rect 959 5864 1045 5920
rect 1101 5864 1170 5920
rect 830 5778 1170 5864
rect 830 5722 903 5778
rect 959 5722 1045 5778
rect 1101 5722 1170 5778
rect 830 5636 1170 5722
rect 830 5580 903 5636
rect 959 5580 1045 5636
rect 1101 5580 1170 5636
rect 830 5494 1170 5580
rect 830 5438 903 5494
rect 959 5438 1045 5494
rect 1101 5438 1170 5494
rect 830 5352 1170 5438
rect 830 5296 903 5352
rect 959 5296 1045 5352
rect 1101 5296 1170 5352
rect 830 5210 1170 5296
rect 830 5154 903 5210
rect 959 5154 1045 5210
rect 1101 5154 1170 5210
rect 830 5068 1170 5154
rect 830 5012 903 5068
rect 959 5012 1045 5068
rect 1101 5012 1170 5068
rect 830 4926 1170 5012
rect 830 4870 903 4926
rect 959 4870 1045 4926
rect 1101 4870 1170 4926
rect 830 4784 1170 4870
rect 830 4728 903 4784
rect 959 4728 1045 4784
rect 1101 4728 1170 4784
rect 830 4642 1170 4728
rect 830 4586 903 4642
rect 959 4586 1045 4642
rect 1101 4586 1170 4642
rect 830 4500 1170 4586
rect 830 4444 903 4500
rect 959 4444 1045 4500
rect 1101 4444 1170 4500
rect 830 4358 1170 4444
rect 830 4302 903 4358
rect 959 4302 1045 4358
rect 1101 4302 1170 4358
rect 830 4216 1170 4302
rect 830 4160 903 4216
rect 959 4160 1045 4216
rect 1101 4160 1170 4216
rect 830 4074 1170 4160
rect 830 4018 903 4074
rect 959 4018 1045 4074
rect 1101 4018 1170 4074
rect 830 3932 1170 4018
rect 830 3876 903 3932
rect 959 3876 1045 3932
rect 1101 3876 1170 3932
rect 830 3790 1170 3876
rect 830 3734 903 3790
rect 959 3734 1045 3790
rect 1101 3734 1170 3790
rect 830 3648 1170 3734
rect 830 3592 903 3648
rect 959 3592 1045 3648
rect 1101 3592 1170 3648
rect 830 3506 1170 3592
rect 830 3450 903 3506
rect 959 3450 1045 3506
rect 1101 3450 1170 3506
rect 830 3364 1170 3450
rect 830 3308 903 3364
rect 959 3308 1045 3364
rect 1101 3308 1170 3364
rect 830 3222 1170 3308
rect 830 3166 903 3222
rect 959 3166 1045 3222
rect 1101 3166 1170 3222
rect 830 3080 1170 3166
rect 830 3024 903 3080
rect 959 3024 1045 3080
rect 1101 3024 1170 3080
rect 830 2938 1170 3024
rect 830 2882 903 2938
rect 959 2882 1045 2938
rect 1101 2882 1170 2938
rect 830 2796 1170 2882
rect 830 2740 903 2796
rect 959 2740 1045 2796
rect 1101 2740 1170 2796
rect 830 2654 1170 2740
rect 830 2598 903 2654
rect 959 2598 1045 2654
rect 1101 2598 1170 2654
rect 830 2512 1170 2598
rect 830 2456 903 2512
rect 959 2456 1045 2512
rect 1101 2456 1170 2512
rect 830 2370 1170 2456
rect 830 2314 903 2370
rect 959 2314 1045 2370
rect 1101 2314 1170 2370
rect 830 2228 1170 2314
rect 830 2172 903 2228
rect 959 2172 1045 2228
rect 1101 2172 1170 2228
rect 830 2086 1170 2172
rect 830 2030 903 2086
rect 959 2030 1045 2086
rect 1101 2030 1170 2086
rect 830 1944 1170 2030
rect 830 1888 903 1944
rect 959 1888 1045 1944
rect 1101 1888 1170 1944
rect 830 1802 1170 1888
rect 830 1746 903 1802
rect 959 1746 1045 1802
rect 1101 1746 1170 1802
rect 830 1660 1170 1746
rect 830 1604 903 1660
rect 959 1604 1045 1660
rect 1101 1604 1170 1660
rect 830 1518 1170 1604
rect 830 1462 903 1518
rect 959 1462 1045 1518
rect 1101 1462 1170 1518
rect 830 1376 1170 1462
rect 830 1320 903 1376
rect 959 1320 1045 1376
rect 1101 1320 1170 1376
rect 830 1234 1170 1320
rect 830 1178 903 1234
rect 959 1178 1045 1234
rect 1101 1178 1170 1234
rect 830 1092 1170 1178
rect 830 1036 903 1092
rect 959 1036 1045 1092
rect 1101 1036 1170 1092
rect 830 950 1170 1036
rect 830 894 903 950
rect 959 894 1045 950
rect 1101 894 1170 950
rect 830 808 1170 894
rect 830 752 903 808
rect 959 752 1045 808
rect 1101 752 1170 808
rect 830 666 1170 752
rect 830 610 903 666
rect 959 610 1045 666
rect 1101 610 1170 666
rect 830 524 1170 610
rect 830 468 903 524
rect 959 468 1045 524
rect 1101 468 1170 524
rect 830 400 1170 468
rect 1370 12310 1710 12400
rect 1370 12254 1444 12310
rect 1500 12254 1586 12310
rect 1642 12254 1710 12310
rect 1370 12168 1710 12254
rect 1370 12112 1444 12168
rect 1500 12112 1586 12168
rect 1642 12112 1710 12168
rect 1370 12026 1710 12112
rect 1370 11970 1444 12026
rect 1500 11970 1586 12026
rect 1642 11970 1710 12026
rect 1370 11884 1710 11970
rect 1370 11828 1444 11884
rect 1500 11828 1586 11884
rect 1642 11828 1710 11884
rect 1370 11742 1710 11828
rect 1370 11686 1444 11742
rect 1500 11686 1586 11742
rect 1642 11686 1710 11742
rect 1370 11600 1710 11686
rect 1370 11544 1444 11600
rect 1500 11544 1586 11600
rect 1642 11544 1710 11600
rect 1370 11458 1710 11544
rect 1370 11402 1444 11458
rect 1500 11402 1586 11458
rect 1642 11402 1710 11458
rect 1370 11316 1710 11402
rect 1370 11260 1444 11316
rect 1500 11260 1586 11316
rect 1642 11260 1710 11316
rect 1370 11174 1710 11260
rect 1370 11118 1444 11174
rect 1500 11118 1586 11174
rect 1642 11118 1710 11174
rect 1370 11032 1710 11118
rect 1370 10976 1444 11032
rect 1500 10976 1586 11032
rect 1642 10976 1710 11032
rect 1370 10890 1710 10976
rect 1370 10834 1444 10890
rect 1500 10834 1586 10890
rect 1642 10834 1710 10890
rect 1370 10748 1710 10834
rect 1370 10692 1444 10748
rect 1500 10692 1586 10748
rect 1642 10692 1710 10748
rect 1370 10606 1710 10692
rect 1370 10550 1444 10606
rect 1500 10550 1586 10606
rect 1642 10550 1710 10606
rect 1370 10464 1710 10550
rect 1370 10408 1444 10464
rect 1500 10408 1586 10464
rect 1642 10408 1710 10464
rect 1370 10322 1710 10408
rect 1370 10266 1444 10322
rect 1500 10266 1586 10322
rect 1642 10266 1710 10322
rect 1370 10180 1710 10266
rect 1370 10124 1444 10180
rect 1500 10124 1586 10180
rect 1642 10124 1710 10180
rect 1370 10038 1710 10124
rect 1370 9982 1444 10038
rect 1500 9982 1586 10038
rect 1642 9982 1710 10038
rect 1370 9896 1710 9982
rect 1370 9840 1444 9896
rect 1500 9840 1586 9896
rect 1642 9840 1710 9896
rect 1370 9754 1710 9840
rect 1370 9698 1444 9754
rect 1500 9698 1586 9754
rect 1642 9698 1710 9754
rect 1370 9612 1710 9698
rect 1370 9556 1444 9612
rect 1500 9556 1586 9612
rect 1642 9556 1710 9612
rect 1370 9470 1710 9556
rect 1370 9414 1444 9470
rect 1500 9414 1586 9470
rect 1642 9414 1710 9470
rect 1370 9328 1710 9414
rect 1370 9272 1444 9328
rect 1500 9272 1586 9328
rect 1642 9272 1710 9328
rect 1370 9186 1710 9272
rect 1370 9130 1444 9186
rect 1500 9130 1586 9186
rect 1642 9130 1710 9186
rect 1370 9044 1710 9130
rect 1370 8988 1444 9044
rect 1500 8988 1586 9044
rect 1642 8988 1710 9044
rect 1370 8902 1710 8988
rect 1370 8846 1444 8902
rect 1500 8846 1586 8902
rect 1642 8846 1710 8902
rect 1370 8760 1710 8846
rect 1370 8704 1444 8760
rect 1500 8704 1586 8760
rect 1642 8704 1710 8760
rect 1370 8618 1710 8704
rect 1370 8562 1444 8618
rect 1500 8562 1586 8618
rect 1642 8562 1710 8618
rect 1370 8476 1710 8562
rect 1370 8420 1444 8476
rect 1500 8420 1586 8476
rect 1642 8420 1710 8476
rect 1370 8334 1710 8420
rect 1370 8278 1444 8334
rect 1500 8278 1586 8334
rect 1642 8278 1710 8334
rect 1370 8192 1710 8278
rect 1370 8136 1444 8192
rect 1500 8136 1586 8192
rect 1642 8136 1710 8192
rect 1370 8050 1710 8136
rect 1370 7994 1444 8050
rect 1500 7994 1586 8050
rect 1642 7994 1710 8050
rect 1370 7908 1710 7994
rect 1370 7852 1444 7908
rect 1500 7852 1586 7908
rect 1642 7852 1710 7908
rect 1370 7766 1710 7852
rect 1370 7710 1444 7766
rect 1500 7710 1586 7766
rect 1642 7710 1710 7766
rect 1370 7624 1710 7710
rect 1370 7568 1444 7624
rect 1500 7568 1586 7624
rect 1642 7568 1710 7624
rect 1370 7482 1710 7568
rect 1370 7426 1444 7482
rect 1500 7426 1586 7482
rect 1642 7426 1710 7482
rect 1370 7340 1710 7426
rect 1370 7284 1444 7340
rect 1500 7284 1586 7340
rect 1642 7284 1710 7340
rect 1370 7198 1710 7284
rect 1370 7142 1444 7198
rect 1500 7142 1586 7198
rect 1642 7142 1710 7198
rect 1370 7056 1710 7142
rect 1370 7000 1444 7056
rect 1500 7000 1586 7056
rect 1642 7000 1710 7056
rect 1370 6914 1710 7000
rect 1370 6858 1444 6914
rect 1500 6858 1586 6914
rect 1642 6858 1710 6914
rect 1370 6772 1710 6858
rect 1370 6716 1444 6772
rect 1500 6716 1586 6772
rect 1642 6716 1710 6772
rect 1370 6630 1710 6716
rect 1370 6574 1444 6630
rect 1500 6574 1586 6630
rect 1642 6574 1710 6630
rect 1370 6488 1710 6574
rect 1370 6432 1444 6488
rect 1500 6432 1586 6488
rect 1642 6432 1710 6488
rect 1370 6346 1710 6432
rect 1370 6290 1444 6346
rect 1500 6290 1586 6346
rect 1642 6290 1710 6346
rect 1370 6204 1710 6290
rect 1370 6148 1444 6204
rect 1500 6148 1586 6204
rect 1642 6148 1710 6204
rect 1370 6062 1710 6148
rect 1370 6006 1444 6062
rect 1500 6006 1586 6062
rect 1642 6006 1710 6062
rect 1370 5920 1710 6006
rect 1370 5864 1444 5920
rect 1500 5864 1586 5920
rect 1642 5864 1710 5920
rect 1370 5778 1710 5864
rect 1370 5722 1444 5778
rect 1500 5722 1586 5778
rect 1642 5722 1710 5778
rect 1370 5636 1710 5722
rect 1370 5580 1444 5636
rect 1500 5580 1586 5636
rect 1642 5580 1710 5636
rect 1370 5494 1710 5580
rect 1370 5438 1444 5494
rect 1500 5438 1586 5494
rect 1642 5438 1710 5494
rect 1370 5352 1710 5438
rect 1370 5296 1444 5352
rect 1500 5296 1586 5352
rect 1642 5296 1710 5352
rect 1370 5210 1710 5296
rect 1370 5154 1444 5210
rect 1500 5154 1586 5210
rect 1642 5154 1710 5210
rect 1370 5068 1710 5154
rect 1370 5012 1444 5068
rect 1500 5012 1586 5068
rect 1642 5012 1710 5068
rect 1370 4926 1710 5012
rect 1370 4870 1444 4926
rect 1500 4870 1586 4926
rect 1642 4870 1710 4926
rect 1370 4784 1710 4870
rect 1370 4728 1444 4784
rect 1500 4728 1586 4784
rect 1642 4728 1710 4784
rect 1370 4642 1710 4728
rect 1370 4586 1444 4642
rect 1500 4586 1586 4642
rect 1642 4586 1710 4642
rect 1370 4500 1710 4586
rect 1370 4444 1444 4500
rect 1500 4444 1586 4500
rect 1642 4444 1710 4500
rect 1370 4358 1710 4444
rect 1370 4302 1444 4358
rect 1500 4302 1586 4358
rect 1642 4302 1710 4358
rect 1370 4216 1710 4302
rect 1370 4160 1444 4216
rect 1500 4160 1586 4216
rect 1642 4160 1710 4216
rect 1370 4074 1710 4160
rect 1370 4018 1444 4074
rect 1500 4018 1586 4074
rect 1642 4018 1710 4074
rect 1370 3932 1710 4018
rect 1370 3876 1444 3932
rect 1500 3876 1586 3932
rect 1642 3876 1710 3932
rect 1370 3790 1710 3876
rect 1370 3734 1444 3790
rect 1500 3734 1586 3790
rect 1642 3734 1710 3790
rect 1370 3648 1710 3734
rect 1370 3592 1444 3648
rect 1500 3592 1586 3648
rect 1642 3592 1710 3648
rect 1370 3506 1710 3592
rect 1370 3450 1444 3506
rect 1500 3450 1586 3506
rect 1642 3450 1710 3506
rect 1370 3364 1710 3450
rect 1370 3308 1444 3364
rect 1500 3308 1586 3364
rect 1642 3308 1710 3364
rect 1370 3222 1710 3308
rect 1370 3166 1444 3222
rect 1500 3166 1586 3222
rect 1642 3166 1710 3222
rect 1370 3080 1710 3166
rect 1370 3024 1444 3080
rect 1500 3024 1586 3080
rect 1642 3024 1710 3080
rect 1370 2938 1710 3024
rect 1370 2882 1444 2938
rect 1500 2882 1586 2938
rect 1642 2882 1710 2938
rect 1370 2796 1710 2882
rect 1370 2740 1444 2796
rect 1500 2740 1586 2796
rect 1642 2740 1710 2796
rect 1370 2654 1710 2740
rect 1370 2598 1444 2654
rect 1500 2598 1586 2654
rect 1642 2598 1710 2654
rect 1370 2512 1710 2598
rect 1370 2456 1444 2512
rect 1500 2456 1586 2512
rect 1642 2456 1710 2512
rect 1370 2370 1710 2456
rect 1370 2314 1444 2370
rect 1500 2314 1586 2370
rect 1642 2314 1710 2370
rect 1370 2228 1710 2314
rect 1370 2172 1444 2228
rect 1500 2172 1586 2228
rect 1642 2172 1710 2228
rect 1370 2086 1710 2172
rect 1370 2030 1444 2086
rect 1500 2030 1586 2086
rect 1642 2030 1710 2086
rect 1370 1944 1710 2030
rect 1370 1888 1444 1944
rect 1500 1888 1586 1944
rect 1642 1888 1710 1944
rect 1370 1802 1710 1888
rect 1370 1746 1444 1802
rect 1500 1746 1586 1802
rect 1642 1746 1710 1802
rect 1370 1660 1710 1746
rect 1370 1604 1444 1660
rect 1500 1604 1586 1660
rect 1642 1604 1710 1660
rect 1370 1518 1710 1604
rect 1370 1462 1444 1518
rect 1500 1462 1586 1518
rect 1642 1462 1710 1518
rect 1370 1376 1710 1462
rect 1370 1320 1444 1376
rect 1500 1320 1586 1376
rect 1642 1320 1710 1376
rect 1370 1234 1710 1320
rect 1370 1178 1444 1234
rect 1500 1178 1586 1234
rect 1642 1178 1710 1234
rect 1370 1092 1710 1178
rect 1370 1036 1444 1092
rect 1500 1036 1586 1092
rect 1642 1036 1710 1092
rect 1370 950 1710 1036
rect 1370 894 1444 950
rect 1500 894 1586 950
rect 1642 894 1710 950
rect 1370 808 1710 894
rect 1370 752 1444 808
rect 1500 752 1586 808
rect 1642 752 1710 808
rect 1370 666 1710 752
rect 1370 610 1444 666
rect 1500 610 1586 666
rect 1642 610 1710 666
rect 1370 524 1710 610
rect 1370 468 1444 524
rect 1500 468 1586 524
rect 1642 468 1710 524
rect 1370 400 1710 468
rect 1910 12310 2250 12400
rect 1910 12254 1984 12310
rect 2040 12254 2126 12310
rect 2182 12254 2250 12310
rect 1910 12168 2250 12254
rect 1910 12112 1984 12168
rect 2040 12112 2126 12168
rect 2182 12112 2250 12168
rect 1910 12026 2250 12112
rect 1910 11970 1984 12026
rect 2040 11970 2126 12026
rect 2182 11970 2250 12026
rect 1910 11884 2250 11970
rect 1910 11828 1984 11884
rect 2040 11828 2126 11884
rect 2182 11828 2250 11884
rect 1910 11742 2250 11828
rect 1910 11686 1984 11742
rect 2040 11686 2126 11742
rect 2182 11686 2250 11742
rect 1910 11600 2250 11686
rect 1910 11544 1984 11600
rect 2040 11544 2126 11600
rect 2182 11544 2250 11600
rect 1910 11458 2250 11544
rect 1910 11402 1984 11458
rect 2040 11402 2126 11458
rect 2182 11402 2250 11458
rect 1910 11316 2250 11402
rect 1910 11260 1984 11316
rect 2040 11260 2126 11316
rect 2182 11260 2250 11316
rect 1910 11174 2250 11260
rect 1910 11118 1984 11174
rect 2040 11118 2126 11174
rect 2182 11118 2250 11174
rect 1910 11032 2250 11118
rect 1910 10976 1984 11032
rect 2040 10976 2126 11032
rect 2182 10976 2250 11032
rect 1910 10890 2250 10976
rect 1910 10834 1984 10890
rect 2040 10834 2126 10890
rect 2182 10834 2250 10890
rect 1910 10748 2250 10834
rect 1910 10692 1984 10748
rect 2040 10692 2126 10748
rect 2182 10692 2250 10748
rect 1910 10606 2250 10692
rect 1910 10550 1984 10606
rect 2040 10550 2126 10606
rect 2182 10550 2250 10606
rect 1910 10464 2250 10550
rect 1910 10408 1984 10464
rect 2040 10408 2126 10464
rect 2182 10408 2250 10464
rect 1910 10322 2250 10408
rect 1910 10266 1984 10322
rect 2040 10266 2126 10322
rect 2182 10266 2250 10322
rect 1910 10180 2250 10266
rect 1910 10124 1984 10180
rect 2040 10124 2126 10180
rect 2182 10124 2250 10180
rect 1910 10038 2250 10124
rect 1910 9982 1984 10038
rect 2040 9982 2126 10038
rect 2182 9982 2250 10038
rect 1910 9896 2250 9982
rect 1910 9840 1984 9896
rect 2040 9840 2126 9896
rect 2182 9840 2250 9896
rect 1910 9754 2250 9840
rect 1910 9698 1984 9754
rect 2040 9698 2126 9754
rect 2182 9698 2250 9754
rect 1910 9612 2250 9698
rect 1910 9556 1984 9612
rect 2040 9556 2126 9612
rect 2182 9556 2250 9612
rect 1910 9470 2250 9556
rect 1910 9414 1984 9470
rect 2040 9414 2126 9470
rect 2182 9414 2250 9470
rect 1910 9328 2250 9414
rect 1910 9272 1984 9328
rect 2040 9272 2126 9328
rect 2182 9272 2250 9328
rect 1910 9186 2250 9272
rect 1910 9130 1984 9186
rect 2040 9130 2126 9186
rect 2182 9130 2250 9186
rect 1910 9044 2250 9130
rect 1910 8988 1984 9044
rect 2040 8988 2126 9044
rect 2182 8988 2250 9044
rect 1910 8902 2250 8988
rect 1910 8846 1984 8902
rect 2040 8846 2126 8902
rect 2182 8846 2250 8902
rect 1910 8760 2250 8846
rect 1910 8704 1984 8760
rect 2040 8704 2126 8760
rect 2182 8704 2250 8760
rect 1910 8618 2250 8704
rect 1910 8562 1984 8618
rect 2040 8562 2126 8618
rect 2182 8562 2250 8618
rect 1910 8476 2250 8562
rect 1910 8420 1984 8476
rect 2040 8420 2126 8476
rect 2182 8420 2250 8476
rect 1910 8334 2250 8420
rect 1910 8278 1984 8334
rect 2040 8278 2126 8334
rect 2182 8278 2250 8334
rect 1910 8192 2250 8278
rect 1910 8136 1984 8192
rect 2040 8136 2126 8192
rect 2182 8136 2250 8192
rect 1910 8050 2250 8136
rect 1910 7994 1984 8050
rect 2040 7994 2126 8050
rect 2182 7994 2250 8050
rect 1910 7908 2250 7994
rect 1910 7852 1984 7908
rect 2040 7852 2126 7908
rect 2182 7852 2250 7908
rect 1910 7766 2250 7852
rect 1910 7710 1984 7766
rect 2040 7710 2126 7766
rect 2182 7710 2250 7766
rect 1910 7624 2250 7710
rect 1910 7568 1984 7624
rect 2040 7568 2126 7624
rect 2182 7568 2250 7624
rect 1910 7482 2250 7568
rect 1910 7426 1984 7482
rect 2040 7426 2126 7482
rect 2182 7426 2250 7482
rect 1910 7340 2250 7426
rect 1910 7284 1984 7340
rect 2040 7284 2126 7340
rect 2182 7284 2250 7340
rect 1910 7198 2250 7284
rect 1910 7142 1984 7198
rect 2040 7142 2126 7198
rect 2182 7142 2250 7198
rect 1910 7056 2250 7142
rect 1910 7000 1984 7056
rect 2040 7000 2126 7056
rect 2182 7000 2250 7056
rect 1910 6914 2250 7000
rect 1910 6858 1984 6914
rect 2040 6858 2126 6914
rect 2182 6858 2250 6914
rect 1910 6772 2250 6858
rect 1910 6716 1984 6772
rect 2040 6716 2126 6772
rect 2182 6716 2250 6772
rect 1910 6630 2250 6716
rect 1910 6574 1984 6630
rect 2040 6574 2126 6630
rect 2182 6574 2250 6630
rect 1910 6488 2250 6574
rect 1910 6432 1984 6488
rect 2040 6432 2126 6488
rect 2182 6432 2250 6488
rect 1910 6346 2250 6432
rect 1910 6290 1984 6346
rect 2040 6290 2126 6346
rect 2182 6290 2250 6346
rect 1910 6204 2250 6290
rect 1910 6148 1984 6204
rect 2040 6148 2126 6204
rect 2182 6148 2250 6204
rect 1910 6062 2250 6148
rect 1910 6006 1984 6062
rect 2040 6006 2126 6062
rect 2182 6006 2250 6062
rect 1910 5920 2250 6006
rect 1910 5864 1984 5920
rect 2040 5864 2126 5920
rect 2182 5864 2250 5920
rect 1910 5778 2250 5864
rect 1910 5722 1984 5778
rect 2040 5722 2126 5778
rect 2182 5722 2250 5778
rect 1910 5636 2250 5722
rect 1910 5580 1984 5636
rect 2040 5580 2126 5636
rect 2182 5580 2250 5636
rect 1910 5494 2250 5580
rect 1910 5438 1984 5494
rect 2040 5438 2126 5494
rect 2182 5438 2250 5494
rect 1910 5352 2250 5438
rect 1910 5296 1984 5352
rect 2040 5296 2126 5352
rect 2182 5296 2250 5352
rect 1910 5210 2250 5296
rect 1910 5154 1984 5210
rect 2040 5154 2126 5210
rect 2182 5154 2250 5210
rect 1910 5068 2250 5154
rect 1910 5012 1984 5068
rect 2040 5012 2126 5068
rect 2182 5012 2250 5068
rect 1910 4926 2250 5012
rect 1910 4870 1984 4926
rect 2040 4870 2126 4926
rect 2182 4870 2250 4926
rect 1910 4784 2250 4870
rect 1910 4728 1984 4784
rect 2040 4728 2126 4784
rect 2182 4728 2250 4784
rect 1910 4642 2250 4728
rect 1910 4586 1984 4642
rect 2040 4586 2126 4642
rect 2182 4586 2250 4642
rect 1910 4500 2250 4586
rect 1910 4444 1984 4500
rect 2040 4444 2126 4500
rect 2182 4444 2250 4500
rect 1910 4358 2250 4444
rect 1910 4302 1984 4358
rect 2040 4302 2126 4358
rect 2182 4302 2250 4358
rect 1910 4216 2250 4302
rect 1910 4160 1984 4216
rect 2040 4160 2126 4216
rect 2182 4160 2250 4216
rect 1910 4074 2250 4160
rect 1910 4018 1984 4074
rect 2040 4018 2126 4074
rect 2182 4018 2250 4074
rect 1910 3932 2250 4018
rect 1910 3876 1984 3932
rect 2040 3876 2126 3932
rect 2182 3876 2250 3932
rect 1910 3790 2250 3876
rect 1910 3734 1984 3790
rect 2040 3734 2126 3790
rect 2182 3734 2250 3790
rect 1910 3648 2250 3734
rect 1910 3592 1984 3648
rect 2040 3592 2126 3648
rect 2182 3592 2250 3648
rect 1910 3506 2250 3592
rect 1910 3450 1984 3506
rect 2040 3450 2126 3506
rect 2182 3450 2250 3506
rect 1910 3364 2250 3450
rect 1910 3308 1984 3364
rect 2040 3308 2126 3364
rect 2182 3308 2250 3364
rect 1910 3222 2250 3308
rect 1910 3166 1984 3222
rect 2040 3166 2126 3222
rect 2182 3166 2250 3222
rect 1910 3080 2250 3166
rect 1910 3024 1984 3080
rect 2040 3024 2126 3080
rect 2182 3024 2250 3080
rect 1910 2938 2250 3024
rect 1910 2882 1984 2938
rect 2040 2882 2126 2938
rect 2182 2882 2250 2938
rect 1910 2796 2250 2882
rect 1910 2740 1984 2796
rect 2040 2740 2126 2796
rect 2182 2740 2250 2796
rect 1910 2654 2250 2740
rect 1910 2598 1984 2654
rect 2040 2598 2126 2654
rect 2182 2598 2250 2654
rect 1910 2512 2250 2598
rect 1910 2456 1984 2512
rect 2040 2456 2126 2512
rect 2182 2456 2250 2512
rect 1910 2370 2250 2456
rect 1910 2314 1984 2370
rect 2040 2314 2126 2370
rect 2182 2314 2250 2370
rect 1910 2228 2250 2314
rect 1910 2172 1984 2228
rect 2040 2172 2126 2228
rect 2182 2172 2250 2228
rect 1910 2086 2250 2172
rect 1910 2030 1984 2086
rect 2040 2030 2126 2086
rect 2182 2030 2250 2086
rect 1910 1944 2250 2030
rect 1910 1888 1984 1944
rect 2040 1888 2126 1944
rect 2182 1888 2250 1944
rect 1910 1802 2250 1888
rect 1910 1746 1984 1802
rect 2040 1746 2126 1802
rect 2182 1746 2250 1802
rect 1910 1660 2250 1746
rect 1910 1604 1984 1660
rect 2040 1604 2126 1660
rect 2182 1604 2250 1660
rect 1910 1518 2250 1604
rect 1910 1462 1984 1518
rect 2040 1462 2126 1518
rect 2182 1462 2250 1518
rect 1910 1376 2250 1462
rect 1910 1320 1984 1376
rect 2040 1320 2126 1376
rect 2182 1320 2250 1376
rect 1910 1234 2250 1320
rect 1910 1178 1984 1234
rect 2040 1178 2126 1234
rect 2182 1178 2250 1234
rect 1910 1092 2250 1178
rect 1910 1036 1984 1092
rect 2040 1036 2126 1092
rect 2182 1036 2250 1092
rect 1910 950 2250 1036
rect 1910 894 1984 950
rect 2040 894 2126 950
rect 2182 894 2250 950
rect 1910 808 2250 894
rect 1910 752 1984 808
rect 2040 752 2126 808
rect 2182 752 2250 808
rect 1910 666 2250 752
rect 1910 610 1984 666
rect 2040 610 2126 666
rect 2182 610 2250 666
rect 1910 524 2250 610
rect 1910 468 1984 524
rect 2040 468 2126 524
rect 2182 468 2250 524
rect 1910 400 2250 468
rect 2450 12310 2790 12400
rect 2450 12254 2521 12310
rect 2577 12254 2663 12310
rect 2719 12254 2790 12310
rect 2450 12168 2790 12254
rect 2450 12112 2521 12168
rect 2577 12112 2663 12168
rect 2719 12112 2790 12168
rect 2450 12026 2790 12112
rect 2450 11970 2521 12026
rect 2577 11970 2663 12026
rect 2719 11970 2790 12026
rect 2450 11884 2790 11970
rect 2450 11828 2521 11884
rect 2577 11828 2663 11884
rect 2719 11828 2790 11884
rect 2450 11742 2790 11828
rect 2450 11686 2521 11742
rect 2577 11686 2663 11742
rect 2719 11686 2790 11742
rect 2450 11600 2790 11686
rect 2450 11544 2521 11600
rect 2577 11544 2663 11600
rect 2719 11544 2790 11600
rect 2450 11458 2790 11544
rect 2450 11402 2521 11458
rect 2577 11402 2663 11458
rect 2719 11402 2790 11458
rect 2450 11316 2790 11402
rect 2450 11260 2521 11316
rect 2577 11260 2663 11316
rect 2719 11260 2790 11316
rect 2450 11174 2790 11260
rect 2450 11118 2521 11174
rect 2577 11118 2663 11174
rect 2719 11118 2790 11174
rect 2450 11032 2790 11118
rect 2450 10976 2521 11032
rect 2577 10976 2663 11032
rect 2719 10976 2790 11032
rect 2450 10890 2790 10976
rect 2450 10834 2521 10890
rect 2577 10834 2663 10890
rect 2719 10834 2790 10890
rect 2450 10748 2790 10834
rect 2450 10692 2521 10748
rect 2577 10692 2663 10748
rect 2719 10692 2790 10748
rect 2450 10606 2790 10692
rect 2450 10550 2521 10606
rect 2577 10550 2663 10606
rect 2719 10550 2790 10606
rect 2450 10464 2790 10550
rect 2450 10408 2521 10464
rect 2577 10408 2663 10464
rect 2719 10408 2790 10464
rect 2450 10322 2790 10408
rect 2450 10266 2521 10322
rect 2577 10266 2663 10322
rect 2719 10266 2790 10322
rect 2450 10180 2790 10266
rect 2450 10124 2521 10180
rect 2577 10124 2663 10180
rect 2719 10124 2790 10180
rect 2450 10038 2790 10124
rect 2450 9982 2521 10038
rect 2577 9982 2663 10038
rect 2719 9982 2790 10038
rect 2450 9896 2790 9982
rect 2450 9840 2521 9896
rect 2577 9840 2663 9896
rect 2719 9840 2790 9896
rect 2450 9754 2790 9840
rect 2450 9698 2521 9754
rect 2577 9698 2663 9754
rect 2719 9698 2790 9754
rect 2450 9612 2790 9698
rect 2450 9556 2521 9612
rect 2577 9556 2663 9612
rect 2719 9556 2790 9612
rect 2450 9470 2790 9556
rect 2450 9414 2521 9470
rect 2577 9414 2663 9470
rect 2719 9414 2790 9470
rect 2450 9328 2790 9414
rect 2450 9272 2521 9328
rect 2577 9272 2663 9328
rect 2719 9272 2790 9328
rect 2450 9186 2790 9272
rect 2450 9130 2521 9186
rect 2577 9130 2663 9186
rect 2719 9130 2790 9186
rect 2450 9044 2790 9130
rect 2450 8988 2521 9044
rect 2577 8988 2663 9044
rect 2719 8988 2790 9044
rect 2450 8902 2790 8988
rect 2450 8846 2521 8902
rect 2577 8846 2663 8902
rect 2719 8846 2790 8902
rect 2450 8760 2790 8846
rect 2450 8704 2521 8760
rect 2577 8704 2663 8760
rect 2719 8704 2790 8760
rect 2450 8618 2790 8704
rect 2450 8562 2521 8618
rect 2577 8562 2663 8618
rect 2719 8562 2790 8618
rect 2450 8476 2790 8562
rect 2450 8420 2521 8476
rect 2577 8420 2663 8476
rect 2719 8420 2790 8476
rect 2450 8334 2790 8420
rect 2450 8278 2521 8334
rect 2577 8278 2663 8334
rect 2719 8278 2790 8334
rect 2450 8192 2790 8278
rect 2450 8136 2521 8192
rect 2577 8136 2663 8192
rect 2719 8136 2790 8192
rect 2450 8050 2790 8136
rect 2450 7994 2521 8050
rect 2577 7994 2663 8050
rect 2719 7994 2790 8050
rect 2450 7908 2790 7994
rect 2450 7852 2521 7908
rect 2577 7852 2663 7908
rect 2719 7852 2790 7908
rect 2450 7766 2790 7852
rect 2450 7710 2521 7766
rect 2577 7710 2663 7766
rect 2719 7710 2790 7766
rect 2450 7624 2790 7710
rect 2450 7568 2521 7624
rect 2577 7568 2663 7624
rect 2719 7568 2790 7624
rect 2450 7482 2790 7568
rect 2450 7426 2521 7482
rect 2577 7426 2663 7482
rect 2719 7426 2790 7482
rect 2450 7340 2790 7426
rect 2450 7284 2521 7340
rect 2577 7284 2663 7340
rect 2719 7284 2790 7340
rect 2450 7198 2790 7284
rect 2450 7142 2521 7198
rect 2577 7142 2663 7198
rect 2719 7142 2790 7198
rect 2450 7056 2790 7142
rect 2450 7000 2521 7056
rect 2577 7000 2663 7056
rect 2719 7000 2790 7056
rect 2450 6914 2790 7000
rect 2450 6858 2521 6914
rect 2577 6858 2663 6914
rect 2719 6858 2790 6914
rect 2450 6772 2790 6858
rect 2450 6716 2521 6772
rect 2577 6716 2663 6772
rect 2719 6716 2790 6772
rect 2450 6630 2790 6716
rect 2450 6574 2521 6630
rect 2577 6574 2663 6630
rect 2719 6574 2790 6630
rect 2450 6488 2790 6574
rect 2450 6432 2521 6488
rect 2577 6432 2663 6488
rect 2719 6432 2790 6488
rect 2450 6346 2790 6432
rect 2450 6290 2521 6346
rect 2577 6290 2663 6346
rect 2719 6290 2790 6346
rect 2450 6204 2790 6290
rect 2450 6148 2521 6204
rect 2577 6148 2663 6204
rect 2719 6148 2790 6204
rect 2450 6062 2790 6148
rect 2450 6006 2521 6062
rect 2577 6006 2663 6062
rect 2719 6006 2790 6062
rect 2450 5920 2790 6006
rect 2450 5864 2521 5920
rect 2577 5864 2663 5920
rect 2719 5864 2790 5920
rect 2450 5778 2790 5864
rect 2450 5722 2521 5778
rect 2577 5722 2663 5778
rect 2719 5722 2790 5778
rect 2450 5636 2790 5722
rect 2450 5580 2521 5636
rect 2577 5580 2663 5636
rect 2719 5580 2790 5636
rect 2450 5494 2790 5580
rect 2450 5438 2521 5494
rect 2577 5438 2663 5494
rect 2719 5438 2790 5494
rect 2450 5352 2790 5438
rect 2450 5296 2521 5352
rect 2577 5296 2663 5352
rect 2719 5296 2790 5352
rect 2450 5210 2790 5296
rect 2450 5154 2521 5210
rect 2577 5154 2663 5210
rect 2719 5154 2790 5210
rect 2450 5068 2790 5154
rect 2450 5012 2521 5068
rect 2577 5012 2663 5068
rect 2719 5012 2790 5068
rect 2450 4926 2790 5012
rect 2450 4870 2521 4926
rect 2577 4870 2663 4926
rect 2719 4870 2790 4926
rect 2450 4784 2790 4870
rect 2450 4728 2521 4784
rect 2577 4728 2663 4784
rect 2719 4728 2790 4784
rect 2450 4642 2790 4728
rect 2450 4586 2521 4642
rect 2577 4586 2663 4642
rect 2719 4586 2790 4642
rect 2450 4500 2790 4586
rect 2450 4444 2521 4500
rect 2577 4444 2663 4500
rect 2719 4444 2790 4500
rect 2450 4358 2790 4444
rect 2450 4302 2521 4358
rect 2577 4302 2663 4358
rect 2719 4302 2790 4358
rect 2450 4216 2790 4302
rect 2450 4160 2521 4216
rect 2577 4160 2663 4216
rect 2719 4160 2790 4216
rect 2450 4074 2790 4160
rect 2450 4018 2521 4074
rect 2577 4018 2663 4074
rect 2719 4018 2790 4074
rect 2450 3932 2790 4018
rect 2450 3876 2521 3932
rect 2577 3876 2663 3932
rect 2719 3876 2790 3932
rect 2450 3790 2790 3876
rect 2450 3734 2521 3790
rect 2577 3734 2663 3790
rect 2719 3734 2790 3790
rect 2450 3648 2790 3734
rect 2450 3592 2521 3648
rect 2577 3592 2663 3648
rect 2719 3592 2790 3648
rect 2450 3506 2790 3592
rect 2450 3450 2521 3506
rect 2577 3450 2663 3506
rect 2719 3450 2790 3506
rect 2450 3364 2790 3450
rect 2450 3308 2521 3364
rect 2577 3308 2663 3364
rect 2719 3308 2790 3364
rect 2450 3222 2790 3308
rect 2450 3166 2521 3222
rect 2577 3166 2663 3222
rect 2719 3166 2790 3222
rect 2450 3080 2790 3166
rect 2450 3024 2521 3080
rect 2577 3024 2663 3080
rect 2719 3024 2790 3080
rect 2450 2938 2790 3024
rect 2450 2882 2521 2938
rect 2577 2882 2663 2938
rect 2719 2882 2790 2938
rect 2450 2796 2790 2882
rect 2450 2740 2521 2796
rect 2577 2740 2663 2796
rect 2719 2740 2790 2796
rect 2450 2654 2790 2740
rect 2450 2598 2521 2654
rect 2577 2598 2663 2654
rect 2719 2598 2790 2654
rect 2450 2512 2790 2598
rect 2450 2456 2521 2512
rect 2577 2456 2663 2512
rect 2719 2456 2790 2512
rect 2450 2370 2790 2456
rect 2450 2314 2521 2370
rect 2577 2314 2663 2370
rect 2719 2314 2790 2370
rect 2450 2228 2790 2314
rect 2450 2172 2521 2228
rect 2577 2172 2663 2228
rect 2719 2172 2790 2228
rect 2450 2086 2790 2172
rect 2450 2030 2521 2086
rect 2577 2030 2663 2086
rect 2719 2030 2790 2086
rect 2450 1944 2790 2030
rect 2450 1888 2521 1944
rect 2577 1888 2663 1944
rect 2719 1888 2790 1944
rect 2450 1802 2790 1888
rect 2450 1746 2521 1802
rect 2577 1746 2663 1802
rect 2719 1746 2790 1802
rect 2450 1660 2790 1746
rect 2450 1604 2521 1660
rect 2577 1604 2663 1660
rect 2719 1604 2790 1660
rect 2450 1518 2790 1604
rect 2450 1462 2521 1518
rect 2577 1462 2663 1518
rect 2719 1462 2790 1518
rect 2450 1376 2790 1462
rect 2450 1320 2521 1376
rect 2577 1320 2663 1376
rect 2719 1320 2790 1376
rect 2450 1234 2790 1320
rect 2450 1178 2521 1234
rect 2577 1178 2663 1234
rect 2719 1178 2790 1234
rect 2450 1092 2790 1178
rect 2450 1036 2521 1092
rect 2577 1036 2663 1092
rect 2719 1036 2790 1092
rect 2450 950 2790 1036
rect 2450 894 2521 950
rect 2577 894 2663 950
rect 2719 894 2790 950
rect 2450 808 2790 894
rect 2450 752 2521 808
rect 2577 752 2663 808
rect 2719 752 2790 808
rect 2450 666 2790 752
rect 2450 610 2521 666
rect 2577 610 2663 666
rect 2719 610 2790 666
rect 2450 524 2790 610
rect 2450 468 2521 524
rect 2577 468 2663 524
rect 2719 468 2790 524
rect 2450 400 2790 468
rect 2990 12310 3330 12400
rect 2990 12254 3058 12310
rect 3114 12254 3200 12310
rect 3256 12254 3330 12310
rect 2990 12168 3330 12254
rect 2990 12112 3058 12168
rect 3114 12112 3200 12168
rect 3256 12112 3330 12168
rect 2990 12026 3330 12112
rect 2990 11970 3058 12026
rect 3114 11970 3200 12026
rect 3256 11970 3330 12026
rect 2990 11884 3330 11970
rect 2990 11828 3058 11884
rect 3114 11828 3200 11884
rect 3256 11828 3330 11884
rect 2990 11742 3330 11828
rect 2990 11686 3058 11742
rect 3114 11686 3200 11742
rect 3256 11686 3330 11742
rect 2990 11600 3330 11686
rect 2990 11544 3058 11600
rect 3114 11544 3200 11600
rect 3256 11544 3330 11600
rect 2990 11458 3330 11544
rect 2990 11402 3058 11458
rect 3114 11402 3200 11458
rect 3256 11402 3330 11458
rect 2990 11316 3330 11402
rect 2990 11260 3058 11316
rect 3114 11260 3200 11316
rect 3256 11260 3330 11316
rect 2990 11174 3330 11260
rect 2990 11118 3058 11174
rect 3114 11118 3200 11174
rect 3256 11118 3330 11174
rect 2990 11032 3330 11118
rect 2990 10976 3058 11032
rect 3114 10976 3200 11032
rect 3256 10976 3330 11032
rect 2990 10890 3330 10976
rect 2990 10834 3058 10890
rect 3114 10834 3200 10890
rect 3256 10834 3330 10890
rect 2990 10748 3330 10834
rect 2990 10692 3058 10748
rect 3114 10692 3200 10748
rect 3256 10692 3330 10748
rect 2990 10606 3330 10692
rect 2990 10550 3058 10606
rect 3114 10550 3200 10606
rect 3256 10550 3330 10606
rect 2990 10464 3330 10550
rect 2990 10408 3058 10464
rect 3114 10408 3200 10464
rect 3256 10408 3330 10464
rect 2990 10322 3330 10408
rect 2990 10266 3058 10322
rect 3114 10266 3200 10322
rect 3256 10266 3330 10322
rect 2990 10180 3330 10266
rect 2990 10124 3058 10180
rect 3114 10124 3200 10180
rect 3256 10124 3330 10180
rect 2990 10038 3330 10124
rect 2990 9982 3058 10038
rect 3114 9982 3200 10038
rect 3256 9982 3330 10038
rect 2990 9896 3330 9982
rect 2990 9840 3058 9896
rect 3114 9840 3200 9896
rect 3256 9840 3330 9896
rect 2990 9754 3330 9840
rect 2990 9698 3058 9754
rect 3114 9698 3200 9754
rect 3256 9698 3330 9754
rect 2990 9612 3330 9698
rect 2990 9556 3058 9612
rect 3114 9556 3200 9612
rect 3256 9556 3330 9612
rect 2990 9470 3330 9556
rect 2990 9414 3058 9470
rect 3114 9414 3200 9470
rect 3256 9414 3330 9470
rect 2990 9328 3330 9414
rect 2990 9272 3058 9328
rect 3114 9272 3200 9328
rect 3256 9272 3330 9328
rect 2990 9186 3330 9272
rect 2990 9130 3058 9186
rect 3114 9130 3200 9186
rect 3256 9130 3330 9186
rect 2990 9044 3330 9130
rect 2990 8988 3058 9044
rect 3114 8988 3200 9044
rect 3256 8988 3330 9044
rect 2990 8902 3330 8988
rect 2990 8846 3058 8902
rect 3114 8846 3200 8902
rect 3256 8846 3330 8902
rect 2990 8760 3330 8846
rect 2990 8704 3058 8760
rect 3114 8704 3200 8760
rect 3256 8704 3330 8760
rect 2990 8618 3330 8704
rect 2990 8562 3058 8618
rect 3114 8562 3200 8618
rect 3256 8562 3330 8618
rect 2990 8476 3330 8562
rect 2990 8420 3058 8476
rect 3114 8420 3200 8476
rect 3256 8420 3330 8476
rect 2990 8334 3330 8420
rect 2990 8278 3058 8334
rect 3114 8278 3200 8334
rect 3256 8278 3330 8334
rect 2990 8192 3330 8278
rect 2990 8136 3058 8192
rect 3114 8136 3200 8192
rect 3256 8136 3330 8192
rect 2990 8050 3330 8136
rect 2990 7994 3058 8050
rect 3114 7994 3200 8050
rect 3256 7994 3330 8050
rect 2990 7908 3330 7994
rect 2990 7852 3058 7908
rect 3114 7852 3200 7908
rect 3256 7852 3330 7908
rect 2990 7766 3330 7852
rect 2990 7710 3058 7766
rect 3114 7710 3200 7766
rect 3256 7710 3330 7766
rect 2990 7624 3330 7710
rect 2990 7568 3058 7624
rect 3114 7568 3200 7624
rect 3256 7568 3330 7624
rect 2990 7482 3330 7568
rect 2990 7426 3058 7482
rect 3114 7426 3200 7482
rect 3256 7426 3330 7482
rect 2990 7340 3330 7426
rect 2990 7284 3058 7340
rect 3114 7284 3200 7340
rect 3256 7284 3330 7340
rect 2990 7198 3330 7284
rect 2990 7142 3058 7198
rect 3114 7142 3200 7198
rect 3256 7142 3330 7198
rect 2990 7056 3330 7142
rect 2990 7000 3058 7056
rect 3114 7000 3200 7056
rect 3256 7000 3330 7056
rect 2990 6914 3330 7000
rect 2990 6858 3058 6914
rect 3114 6858 3200 6914
rect 3256 6858 3330 6914
rect 2990 6772 3330 6858
rect 2990 6716 3058 6772
rect 3114 6716 3200 6772
rect 3256 6716 3330 6772
rect 2990 6630 3330 6716
rect 2990 6574 3058 6630
rect 3114 6574 3200 6630
rect 3256 6574 3330 6630
rect 2990 6488 3330 6574
rect 2990 6432 3058 6488
rect 3114 6432 3200 6488
rect 3256 6432 3330 6488
rect 2990 6346 3330 6432
rect 2990 6290 3058 6346
rect 3114 6290 3200 6346
rect 3256 6290 3330 6346
rect 2990 6204 3330 6290
rect 2990 6148 3058 6204
rect 3114 6148 3200 6204
rect 3256 6148 3330 6204
rect 2990 6062 3330 6148
rect 2990 6006 3058 6062
rect 3114 6006 3200 6062
rect 3256 6006 3330 6062
rect 2990 5920 3330 6006
rect 2990 5864 3058 5920
rect 3114 5864 3200 5920
rect 3256 5864 3330 5920
rect 2990 5778 3330 5864
rect 2990 5722 3058 5778
rect 3114 5722 3200 5778
rect 3256 5722 3330 5778
rect 2990 5636 3330 5722
rect 2990 5580 3058 5636
rect 3114 5580 3200 5636
rect 3256 5580 3330 5636
rect 2990 5494 3330 5580
rect 2990 5438 3058 5494
rect 3114 5438 3200 5494
rect 3256 5438 3330 5494
rect 2990 5352 3330 5438
rect 2990 5296 3058 5352
rect 3114 5296 3200 5352
rect 3256 5296 3330 5352
rect 2990 5210 3330 5296
rect 2990 5154 3058 5210
rect 3114 5154 3200 5210
rect 3256 5154 3330 5210
rect 2990 5068 3330 5154
rect 2990 5012 3058 5068
rect 3114 5012 3200 5068
rect 3256 5012 3330 5068
rect 2990 4926 3330 5012
rect 2990 4870 3058 4926
rect 3114 4870 3200 4926
rect 3256 4870 3330 4926
rect 2990 4784 3330 4870
rect 2990 4728 3058 4784
rect 3114 4728 3200 4784
rect 3256 4728 3330 4784
rect 2990 4642 3330 4728
rect 2990 4586 3058 4642
rect 3114 4586 3200 4642
rect 3256 4586 3330 4642
rect 2990 4500 3330 4586
rect 2990 4444 3058 4500
rect 3114 4444 3200 4500
rect 3256 4444 3330 4500
rect 2990 4358 3330 4444
rect 2990 4302 3058 4358
rect 3114 4302 3200 4358
rect 3256 4302 3330 4358
rect 2990 4216 3330 4302
rect 2990 4160 3058 4216
rect 3114 4160 3200 4216
rect 3256 4160 3330 4216
rect 2990 4074 3330 4160
rect 2990 4018 3058 4074
rect 3114 4018 3200 4074
rect 3256 4018 3330 4074
rect 2990 3932 3330 4018
rect 2990 3876 3058 3932
rect 3114 3876 3200 3932
rect 3256 3876 3330 3932
rect 2990 3790 3330 3876
rect 2990 3734 3058 3790
rect 3114 3734 3200 3790
rect 3256 3734 3330 3790
rect 2990 3648 3330 3734
rect 2990 3592 3058 3648
rect 3114 3592 3200 3648
rect 3256 3592 3330 3648
rect 2990 3506 3330 3592
rect 2990 3450 3058 3506
rect 3114 3450 3200 3506
rect 3256 3450 3330 3506
rect 2990 3364 3330 3450
rect 2990 3308 3058 3364
rect 3114 3308 3200 3364
rect 3256 3308 3330 3364
rect 2990 3222 3330 3308
rect 2990 3166 3058 3222
rect 3114 3166 3200 3222
rect 3256 3166 3330 3222
rect 2990 3080 3330 3166
rect 2990 3024 3058 3080
rect 3114 3024 3200 3080
rect 3256 3024 3330 3080
rect 2990 2938 3330 3024
rect 2990 2882 3058 2938
rect 3114 2882 3200 2938
rect 3256 2882 3330 2938
rect 2990 2796 3330 2882
rect 2990 2740 3058 2796
rect 3114 2740 3200 2796
rect 3256 2740 3330 2796
rect 2990 2654 3330 2740
rect 2990 2598 3058 2654
rect 3114 2598 3200 2654
rect 3256 2598 3330 2654
rect 2990 2512 3330 2598
rect 2990 2456 3058 2512
rect 3114 2456 3200 2512
rect 3256 2456 3330 2512
rect 2990 2370 3330 2456
rect 2990 2314 3058 2370
rect 3114 2314 3200 2370
rect 3256 2314 3330 2370
rect 2990 2228 3330 2314
rect 2990 2172 3058 2228
rect 3114 2172 3200 2228
rect 3256 2172 3330 2228
rect 2990 2086 3330 2172
rect 2990 2030 3058 2086
rect 3114 2030 3200 2086
rect 3256 2030 3330 2086
rect 2990 1944 3330 2030
rect 2990 1888 3058 1944
rect 3114 1888 3200 1944
rect 3256 1888 3330 1944
rect 2990 1802 3330 1888
rect 2990 1746 3058 1802
rect 3114 1746 3200 1802
rect 3256 1746 3330 1802
rect 2990 1660 3330 1746
rect 2990 1604 3058 1660
rect 3114 1604 3200 1660
rect 3256 1604 3330 1660
rect 2990 1518 3330 1604
rect 2990 1462 3058 1518
rect 3114 1462 3200 1518
rect 3256 1462 3330 1518
rect 2990 1376 3330 1462
rect 2990 1320 3058 1376
rect 3114 1320 3200 1376
rect 3256 1320 3330 1376
rect 2990 1234 3330 1320
rect 2990 1178 3058 1234
rect 3114 1178 3200 1234
rect 3256 1178 3330 1234
rect 2990 1092 3330 1178
rect 2990 1036 3058 1092
rect 3114 1036 3200 1092
rect 3256 1036 3330 1092
rect 2990 950 3330 1036
rect 2990 894 3058 950
rect 3114 894 3200 950
rect 3256 894 3330 950
rect 2990 808 3330 894
rect 2990 752 3058 808
rect 3114 752 3200 808
rect 3256 752 3330 808
rect 2990 666 3330 752
rect 2990 610 3058 666
rect 3114 610 3200 666
rect 3256 610 3330 666
rect 2990 524 3330 610
rect 2990 468 3058 524
rect 3114 468 3200 524
rect 3256 468 3330 524
rect 2990 400 3330 468
rect 3530 12310 3870 12400
rect 3530 12254 3602 12310
rect 3658 12254 3744 12310
rect 3800 12254 3870 12310
rect 3530 12168 3870 12254
rect 3530 12112 3602 12168
rect 3658 12112 3744 12168
rect 3800 12112 3870 12168
rect 3530 12026 3870 12112
rect 3530 11970 3602 12026
rect 3658 11970 3744 12026
rect 3800 11970 3870 12026
rect 3530 11884 3870 11970
rect 3530 11828 3602 11884
rect 3658 11828 3744 11884
rect 3800 11828 3870 11884
rect 3530 11742 3870 11828
rect 3530 11686 3602 11742
rect 3658 11686 3744 11742
rect 3800 11686 3870 11742
rect 3530 11600 3870 11686
rect 3530 11544 3602 11600
rect 3658 11544 3744 11600
rect 3800 11544 3870 11600
rect 3530 11458 3870 11544
rect 3530 11402 3602 11458
rect 3658 11402 3744 11458
rect 3800 11402 3870 11458
rect 3530 11316 3870 11402
rect 3530 11260 3602 11316
rect 3658 11260 3744 11316
rect 3800 11260 3870 11316
rect 3530 11174 3870 11260
rect 3530 11118 3602 11174
rect 3658 11118 3744 11174
rect 3800 11118 3870 11174
rect 3530 11032 3870 11118
rect 3530 10976 3602 11032
rect 3658 10976 3744 11032
rect 3800 10976 3870 11032
rect 3530 10890 3870 10976
rect 3530 10834 3602 10890
rect 3658 10834 3744 10890
rect 3800 10834 3870 10890
rect 3530 10748 3870 10834
rect 3530 10692 3602 10748
rect 3658 10692 3744 10748
rect 3800 10692 3870 10748
rect 3530 10606 3870 10692
rect 3530 10550 3602 10606
rect 3658 10550 3744 10606
rect 3800 10550 3870 10606
rect 3530 10464 3870 10550
rect 3530 10408 3602 10464
rect 3658 10408 3744 10464
rect 3800 10408 3870 10464
rect 3530 10322 3870 10408
rect 3530 10266 3602 10322
rect 3658 10266 3744 10322
rect 3800 10266 3870 10322
rect 3530 10180 3870 10266
rect 3530 10124 3602 10180
rect 3658 10124 3744 10180
rect 3800 10124 3870 10180
rect 3530 10038 3870 10124
rect 3530 9982 3602 10038
rect 3658 9982 3744 10038
rect 3800 9982 3870 10038
rect 3530 9896 3870 9982
rect 3530 9840 3602 9896
rect 3658 9840 3744 9896
rect 3800 9840 3870 9896
rect 3530 9754 3870 9840
rect 3530 9698 3602 9754
rect 3658 9698 3744 9754
rect 3800 9698 3870 9754
rect 3530 9612 3870 9698
rect 3530 9556 3602 9612
rect 3658 9556 3744 9612
rect 3800 9556 3870 9612
rect 3530 9470 3870 9556
rect 3530 9414 3602 9470
rect 3658 9414 3744 9470
rect 3800 9414 3870 9470
rect 3530 9328 3870 9414
rect 3530 9272 3602 9328
rect 3658 9272 3744 9328
rect 3800 9272 3870 9328
rect 3530 9186 3870 9272
rect 3530 9130 3602 9186
rect 3658 9130 3744 9186
rect 3800 9130 3870 9186
rect 3530 9044 3870 9130
rect 3530 8988 3602 9044
rect 3658 8988 3744 9044
rect 3800 8988 3870 9044
rect 3530 8902 3870 8988
rect 3530 8846 3602 8902
rect 3658 8846 3744 8902
rect 3800 8846 3870 8902
rect 3530 8760 3870 8846
rect 3530 8704 3602 8760
rect 3658 8704 3744 8760
rect 3800 8704 3870 8760
rect 3530 8618 3870 8704
rect 3530 8562 3602 8618
rect 3658 8562 3744 8618
rect 3800 8562 3870 8618
rect 3530 8476 3870 8562
rect 3530 8420 3602 8476
rect 3658 8420 3744 8476
rect 3800 8420 3870 8476
rect 3530 8334 3870 8420
rect 3530 8278 3602 8334
rect 3658 8278 3744 8334
rect 3800 8278 3870 8334
rect 3530 8192 3870 8278
rect 3530 8136 3602 8192
rect 3658 8136 3744 8192
rect 3800 8136 3870 8192
rect 3530 8050 3870 8136
rect 3530 7994 3602 8050
rect 3658 7994 3744 8050
rect 3800 7994 3870 8050
rect 3530 7908 3870 7994
rect 3530 7852 3602 7908
rect 3658 7852 3744 7908
rect 3800 7852 3870 7908
rect 3530 7766 3870 7852
rect 3530 7710 3602 7766
rect 3658 7710 3744 7766
rect 3800 7710 3870 7766
rect 3530 7624 3870 7710
rect 3530 7568 3602 7624
rect 3658 7568 3744 7624
rect 3800 7568 3870 7624
rect 3530 7482 3870 7568
rect 3530 7426 3602 7482
rect 3658 7426 3744 7482
rect 3800 7426 3870 7482
rect 3530 7340 3870 7426
rect 3530 7284 3602 7340
rect 3658 7284 3744 7340
rect 3800 7284 3870 7340
rect 3530 7198 3870 7284
rect 3530 7142 3602 7198
rect 3658 7142 3744 7198
rect 3800 7142 3870 7198
rect 3530 7056 3870 7142
rect 3530 7000 3602 7056
rect 3658 7000 3744 7056
rect 3800 7000 3870 7056
rect 3530 6914 3870 7000
rect 3530 6858 3602 6914
rect 3658 6858 3744 6914
rect 3800 6858 3870 6914
rect 3530 6772 3870 6858
rect 3530 6716 3602 6772
rect 3658 6716 3744 6772
rect 3800 6716 3870 6772
rect 3530 6630 3870 6716
rect 3530 6574 3602 6630
rect 3658 6574 3744 6630
rect 3800 6574 3870 6630
rect 3530 6488 3870 6574
rect 3530 6432 3602 6488
rect 3658 6432 3744 6488
rect 3800 6432 3870 6488
rect 3530 6346 3870 6432
rect 3530 6290 3602 6346
rect 3658 6290 3744 6346
rect 3800 6290 3870 6346
rect 3530 6204 3870 6290
rect 3530 6148 3602 6204
rect 3658 6148 3744 6204
rect 3800 6148 3870 6204
rect 3530 6062 3870 6148
rect 3530 6006 3602 6062
rect 3658 6006 3744 6062
rect 3800 6006 3870 6062
rect 3530 5920 3870 6006
rect 3530 5864 3602 5920
rect 3658 5864 3744 5920
rect 3800 5864 3870 5920
rect 3530 5778 3870 5864
rect 3530 5722 3602 5778
rect 3658 5722 3744 5778
rect 3800 5722 3870 5778
rect 3530 5636 3870 5722
rect 3530 5580 3602 5636
rect 3658 5580 3744 5636
rect 3800 5580 3870 5636
rect 3530 5494 3870 5580
rect 3530 5438 3602 5494
rect 3658 5438 3744 5494
rect 3800 5438 3870 5494
rect 3530 5352 3870 5438
rect 3530 5296 3602 5352
rect 3658 5296 3744 5352
rect 3800 5296 3870 5352
rect 3530 5210 3870 5296
rect 3530 5154 3602 5210
rect 3658 5154 3744 5210
rect 3800 5154 3870 5210
rect 3530 5068 3870 5154
rect 3530 5012 3602 5068
rect 3658 5012 3744 5068
rect 3800 5012 3870 5068
rect 3530 4926 3870 5012
rect 3530 4870 3602 4926
rect 3658 4870 3744 4926
rect 3800 4870 3870 4926
rect 3530 4784 3870 4870
rect 3530 4728 3602 4784
rect 3658 4728 3744 4784
rect 3800 4728 3870 4784
rect 3530 4642 3870 4728
rect 3530 4586 3602 4642
rect 3658 4586 3744 4642
rect 3800 4586 3870 4642
rect 3530 4500 3870 4586
rect 3530 4444 3602 4500
rect 3658 4444 3744 4500
rect 3800 4444 3870 4500
rect 3530 4358 3870 4444
rect 3530 4302 3602 4358
rect 3658 4302 3744 4358
rect 3800 4302 3870 4358
rect 3530 4216 3870 4302
rect 3530 4160 3602 4216
rect 3658 4160 3744 4216
rect 3800 4160 3870 4216
rect 3530 4074 3870 4160
rect 3530 4018 3602 4074
rect 3658 4018 3744 4074
rect 3800 4018 3870 4074
rect 3530 3932 3870 4018
rect 3530 3876 3602 3932
rect 3658 3876 3744 3932
rect 3800 3876 3870 3932
rect 3530 3790 3870 3876
rect 3530 3734 3602 3790
rect 3658 3734 3744 3790
rect 3800 3734 3870 3790
rect 3530 3648 3870 3734
rect 3530 3592 3602 3648
rect 3658 3592 3744 3648
rect 3800 3592 3870 3648
rect 3530 3506 3870 3592
rect 3530 3450 3602 3506
rect 3658 3450 3744 3506
rect 3800 3450 3870 3506
rect 3530 3364 3870 3450
rect 3530 3308 3602 3364
rect 3658 3308 3744 3364
rect 3800 3308 3870 3364
rect 3530 3222 3870 3308
rect 3530 3166 3602 3222
rect 3658 3166 3744 3222
rect 3800 3166 3870 3222
rect 3530 3080 3870 3166
rect 3530 3024 3602 3080
rect 3658 3024 3744 3080
rect 3800 3024 3870 3080
rect 3530 2938 3870 3024
rect 3530 2882 3602 2938
rect 3658 2882 3744 2938
rect 3800 2882 3870 2938
rect 3530 2796 3870 2882
rect 3530 2740 3602 2796
rect 3658 2740 3744 2796
rect 3800 2740 3870 2796
rect 3530 2654 3870 2740
rect 3530 2598 3602 2654
rect 3658 2598 3744 2654
rect 3800 2598 3870 2654
rect 3530 2512 3870 2598
rect 3530 2456 3602 2512
rect 3658 2456 3744 2512
rect 3800 2456 3870 2512
rect 3530 2370 3870 2456
rect 3530 2314 3602 2370
rect 3658 2314 3744 2370
rect 3800 2314 3870 2370
rect 3530 2228 3870 2314
rect 3530 2172 3602 2228
rect 3658 2172 3744 2228
rect 3800 2172 3870 2228
rect 3530 2086 3870 2172
rect 3530 2030 3602 2086
rect 3658 2030 3744 2086
rect 3800 2030 3870 2086
rect 3530 1944 3870 2030
rect 3530 1888 3602 1944
rect 3658 1888 3744 1944
rect 3800 1888 3870 1944
rect 3530 1802 3870 1888
rect 3530 1746 3602 1802
rect 3658 1746 3744 1802
rect 3800 1746 3870 1802
rect 3530 1660 3870 1746
rect 3530 1604 3602 1660
rect 3658 1604 3744 1660
rect 3800 1604 3870 1660
rect 3530 1518 3870 1604
rect 3530 1462 3602 1518
rect 3658 1462 3744 1518
rect 3800 1462 3870 1518
rect 3530 1376 3870 1462
rect 3530 1320 3602 1376
rect 3658 1320 3744 1376
rect 3800 1320 3870 1376
rect 3530 1234 3870 1320
rect 3530 1178 3602 1234
rect 3658 1178 3744 1234
rect 3800 1178 3870 1234
rect 3530 1092 3870 1178
rect 3530 1036 3602 1092
rect 3658 1036 3744 1092
rect 3800 1036 3870 1092
rect 3530 950 3870 1036
rect 3530 894 3602 950
rect 3658 894 3744 950
rect 3800 894 3870 950
rect 3530 808 3870 894
rect 3530 752 3602 808
rect 3658 752 3744 808
rect 3800 752 3870 808
rect 3530 666 3870 752
rect 3530 610 3602 666
rect 3658 610 3744 666
rect 3800 610 3870 666
rect 3530 524 3870 610
rect 3530 468 3602 524
rect 3658 468 3744 524
rect 3800 468 3870 524
rect 3530 400 3870 468
rect 4070 12310 4410 12400
rect 4070 12254 4138 12310
rect 4194 12254 4280 12310
rect 4336 12254 4410 12310
rect 4070 12168 4410 12254
rect 4070 12112 4138 12168
rect 4194 12112 4280 12168
rect 4336 12112 4410 12168
rect 4070 12026 4410 12112
rect 4070 11970 4138 12026
rect 4194 11970 4280 12026
rect 4336 11970 4410 12026
rect 4070 11884 4410 11970
rect 4070 11828 4138 11884
rect 4194 11828 4280 11884
rect 4336 11828 4410 11884
rect 4070 11742 4410 11828
rect 4070 11686 4138 11742
rect 4194 11686 4280 11742
rect 4336 11686 4410 11742
rect 4070 11600 4410 11686
rect 4070 11544 4138 11600
rect 4194 11544 4280 11600
rect 4336 11544 4410 11600
rect 4070 11458 4410 11544
rect 4070 11402 4138 11458
rect 4194 11402 4280 11458
rect 4336 11402 4410 11458
rect 4070 11316 4410 11402
rect 4070 11260 4138 11316
rect 4194 11260 4280 11316
rect 4336 11260 4410 11316
rect 4070 11174 4410 11260
rect 4070 11118 4138 11174
rect 4194 11118 4280 11174
rect 4336 11118 4410 11174
rect 4070 11032 4410 11118
rect 4070 10976 4138 11032
rect 4194 10976 4280 11032
rect 4336 10976 4410 11032
rect 4070 10890 4410 10976
rect 4070 10834 4138 10890
rect 4194 10834 4280 10890
rect 4336 10834 4410 10890
rect 4070 10748 4410 10834
rect 4070 10692 4138 10748
rect 4194 10692 4280 10748
rect 4336 10692 4410 10748
rect 4070 10606 4410 10692
rect 4070 10550 4138 10606
rect 4194 10550 4280 10606
rect 4336 10550 4410 10606
rect 4070 10464 4410 10550
rect 4070 10408 4138 10464
rect 4194 10408 4280 10464
rect 4336 10408 4410 10464
rect 4070 10322 4410 10408
rect 4070 10266 4138 10322
rect 4194 10266 4280 10322
rect 4336 10266 4410 10322
rect 4070 10180 4410 10266
rect 4070 10124 4138 10180
rect 4194 10124 4280 10180
rect 4336 10124 4410 10180
rect 4070 10038 4410 10124
rect 4070 9982 4138 10038
rect 4194 9982 4280 10038
rect 4336 9982 4410 10038
rect 4070 9896 4410 9982
rect 4070 9840 4138 9896
rect 4194 9840 4280 9896
rect 4336 9840 4410 9896
rect 4070 9754 4410 9840
rect 4070 9698 4138 9754
rect 4194 9698 4280 9754
rect 4336 9698 4410 9754
rect 4070 9612 4410 9698
rect 4070 9556 4138 9612
rect 4194 9556 4280 9612
rect 4336 9556 4410 9612
rect 4070 9470 4410 9556
rect 4070 9414 4138 9470
rect 4194 9414 4280 9470
rect 4336 9414 4410 9470
rect 4070 9328 4410 9414
rect 4070 9272 4138 9328
rect 4194 9272 4280 9328
rect 4336 9272 4410 9328
rect 4070 9186 4410 9272
rect 4070 9130 4138 9186
rect 4194 9130 4280 9186
rect 4336 9130 4410 9186
rect 4070 9044 4410 9130
rect 4070 8988 4138 9044
rect 4194 8988 4280 9044
rect 4336 8988 4410 9044
rect 4070 8902 4410 8988
rect 4070 8846 4138 8902
rect 4194 8846 4280 8902
rect 4336 8846 4410 8902
rect 4070 8760 4410 8846
rect 4070 8704 4138 8760
rect 4194 8704 4280 8760
rect 4336 8704 4410 8760
rect 4070 8618 4410 8704
rect 4070 8562 4138 8618
rect 4194 8562 4280 8618
rect 4336 8562 4410 8618
rect 4070 8476 4410 8562
rect 4070 8420 4138 8476
rect 4194 8420 4280 8476
rect 4336 8420 4410 8476
rect 4070 8334 4410 8420
rect 4070 8278 4138 8334
rect 4194 8278 4280 8334
rect 4336 8278 4410 8334
rect 4070 8192 4410 8278
rect 4070 8136 4138 8192
rect 4194 8136 4280 8192
rect 4336 8136 4410 8192
rect 4070 8050 4410 8136
rect 4070 7994 4138 8050
rect 4194 7994 4280 8050
rect 4336 7994 4410 8050
rect 4070 7908 4410 7994
rect 4070 7852 4138 7908
rect 4194 7852 4280 7908
rect 4336 7852 4410 7908
rect 4070 7766 4410 7852
rect 4070 7710 4138 7766
rect 4194 7710 4280 7766
rect 4336 7710 4410 7766
rect 4070 7624 4410 7710
rect 4070 7568 4138 7624
rect 4194 7568 4280 7624
rect 4336 7568 4410 7624
rect 4070 7482 4410 7568
rect 4070 7426 4138 7482
rect 4194 7426 4280 7482
rect 4336 7426 4410 7482
rect 4070 7340 4410 7426
rect 4070 7284 4138 7340
rect 4194 7284 4280 7340
rect 4336 7284 4410 7340
rect 4070 7198 4410 7284
rect 4070 7142 4138 7198
rect 4194 7142 4280 7198
rect 4336 7142 4410 7198
rect 4070 7056 4410 7142
rect 4070 7000 4138 7056
rect 4194 7000 4280 7056
rect 4336 7000 4410 7056
rect 4070 6914 4410 7000
rect 4070 6858 4138 6914
rect 4194 6858 4280 6914
rect 4336 6858 4410 6914
rect 4070 6772 4410 6858
rect 4070 6716 4138 6772
rect 4194 6716 4280 6772
rect 4336 6716 4410 6772
rect 4070 6630 4410 6716
rect 4070 6574 4138 6630
rect 4194 6574 4280 6630
rect 4336 6574 4410 6630
rect 4070 6488 4410 6574
rect 4070 6432 4138 6488
rect 4194 6432 4280 6488
rect 4336 6432 4410 6488
rect 4070 6346 4410 6432
rect 4070 6290 4138 6346
rect 4194 6290 4280 6346
rect 4336 6290 4410 6346
rect 4070 6204 4410 6290
rect 4070 6148 4138 6204
rect 4194 6148 4280 6204
rect 4336 6148 4410 6204
rect 4070 6062 4410 6148
rect 4070 6006 4138 6062
rect 4194 6006 4280 6062
rect 4336 6006 4410 6062
rect 4070 5920 4410 6006
rect 4070 5864 4138 5920
rect 4194 5864 4280 5920
rect 4336 5864 4410 5920
rect 4070 5778 4410 5864
rect 4070 5722 4138 5778
rect 4194 5722 4280 5778
rect 4336 5722 4410 5778
rect 4070 5636 4410 5722
rect 4070 5580 4138 5636
rect 4194 5580 4280 5636
rect 4336 5580 4410 5636
rect 4070 5494 4410 5580
rect 4070 5438 4138 5494
rect 4194 5438 4280 5494
rect 4336 5438 4410 5494
rect 4070 5352 4410 5438
rect 4070 5296 4138 5352
rect 4194 5296 4280 5352
rect 4336 5296 4410 5352
rect 4070 5210 4410 5296
rect 4070 5154 4138 5210
rect 4194 5154 4280 5210
rect 4336 5154 4410 5210
rect 4070 5068 4410 5154
rect 4070 5012 4138 5068
rect 4194 5012 4280 5068
rect 4336 5012 4410 5068
rect 4070 4926 4410 5012
rect 4070 4870 4138 4926
rect 4194 4870 4280 4926
rect 4336 4870 4410 4926
rect 4070 4784 4410 4870
rect 4070 4728 4138 4784
rect 4194 4728 4280 4784
rect 4336 4728 4410 4784
rect 4070 4642 4410 4728
rect 4070 4586 4138 4642
rect 4194 4586 4280 4642
rect 4336 4586 4410 4642
rect 4070 4500 4410 4586
rect 4070 4444 4138 4500
rect 4194 4444 4280 4500
rect 4336 4444 4410 4500
rect 4070 4358 4410 4444
rect 4070 4302 4138 4358
rect 4194 4302 4280 4358
rect 4336 4302 4410 4358
rect 4070 4216 4410 4302
rect 4070 4160 4138 4216
rect 4194 4160 4280 4216
rect 4336 4160 4410 4216
rect 4070 4074 4410 4160
rect 4070 4018 4138 4074
rect 4194 4018 4280 4074
rect 4336 4018 4410 4074
rect 4070 3932 4410 4018
rect 4070 3876 4138 3932
rect 4194 3876 4280 3932
rect 4336 3876 4410 3932
rect 4070 3790 4410 3876
rect 4070 3734 4138 3790
rect 4194 3734 4280 3790
rect 4336 3734 4410 3790
rect 4070 3648 4410 3734
rect 4070 3592 4138 3648
rect 4194 3592 4280 3648
rect 4336 3592 4410 3648
rect 4070 3506 4410 3592
rect 4070 3450 4138 3506
rect 4194 3450 4280 3506
rect 4336 3450 4410 3506
rect 4070 3364 4410 3450
rect 4070 3308 4138 3364
rect 4194 3308 4280 3364
rect 4336 3308 4410 3364
rect 4070 3222 4410 3308
rect 4070 3166 4138 3222
rect 4194 3166 4280 3222
rect 4336 3166 4410 3222
rect 4070 3080 4410 3166
rect 4070 3024 4138 3080
rect 4194 3024 4280 3080
rect 4336 3024 4410 3080
rect 4070 2938 4410 3024
rect 4070 2882 4138 2938
rect 4194 2882 4280 2938
rect 4336 2882 4410 2938
rect 4070 2796 4410 2882
rect 4070 2740 4138 2796
rect 4194 2740 4280 2796
rect 4336 2740 4410 2796
rect 4070 2654 4410 2740
rect 4070 2598 4138 2654
rect 4194 2598 4280 2654
rect 4336 2598 4410 2654
rect 4070 2512 4410 2598
rect 4070 2456 4138 2512
rect 4194 2456 4280 2512
rect 4336 2456 4410 2512
rect 4070 2370 4410 2456
rect 4070 2314 4138 2370
rect 4194 2314 4280 2370
rect 4336 2314 4410 2370
rect 4070 2228 4410 2314
rect 4070 2172 4138 2228
rect 4194 2172 4280 2228
rect 4336 2172 4410 2228
rect 4070 2086 4410 2172
rect 4070 2030 4138 2086
rect 4194 2030 4280 2086
rect 4336 2030 4410 2086
rect 4070 1944 4410 2030
rect 4070 1888 4138 1944
rect 4194 1888 4280 1944
rect 4336 1888 4410 1944
rect 4070 1802 4410 1888
rect 4070 1746 4138 1802
rect 4194 1746 4280 1802
rect 4336 1746 4410 1802
rect 4070 1660 4410 1746
rect 4070 1604 4138 1660
rect 4194 1604 4280 1660
rect 4336 1604 4410 1660
rect 4070 1518 4410 1604
rect 4070 1462 4138 1518
rect 4194 1462 4280 1518
rect 4336 1462 4410 1518
rect 4070 1376 4410 1462
rect 4070 1320 4138 1376
rect 4194 1320 4280 1376
rect 4336 1320 4410 1376
rect 4070 1234 4410 1320
rect 4070 1178 4138 1234
rect 4194 1178 4280 1234
rect 4336 1178 4410 1234
rect 4070 1092 4410 1178
rect 4070 1036 4138 1092
rect 4194 1036 4280 1092
rect 4336 1036 4410 1092
rect 4070 950 4410 1036
rect 4070 894 4138 950
rect 4194 894 4280 950
rect 4336 894 4410 950
rect 4070 808 4410 894
rect 4070 752 4138 808
rect 4194 752 4280 808
rect 4336 752 4410 808
rect 4070 666 4410 752
rect 4070 610 4138 666
rect 4194 610 4280 666
rect 4336 610 4410 666
rect 4070 524 4410 610
rect 4070 468 4138 524
rect 4194 468 4280 524
rect 4336 468 4410 524
rect 4070 400 4410 468
rect 4610 12310 4950 12400
rect 4610 12254 4678 12310
rect 4734 12254 4820 12310
rect 4876 12254 4950 12310
rect 4610 12168 4950 12254
rect 4610 12112 4678 12168
rect 4734 12112 4820 12168
rect 4876 12112 4950 12168
rect 4610 12026 4950 12112
rect 4610 11970 4678 12026
rect 4734 11970 4820 12026
rect 4876 11970 4950 12026
rect 4610 11884 4950 11970
rect 4610 11828 4678 11884
rect 4734 11828 4820 11884
rect 4876 11828 4950 11884
rect 4610 11742 4950 11828
rect 4610 11686 4678 11742
rect 4734 11686 4820 11742
rect 4876 11686 4950 11742
rect 4610 11600 4950 11686
rect 4610 11544 4678 11600
rect 4734 11544 4820 11600
rect 4876 11544 4950 11600
rect 4610 11458 4950 11544
rect 4610 11402 4678 11458
rect 4734 11402 4820 11458
rect 4876 11402 4950 11458
rect 4610 11316 4950 11402
rect 4610 11260 4678 11316
rect 4734 11260 4820 11316
rect 4876 11260 4950 11316
rect 4610 11174 4950 11260
rect 4610 11118 4678 11174
rect 4734 11118 4820 11174
rect 4876 11118 4950 11174
rect 4610 11032 4950 11118
rect 4610 10976 4678 11032
rect 4734 10976 4820 11032
rect 4876 10976 4950 11032
rect 4610 10890 4950 10976
rect 4610 10834 4678 10890
rect 4734 10834 4820 10890
rect 4876 10834 4950 10890
rect 4610 10748 4950 10834
rect 4610 10692 4678 10748
rect 4734 10692 4820 10748
rect 4876 10692 4950 10748
rect 4610 10606 4950 10692
rect 4610 10550 4678 10606
rect 4734 10550 4820 10606
rect 4876 10550 4950 10606
rect 4610 10464 4950 10550
rect 4610 10408 4678 10464
rect 4734 10408 4820 10464
rect 4876 10408 4950 10464
rect 4610 10322 4950 10408
rect 4610 10266 4678 10322
rect 4734 10266 4820 10322
rect 4876 10266 4950 10322
rect 4610 10180 4950 10266
rect 4610 10124 4678 10180
rect 4734 10124 4820 10180
rect 4876 10124 4950 10180
rect 4610 10038 4950 10124
rect 4610 9982 4678 10038
rect 4734 9982 4820 10038
rect 4876 9982 4950 10038
rect 4610 9896 4950 9982
rect 4610 9840 4678 9896
rect 4734 9840 4820 9896
rect 4876 9840 4950 9896
rect 4610 9754 4950 9840
rect 4610 9698 4678 9754
rect 4734 9698 4820 9754
rect 4876 9698 4950 9754
rect 4610 9612 4950 9698
rect 4610 9556 4678 9612
rect 4734 9556 4820 9612
rect 4876 9556 4950 9612
rect 4610 9470 4950 9556
rect 4610 9414 4678 9470
rect 4734 9414 4820 9470
rect 4876 9414 4950 9470
rect 4610 9328 4950 9414
rect 4610 9272 4678 9328
rect 4734 9272 4820 9328
rect 4876 9272 4950 9328
rect 4610 9186 4950 9272
rect 4610 9130 4678 9186
rect 4734 9130 4820 9186
rect 4876 9130 4950 9186
rect 4610 9044 4950 9130
rect 4610 8988 4678 9044
rect 4734 8988 4820 9044
rect 4876 8988 4950 9044
rect 4610 8902 4950 8988
rect 4610 8846 4678 8902
rect 4734 8846 4820 8902
rect 4876 8846 4950 8902
rect 4610 8760 4950 8846
rect 4610 8704 4678 8760
rect 4734 8704 4820 8760
rect 4876 8704 4950 8760
rect 4610 8618 4950 8704
rect 4610 8562 4678 8618
rect 4734 8562 4820 8618
rect 4876 8562 4950 8618
rect 4610 8476 4950 8562
rect 4610 8420 4678 8476
rect 4734 8420 4820 8476
rect 4876 8420 4950 8476
rect 4610 8334 4950 8420
rect 4610 8278 4678 8334
rect 4734 8278 4820 8334
rect 4876 8278 4950 8334
rect 4610 8192 4950 8278
rect 4610 8136 4678 8192
rect 4734 8136 4820 8192
rect 4876 8136 4950 8192
rect 4610 8050 4950 8136
rect 4610 7994 4678 8050
rect 4734 7994 4820 8050
rect 4876 7994 4950 8050
rect 4610 7908 4950 7994
rect 4610 7852 4678 7908
rect 4734 7852 4820 7908
rect 4876 7852 4950 7908
rect 4610 7766 4950 7852
rect 4610 7710 4678 7766
rect 4734 7710 4820 7766
rect 4876 7710 4950 7766
rect 4610 7624 4950 7710
rect 4610 7568 4678 7624
rect 4734 7568 4820 7624
rect 4876 7568 4950 7624
rect 4610 7482 4950 7568
rect 4610 7426 4678 7482
rect 4734 7426 4820 7482
rect 4876 7426 4950 7482
rect 4610 7340 4950 7426
rect 4610 7284 4678 7340
rect 4734 7284 4820 7340
rect 4876 7284 4950 7340
rect 4610 7198 4950 7284
rect 4610 7142 4678 7198
rect 4734 7142 4820 7198
rect 4876 7142 4950 7198
rect 4610 7056 4950 7142
rect 4610 7000 4678 7056
rect 4734 7000 4820 7056
rect 4876 7000 4950 7056
rect 4610 6914 4950 7000
rect 4610 6858 4678 6914
rect 4734 6858 4820 6914
rect 4876 6858 4950 6914
rect 4610 6772 4950 6858
rect 4610 6716 4678 6772
rect 4734 6716 4820 6772
rect 4876 6716 4950 6772
rect 4610 6630 4950 6716
rect 4610 6574 4678 6630
rect 4734 6574 4820 6630
rect 4876 6574 4950 6630
rect 4610 6488 4950 6574
rect 4610 6432 4678 6488
rect 4734 6432 4820 6488
rect 4876 6432 4950 6488
rect 4610 6346 4950 6432
rect 4610 6290 4678 6346
rect 4734 6290 4820 6346
rect 4876 6290 4950 6346
rect 4610 6204 4950 6290
rect 4610 6148 4678 6204
rect 4734 6148 4820 6204
rect 4876 6148 4950 6204
rect 4610 6062 4950 6148
rect 4610 6006 4678 6062
rect 4734 6006 4820 6062
rect 4876 6006 4950 6062
rect 4610 5920 4950 6006
rect 4610 5864 4678 5920
rect 4734 5864 4820 5920
rect 4876 5864 4950 5920
rect 4610 5778 4950 5864
rect 4610 5722 4678 5778
rect 4734 5722 4820 5778
rect 4876 5722 4950 5778
rect 4610 5636 4950 5722
rect 4610 5580 4678 5636
rect 4734 5580 4820 5636
rect 4876 5580 4950 5636
rect 4610 5494 4950 5580
rect 4610 5438 4678 5494
rect 4734 5438 4820 5494
rect 4876 5438 4950 5494
rect 4610 5352 4950 5438
rect 4610 5296 4678 5352
rect 4734 5296 4820 5352
rect 4876 5296 4950 5352
rect 4610 5210 4950 5296
rect 4610 5154 4678 5210
rect 4734 5154 4820 5210
rect 4876 5154 4950 5210
rect 4610 5068 4950 5154
rect 4610 5012 4678 5068
rect 4734 5012 4820 5068
rect 4876 5012 4950 5068
rect 4610 4926 4950 5012
rect 4610 4870 4678 4926
rect 4734 4870 4820 4926
rect 4876 4870 4950 4926
rect 4610 4784 4950 4870
rect 4610 4728 4678 4784
rect 4734 4728 4820 4784
rect 4876 4728 4950 4784
rect 4610 4642 4950 4728
rect 4610 4586 4678 4642
rect 4734 4586 4820 4642
rect 4876 4586 4950 4642
rect 4610 4500 4950 4586
rect 4610 4444 4678 4500
rect 4734 4444 4820 4500
rect 4876 4444 4950 4500
rect 4610 4358 4950 4444
rect 4610 4302 4678 4358
rect 4734 4302 4820 4358
rect 4876 4302 4950 4358
rect 4610 4216 4950 4302
rect 4610 4160 4678 4216
rect 4734 4160 4820 4216
rect 4876 4160 4950 4216
rect 4610 4074 4950 4160
rect 4610 4018 4678 4074
rect 4734 4018 4820 4074
rect 4876 4018 4950 4074
rect 4610 3932 4950 4018
rect 4610 3876 4678 3932
rect 4734 3876 4820 3932
rect 4876 3876 4950 3932
rect 4610 3790 4950 3876
rect 4610 3734 4678 3790
rect 4734 3734 4820 3790
rect 4876 3734 4950 3790
rect 4610 3648 4950 3734
rect 4610 3592 4678 3648
rect 4734 3592 4820 3648
rect 4876 3592 4950 3648
rect 4610 3506 4950 3592
rect 4610 3450 4678 3506
rect 4734 3450 4820 3506
rect 4876 3450 4950 3506
rect 4610 3364 4950 3450
rect 4610 3308 4678 3364
rect 4734 3308 4820 3364
rect 4876 3308 4950 3364
rect 4610 3222 4950 3308
rect 4610 3166 4678 3222
rect 4734 3166 4820 3222
rect 4876 3166 4950 3222
rect 4610 3080 4950 3166
rect 4610 3024 4678 3080
rect 4734 3024 4820 3080
rect 4876 3024 4950 3080
rect 4610 2938 4950 3024
rect 4610 2882 4678 2938
rect 4734 2882 4820 2938
rect 4876 2882 4950 2938
rect 4610 2796 4950 2882
rect 4610 2740 4678 2796
rect 4734 2740 4820 2796
rect 4876 2740 4950 2796
rect 4610 2654 4950 2740
rect 4610 2598 4678 2654
rect 4734 2598 4820 2654
rect 4876 2598 4950 2654
rect 4610 2512 4950 2598
rect 4610 2456 4678 2512
rect 4734 2456 4820 2512
rect 4876 2456 4950 2512
rect 4610 2370 4950 2456
rect 4610 2314 4678 2370
rect 4734 2314 4820 2370
rect 4876 2314 4950 2370
rect 4610 2228 4950 2314
rect 4610 2172 4678 2228
rect 4734 2172 4820 2228
rect 4876 2172 4950 2228
rect 4610 2086 4950 2172
rect 4610 2030 4678 2086
rect 4734 2030 4820 2086
rect 4876 2030 4950 2086
rect 4610 1944 4950 2030
rect 4610 1888 4678 1944
rect 4734 1888 4820 1944
rect 4876 1888 4950 1944
rect 4610 1802 4950 1888
rect 4610 1746 4678 1802
rect 4734 1746 4820 1802
rect 4876 1746 4950 1802
rect 4610 1660 4950 1746
rect 4610 1604 4678 1660
rect 4734 1604 4820 1660
rect 4876 1604 4950 1660
rect 4610 1518 4950 1604
rect 4610 1462 4678 1518
rect 4734 1462 4820 1518
rect 4876 1462 4950 1518
rect 4610 1376 4950 1462
rect 4610 1320 4678 1376
rect 4734 1320 4820 1376
rect 4876 1320 4950 1376
rect 4610 1234 4950 1320
rect 4610 1178 4678 1234
rect 4734 1178 4820 1234
rect 4876 1178 4950 1234
rect 4610 1092 4950 1178
rect 4610 1036 4678 1092
rect 4734 1036 4820 1092
rect 4876 1036 4950 1092
rect 4610 950 4950 1036
rect 4610 894 4678 950
rect 4734 894 4820 950
rect 4876 894 4950 950
rect 4610 808 4950 894
rect 4610 752 4678 808
rect 4734 752 4820 808
rect 4876 752 4950 808
rect 4610 666 4950 752
rect 4610 610 4678 666
rect 4734 610 4820 666
rect 4876 610 4950 666
rect 4610 524 4950 610
rect 4610 468 4678 524
rect 4734 468 4820 524
rect 4876 468 4950 524
rect 4610 400 4950 468
rect 5150 12310 5490 12400
rect 5150 12254 5215 12310
rect 5271 12254 5357 12310
rect 5413 12254 5490 12310
rect 5150 12168 5490 12254
rect 5150 12112 5215 12168
rect 5271 12112 5357 12168
rect 5413 12112 5490 12168
rect 5150 12026 5490 12112
rect 5150 11970 5215 12026
rect 5271 11970 5357 12026
rect 5413 11970 5490 12026
rect 5150 11884 5490 11970
rect 5150 11828 5215 11884
rect 5271 11828 5357 11884
rect 5413 11828 5490 11884
rect 5150 11742 5490 11828
rect 5150 11686 5215 11742
rect 5271 11686 5357 11742
rect 5413 11686 5490 11742
rect 5150 11600 5490 11686
rect 5150 11544 5215 11600
rect 5271 11544 5357 11600
rect 5413 11544 5490 11600
rect 5150 11458 5490 11544
rect 5150 11402 5215 11458
rect 5271 11402 5357 11458
rect 5413 11402 5490 11458
rect 5150 11316 5490 11402
rect 5150 11260 5215 11316
rect 5271 11260 5357 11316
rect 5413 11260 5490 11316
rect 5150 11174 5490 11260
rect 5150 11118 5215 11174
rect 5271 11118 5357 11174
rect 5413 11118 5490 11174
rect 5150 11032 5490 11118
rect 5150 10976 5215 11032
rect 5271 10976 5357 11032
rect 5413 10976 5490 11032
rect 5150 10890 5490 10976
rect 5150 10834 5215 10890
rect 5271 10834 5357 10890
rect 5413 10834 5490 10890
rect 5150 10748 5490 10834
rect 5150 10692 5215 10748
rect 5271 10692 5357 10748
rect 5413 10692 5490 10748
rect 5150 10606 5490 10692
rect 5150 10550 5215 10606
rect 5271 10550 5357 10606
rect 5413 10550 5490 10606
rect 5150 10464 5490 10550
rect 5150 10408 5215 10464
rect 5271 10408 5357 10464
rect 5413 10408 5490 10464
rect 5150 10322 5490 10408
rect 5150 10266 5215 10322
rect 5271 10266 5357 10322
rect 5413 10266 5490 10322
rect 5150 10180 5490 10266
rect 5150 10124 5215 10180
rect 5271 10124 5357 10180
rect 5413 10124 5490 10180
rect 5150 10038 5490 10124
rect 5150 9982 5215 10038
rect 5271 9982 5357 10038
rect 5413 9982 5490 10038
rect 5150 9896 5490 9982
rect 5150 9840 5215 9896
rect 5271 9840 5357 9896
rect 5413 9840 5490 9896
rect 5150 9754 5490 9840
rect 5150 9698 5215 9754
rect 5271 9698 5357 9754
rect 5413 9698 5490 9754
rect 5150 9612 5490 9698
rect 5150 9556 5215 9612
rect 5271 9556 5357 9612
rect 5413 9556 5490 9612
rect 5150 9470 5490 9556
rect 5150 9414 5215 9470
rect 5271 9414 5357 9470
rect 5413 9414 5490 9470
rect 5150 9328 5490 9414
rect 5150 9272 5215 9328
rect 5271 9272 5357 9328
rect 5413 9272 5490 9328
rect 5150 9186 5490 9272
rect 5150 9130 5215 9186
rect 5271 9130 5357 9186
rect 5413 9130 5490 9186
rect 5150 9044 5490 9130
rect 5150 8988 5215 9044
rect 5271 8988 5357 9044
rect 5413 8988 5490 9044
rect 5150 8902 5490 8988
rect 5150 8846 5215 8902
rect 5271 8846 5357 8902
rect 5413 8846 5490 8902
rect 5150 8760 5490 8846
rect 5150 8704 5215 8760
rect 5271 8704 5357 8760
rect 5413 8704 5490 8760
rect 5150 8618 5490 8704
rect 5150 8562 5215 8618
rect 5271 8562 5357 8618
rect 5413 8562 5490 8618
rect 5150 8476 5490 8562
rect 5150 8420 5215 8476
rect 5271 8420 5357 8476
rect 5413 8420 5490 8476
rect 5150 8334 5490 8420
rect 5150 8278 5215 8334
rect 5271 8278 5357 8334
rect 5413 8278 5490 8334
rect 5150 8192 5490 8278
rect 5150 8136 5215 8192
rect 5271 8136 5357 8192
rect 5413 8136 5490 8192
rect 5150 8050 5490 8136
rect 5150 7994 5215 8050
rect 5271 7994 5357 8050
rect 5413 7994 5490 8050
rect 5150 7908 5490 7994
rect 5150 7852 5215 7908
rect 5271 7852 5357 7908
rect 5413 7852 5490 7908
rect 5150 7766 5490 7852
rect 5150 7710 5215 7766
rect 5271 7710 5357 7766
rect 5413 7710 5490 7766
rect 5150 7624 5490 7710
rect 5150 7568 5215 7624
rect 5271 7568 5357 7624
rect 5413 7568 5490 7624
rect 5150 7482 5490 7568
rect 5150 7426 5215 7482
rect 5271 7426 5357 7482
rect 5413 7426 5490 7482
rect 5150 7340 5490 7426
rect 5150 7284 5215 7340
rect 5271 7284 5357 7340
rect 5413 7284 5490 7340
rect 5150 7198 5490 7284
rect 5150 7142 5215 7198
rect 5271 7142 5357 7198
rect 5413 7142 5490 7198
rect 5150 7056 5490 7142
rect 5150 7000 5215 7056
rect 5271 7000 5357 7056
rect 5413 7000 5490 7056
rect 5150 6914 5490 7000
rect 5150 6858 5215 6914
rect 5271 6858 5357 6914
rect 5413 6858 5490 6914
rect 5150 6772 5490 6858
rect 5150 6716 5215 6772
rect 5271 6716 5357 6772
rect 5413 6716 5490 6772
rect 5150 6630 5490 6716
rect 5150 6574 5215 6630
rect 5271 6574 5357 6630
rect 5413 6574 5490 6630
rect 5150 6488 5490 6574
rect 5150 6432 5215 6488
rect 5271 6432 5357 6488
rect 5413 6432 5490 6488
rect 5150 6346 5490 6432
rect 5150 6290 5215 6346
rect 5271 6290 5357 6346
rect 5413 6290 5490 6346
rect 5150 6204 5490 6290
rect 5150 6148 5215 6204
rect 5271 6148 5357 6204
rect 5413 6148 5490 6204
rect 5150 6062 5490 6148
rect 5150 6006 5215 6062
rect 5271 6006 5357 6062
rect 5413 6006 5490 6062
rect 5150 5920 5490 6006
rect 5150 5864 5215 5920
rect 5271 5864 5357 5920
rect 5413 5864 5490 5920
rect 5150 5778 5490 5864
rect 5150 5722 5215 5778
rect 5271 5722 5357 5778
rect 5413 5722 5490 5778
rect 5150 5636 5490 5722
rect 5150 5580 5215 5636
rect 5271 5580 5357 5636
rect 5413 5580 5490 5636
rect 5150 5494 5490 5580
rect 5150 5438 5215 5494
rect 5271 5438 5357 5494
rect 5413 5438 5490 5494
rect 5150 5352 5490 5438
rect 5150 5296 5215 5352
rect 5271 5296 5357 5352
rect 5413 5296 5490 5352
rect 5150 5210 5490 5296
rect 5150 5154 5215 5210
rect 5271 5154 5357 5210
rect 5413 5154 5490 5210
rect 5150 5068 5490 5154
rect 5150 5012 5215 5068
rect 5271 5012 5357 5068
rect 5413 5012 5490 5068
rect 5150 4926 5490 5012
rect 5150 4870 5215 4926
rect 5271 4870 5357 4926
rect 5413 4870 5490 4926
rect 5150 4784 5490 4870
rect 5150 4728 5215 4784
rect 5271 4728 5357 4784
rect 5413 4728 5490 4784
rect 5150 4642 5490 4728
rect 5150 4586 5215 4642
rect 5271 4586 5357 4642
rect 5413 4586 5490 4642
rect 5150 4500 5490 4586
rect 5150 4444 5215 4500
rect 5271 4444 5357 4500
rect 5413 4444 5490 4500
rect 5150 4358 5490 4444
rect 5150 4302 5215 4358
rect 5271 4302 5357 4358
rect 5413 4302 5490 4358
rect 5150 4216 5490 4302
rect 5150 4160 5215 4216
rect 5271 4160 5357 4216
rect 5413 4160 5490 4216
rect 5150 4074 5490 4160
rect 5150 4018 5215 4074
rect 5271 4018 5357 4074
rect 5413 4018 5490 4074
rect 5150 3932 5490 4018
rect 5150 3876 5215 3932
rect 5271 3876 5357 3932
rect 5413 3876 5490 3932
rect 5150 3790 5490 3876
rect 5150 3734 5215 3790
rect 5271 3734 5357 3790
rect 5413 3734 5490 3790
rect 5150 3648 5490 3734
rect 5150 3592 5215 3648
rect 5271 3592 5357 3648
rect 5413 3592 5490 3648
rect 5150 3506 5490 3592
rect 5150 3450 5215 3506
rect 5271 3450 5357 3506
rect 5413 3450 5490 3506
rect 5150 3364 5490 3450
rect 5150 3308 5215 3364
rect 5271 3308 5357 3364
rect 5413 3308 5490 3364
rect 5150 3222 5490 3308
rect 5150 3166 5215 3222
rect 5271 3166 5357 3222
rect 5413 3166 5490 3222
rect 5150 3080 5490 3166
rect 5150 3024 5215 3080
rect 5271 3024 5357 3080
rect 5413 3024 5490 3080
rect 5150 2938 5490 3024
rect 5150 2882 5215 2938
rect 5271 2882 5357 2938
rect 5413 2882 5490 2938
rect 5150 2796 5490 2882
rect 5150 2740 5215 2796
rect 5271 2740 5357 2796
rect 5413 2740 5490 2796
rect 5150 2654 5490 2740
rect 5150 2598 5215 2654
rect 5271 2598 5357 2654
rect 5413 2598 5490 2654
rect 5150 2512 5490 2598
rect 5150 2456 5215 2512
rect 5271 2456 5357 2512
rect 5413 2456 5490 2512
rect 5150 2370 5490 2456
rect 5150 2314 5215 2370
rect 5271 2314 5357 2370
rect 5413 2314 5490 2370
rect 5150 2228 5490 2314
rect 5150 2172 5215 2228
rect 5271 2172 5357 2228
rect 5413 2172 5490 2228
rect 5150 2086 5490 2172
rect 5150 2030 5215 2086
rect 5271 2030 5357 2086
rect 5413 2030 5490 2086
rect 5150 1944 5490 2030
rect 5150 1888 5215 1944
rect 5271 1888 5357 1944
rect 5413 1888 5490 1944
rect 5150 1802 5490 1888
rect 5150 1746 5215 1802
rect 5271 1746 5357 1802
rect 5413 1746 5490 1802
rect 5150 1660 5490 1746
rect 5150 1604 5215 1660
rect 5271 1604 5357 1660
rect 5413 1604 5490 1660
rect 5150 1518 5490 1604
rect 5150 1462 5215 1518
rect 5271 1462 5357 1518
rect 5413 1462 5490 1518
rect 5150 1376 5490 1462
rect 5150 1320 5215 1376
rect 5271 1320 5357 1376
rect 5413 1320 5490 1376
rect 5150 1234 5490 1320
rect 5150 1178 5215 1234
rect 5271 1178 5357 1234
rect 5413 1178 5490 1234
rect 5150 1092 5490 1178
rect 5150 1036 5215 1092
rect 5271 1036 5357 1092
rect 5413 1036 5490 1092
rect 5150 950 5490 1036
rect 5150 894 5215 950
rect 5271 894 5357 950
rect 5413 894 5490 950
rect 5150 808 5490 894
rect 5150 752 5215 808
rect 5271 752 5357 808
rect 5413 752 5490 808
rect 5150 666 5490 752
rect 5150 610 5215 666
rect 5271 610 5357 666
rect 5413 610 5490 666
rect 5150 524 5490 610
rect 5150 468 5215 524
rect 5271 468 5357 524
rect 5413 468 5490 524
rect 5150 400 5490 468
rect 5690 12310 6030 12400
rect 5690 12254 5760 12310
rect 5816 12254 5902 12310
rect 5958 12254 6030 12310
rect 5690 12168 6030 12254
rect 5690 12112 5760 12168
rect 5816 12112 5902 12168
rect 5958 12112 6030 12168
rect 5690 12026 6030 12112
rect 5690 11970 5760 12026
rect 5816 11970 5902 12026
rect 5958 11970 6030 12026
rect 5690 11884 6030 11970
rect 5690 11828 5760 11884
rect 5816 11828 5902 11884
rect 5958 11828 6030 11884
rect 5690 11742 6030 11828
rect 5690 11686 5760 11742
rect 5816 11686 5902 11742
rect 5958 11686 6030 11742
rect 5690 11600 6030 11686
rect 5690 11544 5760 11600
rect 5816 11544 5902 11600
rect 5958 11544 6030 11600
rect 5690 11458 6030 11544
rect 5690 11402 5760 11458
rect 5816 11402 5902 11458
rect 5958 11402 6030 11458
rect 5690 11316 6030 11402
rect 5690 11260 5760 11316
rect 5816 11260 5902 11316
rect 5958 11260 6030 11316
rect 5690 11174 6030 11260
rect 5690 11118 5760 11174
rect 5816 11118 5902 11174
rect 5958 11118 6030 11174
rect 5690 11032 6030 11118
rect 5690 10976 5760 11032
rect 5816 10976 5902 11032
rect 5958 10976 6030 11032
rect 5690 10890 6030 10976
rect 5690 10834 5760 10890
rect 5816 10834 5902 10890
rect 5958 10834 6030 10890
rect 5690 10748 6030 10834
rect 5690 10692 5760 10748
rect 5816 10692 5902 10748
rect 5958 10692 6030 10748
rect 5690 10606 6030 10692
rect 5690 10550 5760 10606
rect 5816 10550 5902 10606
rect 5958 10550 6030 10606
rect 5690 10464 6030 10550
rect 5690 10408 5760 10464
rect 5816 10408 5902 10464
rect 5958 10408 6030 10464
rect 5690 10322 6030 10408
rect 5690 10266 5760 10322
rect 5816 10266 5902 10322
rect 5958 10266 6030 10322
rect 5690 10180 6030 10266
rect 5690 10124 5760 10180
rect 5816 10124 5902 10180
rect 5958 10124 6030 10180
rect 5690 10038 6030 10124
rect 5690 9982 5760 10038
rect 5816 9982 5902 10038
rect 5958 9982 6030 10038
rect 5690 9896 6030 9982
rect 5690 9840 5760 9896
rect 5816 9840 5902 9896
rect 5958 9840 6030 9896
rect 5690 9754 6030 9840
rect 5690 9698 5760 9754
rect 5816 9698 5902 9754
rect 5958 9698 6030 9754
rect 5690 9612 6030 9698
rect 5690 9556 5760 9612
rect 5816 9556 5902 9612
rect 5958 9556 6030 9612
rect 5690 9470 6030 9556
rect 5690 9414 5760 9470
rect 5816 9414 5902 9470
rect 5958 9414 6030 9470
rect 5690 9328 6030 9414
rect 5690 9272 5760 9328
rect 5816 9272 5902 9328
rect 5958 9272 6030 9328
rect 5690 9186 6030 9272
rect 5690 9130 5760 9186
rect 5816 9130 5902 9186
rect 5958 9130 6030 9186
rect 5690 9044 6030 9130
rect 5690 8988 5760 9044
rect 5816 8988 5902 9044
rect 5958 8988 6030 9044
rect 5690 8902 6030 8988
rect 5690 8846 5760 8902
rect 5816 8846 5902 8902
rect 5958 8846 6030 8902
rect 5690 8760 6030 8846
rect 5690 8704 5760 8760
rect 5816 8704 5902 8760
rect 5958 8704 6030 8760
rect 5690 8618 6030 8704
rect 5690 8562 5760 8618
rect 5816 8562 5902 8618
rect 5958 8562 6030 8618
rect 5690 8476 6030 8562
rect 5690 8420 5760 8476
rect 5816 8420 5902 8476
rect 5958 8420 6030 8476
rect 5690 8334 6030 8420
rect 5690 8278 5760 8334
rect 5816 8278 5902 8334
rect 5958 8278 6030 8334
rect 5690 8192 6030 8278
rect 5690 8136 5760 8192
rect 5816 8136 5902 8192
rect 5958 8136 6030 8192
rect 5690 8050 6030 8136
rect 5690 7994 5760 8050
rect 5816 7994 5902 8050
rect 5958 7994 6030 8050
rect 5690 7908 6030 7994
rect 5690 7852 5760 7908
rect 5816 7852 5902 7908
rect 5958 7852 6030 7908
rect 5690 7766 6030 7852
rect 5690 7710 5760 7766
rect 5816 7710 5902 7766
rect 5958 7710 6030 7766
rect 5690 7624 6030 7710
rect 5690 7568 5760 7624
rect 5816 7568 5902 7624
rect 5958 7568 6030 7624
rect 5690 7482 6030 7568
rect 5690 7426 5760 7482
rect 5816 7426 5902 7482
rect 5958 7426 6030 7482
rect 5690 7340 6030 7426
rect 5690 7284 5760 7340
rect 5816 7284 5902 7340
rect 5958 7284 6030 7340
rect 5690 7198 6030 7284
rect 5690 7142 5760 7198
rect 5816 7142 5902 7198
rect 5958 7142 6030 7198
rect 5690 7056 6030 7142
rect 5690 7000 5760 7056
rect 5816 7000 5902 7056
rect 5958 7000 6030 7056
rect 5690 6914 6030 7000
rect 5690 6858 5760 6914
rect 5816 6858 5902 6914
rect 5958 6858 6030 6914
rect 5690 6772 6030 6858
rect 5690 6716 5760 6772
rect 5816 6716 5902 6772
rect 5958 6716 6030 6772
rect 5690 6630 6030 6716
rect 5690 6574 5760 6630
rect 5816 6574 5902 6630
rect 5958 6574 6030 6630
rect 5690 6488 6030 6574
rect 5690 6432 5760 6488
rect 5816 6432 5902 6488
rect 5958 6432 6030 6488
rect 5690 6346 6030 6432
rect 5690 6290 5760 6346
rect 5816 6290 5902 6346
rect 5958 6290 6030 6346
rect 5690 6204 6030 6290
rect 5690 6148 5760 6204
rect 5816 6148 5902 6204
rect 5958 6148 6030 6204
rect 5690 6062 6030 6148
rect 5690 6006 5760 6062
rect 5816 6006 5902 6062
rect 5958 6006 6030 6062
rect 5690 5920 6030 6006
rect 5690 5864 5760 5920
rect 5816 5864 5902 5920
rect 5958 5864 6030 5920
rect 5690 5778 6030 5864
rect 5690 5722 5760 5778
rect 5816 5722 5902 5778
rect 5958 5722 6030 5778
rect 5690 5636 6030 5722
rect 5690 5580 5760 5636
rect 5816 5580 5902 5636
rect 5958 5580 6030 5636
rect 5690 5494 6030 5580
rect 5690 5438 5760 5494
rect 5816 5438 5902 5494
rect 5958 5438 6030 5494
rect 5690 5352 6030 5438
rect 5690 5296 5760 5352
rect 5816 5296 5902 5352
rect 5958 5296 6030 5352
rect 5690 5210 6030 5296
rect 5690 5154 5760 5210
rect 5816 5154 5902 5210
rect 5958 5154 6030 5210
rect 5690 5068 6030 5154
rect 5690 5012 5760 5068
rect 5816 5012 5902 5068
rect 5958 5012 6030 5068
rect 5690 4926 6030 5012
rect 5690 4870 5760 4926
rect 5816 4870 5902 4926
rect 5958 4870 6030 4926
rect 5690 4784 6030 4870
rect 5690 4728 5760 4784
rect 5816 4728 5902 4784
rect 5958 4728 6030 4784
rect 5690 4642 6030 4728
rect 5690 4586 5760 4642
rect 5816 4586 5902 4642
rect 5958 4586 6030 4642
rect 5690 4500 6030 4586
rect 5690 4444 5760 4500
rect 5816 4444 5902 4500
rect 5958 4444 6030 4500
rect 5690 4358 6030 4444
rect 5690 4302 5760 4358
rect 5816 4302 5902 4358
rect 5958 4302 6030 4358
rect 5690 4216 6030 4302
rect 5690 4160 5760 4216
rect 5816 4160 5902 4216
rect 5958 4160 6030 4216
rect 5690 4074 6030 4160
rect 5690 4018 5760 4074
rect 5816 4018 5902 4074
rect 5958 4018 6030 4074
rect 5690 3932 6030 4018
rect 5690 3876 5760 3932
rect 5816 3876 5902 3932
rect 5958 3876 6030 3932
rect 5690 3790 6030 3876
rect 5690 3734 5760 3790
rect 5816 3734 5902 3790
rect 5958 3734 6030 3790
rect 5690 3648 6030 3734
rect 5690 3592 5760 3648
rect 5816 3592 5902 3648
rect 5958 3592 6030 3648
rect 5690 3506 6030 3592
rect 5690 3450 5760 3506
rect 5816 3450 5902 3506
rect 5958 3450 6030 3506
rect 5690 3364 6030 3450
rect 5690 3308 5760 3364
rect 5816 3308 5902 3364
rect 5958 3308 6030 3364
rect 5690 3222 6030 3308
rect 5690 3166 5760 3222
rect 5816 3166 5902 3222
rect 5958 3166 6030 3222
rect 5690 3080 6030 3166
rect 5690 3024 5760 3080
rect 5816 3024 5902 3080
rect 5958 3024 6030 3080
rect 5690 2938 6030 3024
rect 5690 2882 5760 2938
rect 5816 2882 5902 2938
rect 5958 2882 6030 2938
rect 5690 2796 6030 2882
rect 5690 2740 5760 2796
rect 5816 2740 5902 2796
rect 5958 2740 6030 2796
rect 5690 2654 6030 2740
rect 5690 2598 5760 2654
rect 5816 2598 5902 2654
rect 5958 2598 6030 2654
rect 5690 2512 6030 2598
rect 5690 2456 5760 2512
rect 5816 2456 5902 2512
rect 5958 2456 6030 2512
rect 5690 2370 6030 2456
rect 5690 2314 5760 2370
rect 5816 2314 5902 2370
rect 5958 2314 6030 2370
rect 5690 2228 6030 2314
rect 5690 2172 5760 2228
rect 5816 2172 5902 2228
rect 5958 2172 6030 2228
rect 5690 2086 6030 2172
rect 5690 2030 5760 2086
rect 5816 2030 5902 2086
rect 5958 2030 6030 2086
rect 5690 1944 6030 2030
rect 5690 1888 5760 1944
rect 5816 1888 5902 1944
rect 5958 1888 6030 1944
rect 5690 1802 6030 1888
rect 5690 1746 5760 1802
rect 5816 1746 5902 1802
rect 5958 1746 6030 1802
rect 5690 1660 6030 1746
rect 5690 1604 5760 1660
rect 5816 1604 5902 1660
rect 5958 1604 6030 1660
rect 5690 1518 6030 1604
rect 5690 1462 5760 1518
rect 5816 1462 5902 1518
rect 5958 1462 6030 1518
rect 5690 1376 6030 1462
rect 5690 1320 5760 1376
rect 5816 1320 5902 1376
rect 5958 1320 6030 1376
rect 5690 1234 6030 1320
rect 5690 1178 5760 1234
rect 5816 1178 5902 1234
rect 5958 1178 6030 1234
rect 5690 1092 6030 1178
rect 5690 1036 5760 1092
rect 5816 1036 5902 1092
rect 5958 1036 6030 1092
rect 5690 950 6030 1036
rect 5690 894 5760 950
rect 5816 894 5902 950
rect 5958 894 6030 950
rect 5690 808 6030 894
rect 5690 752 5760 808
rect 5816 752 5902 808
rect 5958 752 6030 808
rect 5690 666 6030 752
rect 5690 610 5760 666
rect 5816 610 5902 666
rect 5958 610 6030 666
rect 5690 524 6030 610
rect 5690 468 5760 524
rect 5816 468 5902 524
rect 5958 468 6030 524
rect 5690 400 6030 468
rect 6230 12310 6570 12400
rect 6230 12254 6300 12310
rect 6356 12254 6442 12310
rect 6498 12254 6570 12310
rect 6230 12168 6570 12254
rect 6230 12112 6300 12168
rect 6356 12112 6442 12168
rect 6498 12112 6570 12168
rect 6230 12026 6570 12112
rect 6230 11970 6300 12026
rect 6356 11970 6442 12026
rect 6498 11970 6570 12026
rect 6230 11884 6570 11970
rect 6230 11828 6300 11884
rect 6356 11828 6442 11884
rect 6498 11828 6570 11884
rect 6230 11742 6570 11828
rect 6230 11686 6300 11742
rect 6356 11686 6442 11742
rect 6498 11686 6570 11742
rect 6230 11600 6570 11686
rect 6230 11544 6300 11600
rect 6356 11544 6442 11600
rect 6498 11544 6570 11600
rect 6230 11458 6570 11544
rect 6230 11402 6300 11458
rect 6356 11402 6442 11458
rect 6498 11402 6570 11458
rect 6230 11316 6570 11402
rect 6230 11260 6300 11316
rect 6356 11260 6442 11316
rect 6498 11260 6570 11316
rect 6230 11174 6570 11260
rect 6230 11118 6300 11174
rect 6356 11118 6442 11174
rect 6498 11118 6570 11174
rect 6230 11032 6570 11118
rect 6230 10976 6300 11032
rect 6356 10976 6442 11032
rect 6498 10976 6570 11032
rect 6230 10890 6570 10976
rect 6230 10834 6300 10890
rect 6356 10834 6442 10890
rect 6498 10834 6570 10890
rect 6230 10748 6570 10834
rect 6230 10692 6300 10748
rect 6356 10692 6442 10748
rect 6498 10692 6570 10748
rect 6230 10606 6570 10692
rect 6230 10550 6300 10606
rect 6356 10550 6442 10606
rect 6498 10550 6570 10606
rect 6230 10464 6570 10550
rect 6230 10408 6300 10464
rect 6356 10408 6442 10464
rect 6498 10408 6570 10464
rect 6230 10322 6570 10408
rect 6230 10266 6300 10322
rect 6356 10266 6442 10322
rect 6498 10266 6570 10322
rect 6230 10180 6570 10266
rect 6230 10124 6300 10180
rect 6356 10124 6442 10180
rect 6498 10124 6570 10180
rect 6230 10038 6570 10124
rect 6230 9982 6300 10038
rect 6356 9982 6442 10038
rect 6498 9982 6570 10038
rect 6230 9896 6570 9982
rect 6230 9840 6300 9896
rect 6356 9840 6442 9896
rect 6498 9840 6570 9896
rect 6230 9754 6570 9840
rect 6230 9698 6300 9754
rect 6356 9698 6442 9754
rect 6498 9698 6570 9754
rect 6230 9612 6570 9698
rect 6230 9556 6300 9612
rect 6356 9556 6442 9612
rect 6498 9556 6570 9612
rect 6230 9470 6570 9556
rect 6230 9414 6300 9470
rect 6356 9414 6442 9470
rect 6498 9414 6570 9470
rect 6230 9328 6570 9414
rect 6230 9272 6300 9328
rect 6356 9272 6442 9328
rect 6498 9272 6570 9328
rect 6230 9186 6570 9272
rect 6230 9130 6300 9186
rect 6356 9130 6442 9186
rect 6498 9130 6570 9186
rect 6230 9044 6570 9130
rect 6230 8988 6300 9044
rect 6356 8988 6442 9044
rect 6498 8988 6570 9044
rect 6230 8902 6570 8988
rect 6230 8846 6300 8902
rect 6356 8846 6442 8902
rect 6498 8846 6570 8902
rect 6230 8760 6570 8846
rect 6230 8704 6300 8760
rect 6356 8704 6442 8760
rect 6498 8704 6570 8760
rect 6230 8618 6570 8704
rect 6230 8562 6300 8618
rect 6356 8562 6442 8618
rect 6498 8562 6570 8618
rect 6230 8476 6570 8562
rect 6230 8420 6300 8476
rect 6356 8420 6442 8476
rect 6498 8420 6570 8476
rect 6230 8334 6570 8420
rect 6230 8278 6300 8334
rect 6356 8278 6442 8334
rect 6498 8278 6570 8334
rect 6230 8192 6570 8278
rect 6230 8136 6300 8192
rect 6356 8136 6442 8192
rect 6498 8136 6570 8192
rect 6230 8050 6570 8136
rect 6230 7994 6300 8050
rect 6356 7994 6442 8050
rect 6498 7994 6570 8050
rect 6230 7908 6570 7994
rect 6230 7852 6300 7908
rect 6356 7852 6442 7908
rect 6498 7852 6570 7908
rect 6230 7766 6570 7852
rect 6230 7710 6300 7766
rect 6356 7710 6442 7766
rect 6498 7710 6570 7766
rect 6230 7624 6570 7710
rect 6230 7568 6300 7624
rect 6356 7568 6442 7624
rect 6498 7568 6570 7624
rect 6230 7482 6570 7568
rect 6230 7426 6300 7482
rect 6356 7426 6442 7482
rect 6498 7426 6570 7482
rect 6230 7340 6570 7426
rect 6230 7284 6300 7340
rect 6356 7284 6442 7340
rect 6498 7284 6570 7340
rect 6230 7198 6570 7284
rect 6230 7142 6300 7198
rect 6356 7142 6442 7198
rect 6498 7142 6570 7198
rect 6230 7056 6570 7142
rect 6230 7000 6300 7056
rect 6356 7000 6442 7056
rect 6498 7000 6570 7056
rect 6230 6914 6570 7000
rect 6230 6858 6300 6914
rect 6356 6858 6442 6914
rect 6498 6858 6570 6914
rect 6230 6772 6570 6858
rect 6230 6716 6300 6772
rect 6356 6716 6442 6772
rect 6498 6716 6570 6772
rect 6230 6630 6570 6716
rect 6230 6574 6300 6630
rect 6356 6574 6442 6630
rect 6498 6574 6570 6630
rect 6230 6488 6570 6574
rect 6230 6432 6300 6488
rect 6356 6432 6442 6488
rect 6498 6432 6570 6488
rect 6230 6346 6570 6432
rect 6230 6290 6300 6346
rect 6356 6290 6442 6346
rect 6498 6290 6570 6346
rect 6230 6204 6570 6290
rect 6230 6148 6300 6204
rect 6356 6148 6442 6204
rect 6498 6148 6570 6204
rect 6230 6062 6570 6148
rect 6230 6006 6300 6062
rect 6356 6006 6442 6062
rect 6498 6006 6570 6062
rect 6230 5920 6570 6006
rect 6230 5864 6300 5920
rect 6356 5864 6442 5920
rect 6498 5864 6570 5920
rect 6230 5778 6570 5864
rect 6230 5722 6300 5778
rect 6356 5722 6442 5778
rect 6498 5722 6570 5778
rect 6230 5636 6570 5722
rect 6230 5580 6300 5636
rect 6356 5580 6442 5636
rect 6498 5580 6570 5636
rect 6230 5494 6570 5580
rect 6230 5438 6300 5494
rect 6356 5438 6442 5494
rect 6498 5438 6570 5494
rect 6230 5352 6570 5438
rect 6230 5296 6300 5352
rect 6356 5296 6442 5352
rect 6498 5296 6570 5352
rect 6230 5210 6570 5296
rect 6230 5154 6300 5210
rect 6356 5154 6442 5210
rect 6498 5154 6570 5210
rect 6230 5068 6570 5154
rect 6230 5012 6300 5068
rect 6356 5012 6442 5068
rect 6498 5012 6570 5068
rect 6230 4926 6570 5012
rect 6230 4870 6300 4926
rect 6356 4870 6442 4926
rect 6498 4870 6570 4926
rect 6230 4784 6570 4870
rect 6230 4728 6300 4784
rect 6356 4728 6442 4784
rect 6498 4728 6570 4784
rect 6230 4642 6570 4728
rect 6230 4586 6300 4642
rect 6356 4586 6442 4642
rect 6498 4586 6570 4642
rect 6230 4500 6570 4586
rect 6230 4444 6300 4500
rect 6356 4444 6442 4500
rect 6498 4444 6570 4500
rect 6230 4358 6570 4444
rect 6230 4302 6300 4358
rect 6356 4302 6442 4358
rect 6498 4302 6570 4358
rect 6230 4216 6570 4302
rect 6230 4160 6300 4216
rect 6356 4160 6442 4216
rect 6498 4160 6570 4216
rect 6230 4074 6570 4160
rect 6230 4018 6300 4074
rect 6356 4018 6442 4074
rect 6498 4018 6570 4074
rect 6230 3932 6570 4018
rect 6230 3876 6300 3932
rect 6356 3876 6442 3932
rect 6498 3876 6570 3932
rect 6230 3790 6570 3876
rect 6230 3734 6300 3790
rect 6356 3734 6442 3790
rect 6498 3734 6570 3790
rect 6230 3648 6570 3734
rect 6230 3592 6300 3648
rect 6356 3592 6442 3648
rect 6498 3592 6570 3648
rect 6230 3506 6570 3592
rect 6230 3450 6300 3506
rect 6356 3450 6442 3506
rect 6498 3450 6570 3506
rect 6230 3364 6570 3450
rect 6230 3308 6300 3364
rect 6356 3308 6442 3364
rect 6498 3308 6570 3364
rect 6230 3222 6570 3308
rect 6230 3166 6300 3222
rect 6356 3166 6442 3222
rect 6498 3166 6570 3222
rect 6230 3080 6570 3166
rect 6230 3024 6300 3080
rect 6356 3024 6442 3080
rect 6498 3024 6570 3080
rect 6230 2938 6570 3024
rect 6230 2882 6300 2938
rect 6356 2882 6442 2938
rect 6498 2882 6570 2938
rect 6230 2796 6570 2882
rect 6230 2740 6300 2796
rect 6356 2740 6442 2796
rect 6498 2740 6570 2796
rect 6230 2654 6570 2740
rect 6230 2598 6300 2654
rect 6356 2598 6442 2654
rect 6498 2598 6570 2654
rect 6230 2512 6570 2598
rect 6230 2456 6300 2512
rect 6356 2456 6442 2512
rect 6498 2456 6570 2512
rect 6230 2370 6570 2456
rect 6230 2314 6300 2370
rect 6356 2314 6442 2370
rect 6498 2314 6570 2370
rect 6230 2228 6570 2314
rect 6230 2172 6300 2228
rect 6356 2172 6442 2228
rect 6498 2172 6570 2228
rect 6230 2086 6570 2172
rect 6230 2030 6300 2086
rect 6356 2030 6442 2086
rect 6498 2030 6570 2086
rect 6230 1944 6570 2030
rect 6230 1888 6300 1944
rect 6356 1888 6442 1944
rect 6498 1888 6570 1944
rect 6230 1802 6570 1888
rect 6230 1746 6300 1802
rect 6356 1746 6442 1802
rect 6498 1746 6570 1802
rect 6230 1660 6570 1746
rect 6230 1604 6300 1660
rect 6356 1604 6442 1660
rect 6498 1604 6570 1660
rect 6230 1518 6570 1604
rect 6230 1462 6300 1518
rect 6356 1462 6442 1518
rect 6498 1462 6570 1518
rect 6230 1376 6570 1462
rect 6230 1320 6300 1376
rect 6356 1320 6442 1376
rect 6498 1320 6570 1376
rect 6230 1234 6570 1320
rect 6230 1178 6300 1234
rect 6356 1178 6442 1234
rect 6498 1178 6570 1234
rect 6230 1092 6570 1178
rect 6230 1036 6300 1092
rect 6356 1036 6442 1092
rect 6498 1036 6570 1092
rect 6230 950 6570 1036
rect 6230 894 6300 950
rect 6356 894 6442 950
rect 6498 894 6570 950
rect 6230 808 6570 894
rect 6230 752 6300 808
rect 6356 752 6442 808
rect 6498 752 6570 808
rect 6230 666 6570 752
rect 6230 610 6300 666
rect 6356 610 6442 666
rect 6498 610 6570 666
rect 6230 524 6570 610
rect 6230 468 6300 524
rect 6356 468 6442 524
rect 6498 468 6570 524
rect 6230 400 6570 468
rect 6770 12310 7110 12400
rect 6770 12254 6845 12310
rect 6901 12254 6987 12310
rect 7043 12254 7110 12310
rect 6770 12168 7110 12254
rect 6770 12112 6845 12168
rect 6901 12112 6987 12168
rect 7043 12112 7110 12168
rect 6770 12026 7110 12112
rect 6770 11970 6845 12026
rect 6901 11970 6987 12026
rect 7043 11970 7110 12026
rect 6770 11884 7110 11970
rect 6770 11828 6845 11884
rect 6901 11828 6987 11884
rect 7043 11828 7110 11884
rect 6770 11742 7110 11828
rect 6770 11686 6845 11742
rect 6901 11686 6987 11742
rect 7043 11686 7110 11742
rect 6770 11600 7110 11686
rect 6770 11544 6845 11600
rect 6901 11544 6987 11600
rect 7043 11544 7110 11600
rect 6770 11458 7110 11544
rect 6770 11402 6845 11458
rect 6901 11402 6987 11458
rect 7043 11402 7110 11458
rect 6770 11316 7110 11402
rect 6770 11260 6845 11316
rect 6901 11260 6987 11316
rect 7043 11260 7110 11316
rect 6770 11174 7110 11260
rect 6770 11118 6845 11174
rect 6901 11118 6987 11174
rect 7043 11118 7110 11174
rect 6770 11032 7110 11118
rect 6770 10976 6845 11032
rect 6901 10976 6987 11032
rect 7043 10976 7110 11032
rect 6770 10890 7110 10976
rect 6770 10834 6845 10890
rect 6901 10834 6987 10890
rect 7043 10834 7110 10890
rect 6770 10748 7110 10834
rect 6770 10692 6845 10748
rect 6901 10692 6987 10748
rect 7043 10692 7110 10748
rect 6770 10606 7110 10692
rect 6770 10550 6845 10606
rect 6901 10550 6987 10606
rect 7043 10550 7110 10606
rect 6770 10464 7110 10550
rect 6770 10408 6845 10464
rect 6901 10408 6987 10464
rect 7043 10408 7110 10464
rect 6770 10322 7110 10408
rect 6770 10266 6845 10322
rect 6901 10266 6987 10322
rect 7043 10266 7110 10322
rect 6770 10180 7110 10266
rect 6770 10124 6845 10180
rect 6901 10124 6987 10180
rect 7043 10124 7110 10180
rect 6770 10038 7110 10124
rect 6770 9982 6845 10038
rect 6901 9982 6987 10038
rect 7043 9982 7110 10038
rect 6770 9896 7110 9982
rect 6770 9840 6845 9896
rect 6901 9840 6987 9896
rect 7043 9840 7110 9896
rect 6770 9754 7110 9840
rect 6770 9698 6845 9754
rect 6901 9698 6987 9754
rect 7043 9698 7110 9754
rect 6770 9612 7110 9698
rect 6770 9556 6845 9612
rect 6901 9556 6987 9612
rect 7043 9556 7110 9612
rect 6770 9470 7110 9556
rect 6770 9414 6845 9470
rect 6901 9414 6987 9470
rect 7043 9414 7110 9470
rect 6770 9328 7110 9414
rect 6770 9272 6845 9328
rect 6901 9272 6987 9328
rect 7043 9272 7110 9328
rect 6770 9186 7110 9272
rect 6770 9130 6845 9186
rect 6901 9130 6987 9186
rect 7043 9130 7110 9186
rect 6770 9044 7110 9130
rect 6770 8988 6845 9044
rect 6901 8988 6987 9044
rect 7043 8988 7110 9044
rect 6770 8902 7110 8988
rect 6770 8846 6845 8902
rect 6901 8846 6987 8902
rect 7043 8846 7110 8902
rect 6770 8760 7110 8846
rect 6770 8704 6845 8760
rect 6901 8704 6987 8760
rect 7043 8704 7110 8760
rect 6770 8618 7110 8704
rect 6770 8562 6845 8618
rect 6901 8562 6987 8618
rect 7043 8562 7110 8618
rect 6770 8476 7110 8562
rect 6770 8420 6845 8476
rect 6901 8420 6987 8476
rect 7043 8420 7110 8476
rect 6770 8334 7110 8420
rect 6770 8278 6845 8334
rect 6901 8278 6987 8334
rect 7043 8278 7110 8334
rect 6770 8192 7110 8278
rect 6770 8136 6845 8192
rect 6901 8136 6987 8192
rect 7043 8136 7110 8192
rect 6770 8050 7110 8136
rect 6770 7994 6845 8050
rect 6901 7994 6987 8050
rect 7043 7994 7110 8050
rect 6770 7908 7110 7994
rect 6770 7852 6845 7908
rect 6901 7852 6987 7908
rect 7043 7852 7110 7908
rect 6770 7766 7110 7852
rect 6770 7710 6845 7766
rect 6901 7710 6987 7766
rect 7043 7710 7110 7766
rect 6770 7624 7110 7710
rect 6770 7568 6845 7624
rect 6901 7568 6987 7624
rect 7043 7568 7110 7624
rect 6770 7482 7110 7568
rect 6770 7426 6845 7482
rect 6901 7426 6987 7482
rect 7043 7426 7110 7482
rect 6770 7340 7110 7426
rect 6770 7284 6845 7340
rect 6901 7284 6987 7340
rect 7043 7284 7110 7340
rect 6770 7198 7110 7284
rect 6770 7142 6845 7198
rect 6901 7142 6987 7198
rect 7043 7142 7110 7198
rect 6770 7056 7110 7142
rect 6770 7000 6845 7056
rect 6901 7000 6987 7056
rect 7043 7000 7110 7056
rect 6770 6914 7110 7000
rect 6770 6858 6845 6914
rect 6901 6858 6987 6914
rect 7043 6858 7110 6914
rect 6770 6772 7110 6858
rect 6770 6716 6845 6772
rect 6901 6716 6987 6772
rect 7043 6716 7110 6772
rect 6770 6630 7110 6716
rect 6770 6574 6845 6630
rect 6901 6574 6987 6630
rect 7043 6574 7110 6630
rect 6770 6488 7110 6574
rect 6770 6432 6845 6488
rect 6901 6432 6987 6488
rect 7043 6432 7110 6488
rect 6770 6346 7110 6432
rect 6770 6290 6845 6346
rect 6901 6290 6987 6346
rect 7043 6290 7110 6346
rect 6770 6204 7110 6290
rect 6770 6148 6845 6204
rect 6901 6148 6987 6204
rect 7043 6148 7110 6204
rect 6770 6062 7110 6148
rect 6770 6006 6845 6062
rect 6901 6006 6987 6062
rect 7043 6006 7110 6062
rect 6770 5920 7110 6006
rect 6770 5864 6845 5920
rect 6901 5864 6987 5920
rect 7043 5864 7110 5920
rect 6770 5778 7110 5864
rect 6770 5722 6845 5778
rect 6901 5722 6987 5778
rect 7043 5722 7110 5778
rect 6770 5636 7110 5722
rect 6770 5580 6845 5636
rect 6901 5580 6987 5636
rect 7043 5580 7110 5636
rect 6770 5494 7110 5580
rect 6770 5438 6845 5494
rect 6901 5438 6987 5494
rect 7043 5438 7110 5494
rect 6770 5352 7110 5438
rect 6770 5296 6845 5352
rect 6901 5296 6987 5352
rect 7043 5296 7110 5352
rect 6770 5210 7110 5296
rect 6770 5154 6845 5210
rect 6901 5154 6987 5210
rect 7043 5154 7110 5210
rect 6770 5068 7110 5154
rect 6770 5012 6845 5068
rect 6901 5012 6987 5068
rect 7043 5012 7110 5068
rect 6770 4926 7110 5012
rect 6770 4870 6845 4926
rect 6901 4870 6987 4926
rect 7043 4870 7110 4926
rect 6770 4784 7110 4870
rect 6770 4728 6845 4784
rect 6901 4728 6987 4784
rect 7043 4728 7110 4784
rect 6770 4642 7110 4728
rect 6770 4586 6845 4642
rect 6901 4586 6987 4642
rect 7043 4586 7110 4642
rect 6770 4500 7110 4586
rect 6770 4444 6845 4500
rect 6901 4444 6987 4500
rect 7043 4444 7110 4500
rect 6770 4358 7110 4444
rect 6770 4302 6845 4358
rect 6901 4302 6987 4358
rect 7043 4302 7110 4358
rect 6770 4216 7110 4302
rect 6770 4160 6845 4216
rect 6901 4160 6987 4216
rect 7043 4160 7110 4216
rect 6770 4074 7110 4160
rect 6770 4018 6845 4074
rect 6901 4018 6987 4074
rect 7043 4018 7110 4074
rect 6770 3932 7110 4018
rect 6770 3876 6845 3932
rect 6901 3876 6987 3932
rect 7043 3876 7110 3932
rect 6770 3790 7110 3876
rect 6770 3734 6845 3790
rect 6901 3734 6987 3790
rect 7043 3734 7110 3790
rect 6770 3648 7110 3734
rect 6770 3592 6845 3648
rect 6901 3592 6987 3648
rect 7043 3592 7110 3648
rect 6770 3506 7110 3592
rect 6770 3450 6845 3506
rect 6901 3450 6987 3506
rect 7043 3450 7110 3506
rect 6770 3364 7110 3450
rect 6770 3308 6845 3364
rect 6901 3308 6987 3364
rect 7043 3308 7110 3364
rect 6770 3222 7110 3308
rect 6770 3166 6845 3222
rect 6901 3166 6987 3222
rect 7043 3166 7110 3222
rect 6770 3080 7110 3166
rect 6770 3024 6845 3080
rect 6901 3024 6987 3080
rect 7043 3024 7110 3080
rect 6770 2938 7110 3024
rect 6770 2882 6845 2938
rect 6901 2882 6987 2938
rect 7043 2882 7110 2938
rect 6770 2796 7110 2882
rect 6770 2740 6845 2796
rect 6901 2740 6987 2796
rect 7043 2740 7110 2796
rect 6770 2654 7110 2740
rect 6770 2598 6845 2654
rect 6901 2598 6987 2654
rect 7043 2598 7110 2654
rect 6770 2512 7110 2598
rect 6770 2456 6845 2512
rect 6901 2456 6987 2512
rect 7043 2456 7110 2512
rect 6770 2370 7110 2456
rect 6770 2314 6845 2370
rect 6901 2314 6987 2370
rect 7043 2314 7110 2370
rect 6770 2228 7110 2314
rect 6770 2172 6845 2228
rect 6901 2172 6987 2228
rect 7043 2172 7110 2228
rect 6770 2086 7110 2172
rect 6770 2030 6845 2086
rect 6901 2030 6987 2086
rect 7043 2030 7110 2086
rect 6770 1944 7110 2030
rect 6770 1888 6845 1944
rect 6901 1888 6987 1944
rect 7043 1888 7110 1944
rect 6770 1802 7110 1888
rect 6770 1746 6845 1802
rect 6901 1746 6987 1802
rect 7043 1746 7110 1802
rect 6770 1660 7110 1746
rect 6770 1604 6845 1660
rect 6901 1604 6987 1660
rect 7043 1604 7110 1660
rect 6770 1518 7110 1604
rect 6770 1462 6845 1518
rect 6901 1462 6987 1518
rect 7043 1462 7110 1518
rect 6770 1376 7110 1462
rect 6770 1320 6845 1376
rect 6901 1320 6987 1376
rect 7043 1320 7110 1376
rect 6770 1234 7110 1320
rect 6770 1178 6845 1234
rect 6901 1178 6987 1234
rect 7043 1178 7110 1234
rect 6770 1092 7110 1178
rect 6770 1036 6845 1092
rect 6901 1036 6987 1092
rect 7043 1036 7110 1092
rect 6770 950 7110 1036
rect 6770 894 6845 950
rect 6901 894 6987 950
rect 7043 894 7110 950
rect 6770 808 7110 894
rect 6770 752 6845 808
rect 6901 752 6987 808
rect 7043 752 7110 808
rect 6770 666 7110 752
rect 6770 610 6845 666
rect 6901 610 6987 666
rect 7043 610 7110 666
rect 6770 524 7110 610
rect 6770 468 6845 524
rect 6901 468 6987 524
rect 7043 468 7110 524
rect 6770 400 7110 468
rect 7310 12310 7650 12400
rect 7310 12254 7382 12310
rect 7438 12254 7524 12310
rect 7580 12254 7650 12310
rect 7310 12168 7650 12254
rect 7310 12112 7382 12168
rect 7438 12112 7524 12168
rect 7580 12112 7650 12168
rect 7310 12026 7650 12112
rect 7310 11970 7382 12026
rect 7438 11970 7524 12026
rect 7580 11970 7650 12026
rect 7310 11884 7650 11970
rect 7310 11828 7382 11884
rect 7438 11828 7524 11884
rect 7580 11828 7650 11884
rect 7310 11742 7650 11828
rect 7310 11686 7382 11742
rect 7438 11686 7524 11742
rect 7580 11686 7650 11742
rect 7310 11600 7650 11686
rect 7310 11544 7382 11600
rect 7438 11544 7524 11600
rect 7580 11544 7650 11600
rect 7310 11458 7650 11544
rect 7310 11402 7382 11458
rect 7438 11402 7524 11458
rect 7580 11402 7650 11458
rect 7310 11316 7650 11402
rect 7310 11260 7382 11316
rect 7438 11260 7524 11316
rect 7580 11260 7650 11316
rect 7310 11174 7650 11260
rect 7310 11118 7382 11174
rect 7438 11118 7524 11174
rect 7580 11118 7650 11174
rect 7310 11032 7650 11118
rect 7310 10976 7382 11032
rect 7438 10976 7524 11032
rect 7580 10976 7650 11032
rect 7310 10890 7650 10976
rect 7310 10834 7382 10890
rect 7438 10834 7524 10890
rect 7580 10834 7650 10890
rect 7310 10748 7650 10834
rect 7310 10692 7382 10748
rect 7438 10692 7524 10748
rect 7580 10692 7650 10748
rect 7310 10606 7650 10692
rect 7310 10550 7382 10606
rect 7438 10550 7524 10606
rect 7580 10550 7650 10606
rect 7310 10464 7650 10550
rect 7310 10408 7382 10464
rect 7438 10408 7524 10464
rect 7580 10408 7650 10464
rect 7310 10322 7650 10408
rect 7310 10266 7382 10322
rect 7438 10266 7524 10322
rect 7580 10266 7650 10322
rect 7310 10180 7650 10266
rect 7310 10124 7382 10180
rect 7438 10124 7524 10180
rect 7580 10124 7650 10180
rect 7310 10038 7650 10124
rect 7310 9982 7382 10038
rect 7438 9982 7524 10038
rect 7580 9982 7650 10038
rect 7310 9896 7650 9982
rect 7310 9840 7382 9896
rect 7438 9840 7524 9896
rect 7580 9840 7650 9896
rect 7310 9754 7650 9840
rect 7310 9698 7382 9754
rect 7438 9698 7524 9754
rect 7580 9698 7650 9754
rect 7310 9612 7650 9698
rect 7310 9556 7382 9612
rect 7438 9556 7524 9612
rect 7580 9556 7650 9612
rect 7310 9470 7650 9556
rect 7310 9414 7382 9470
rect 7438 9414 7524 9470
rect 7580 9414 7650 9470
rect 7310 9328 7650 9414
rect 7310 9272 7382 9328
rect 7438 9272 7524 9328
rect 7580 9272 7650 9328
rect 7310 9186 7650 9272
rect 7310 9130 7382 9186
rect 7438 9130 7524 9186
rect 7580 9130 7650 9186
rect 7310 9044 7650 9130
rect 7310 8988 7382 9044
rect 7438 8988 7524 9044
rect 7580 8988 7650 9044
rect 7310 8902 7650 8988
rect 7310 8846 7382 8902
rect 7438 8846 7524 8902
rect 7580 8846 7650 8902
rect 7310 8760 7650 8846
rect 7310 8704 7382 8760
rect 7438 8704 7524 8760
rect 7580 8704 7650 8760
rect 7310 8618 7650 8704
rect 7310 8562 7382 8618
rect 7438 8562 7524 8618
rect 7580 8562 7650 8618
rect 7310 8476 7650 8562
rect 7310 8420 7382 8476
rect 7438 8420 7524 8476
rect 7580 8420 7650 8476
rect 7310 8334 7650 8420
rect 7310 8278 7382 8334
rect 7438 8278 7524 8334
rect 7580 8278 7650 8334
rect 7310 8192 7650 8278
rect 7310 8136 7382 8192
rect 7438 8136 7524 8192
rect 7580 8136 7650 8192
rect 7310 8050 7650 8136
rect 7310 7994 7382 8050
rect 7438 7994 7524 8050
rect 7580 7994 7650 8050
rect 7310 7908 7650 7994
rect 7310 7852 7382 7908
rect 7438 7852 7524 7908
rect 7580 7852 7650 7908
rect 7310 7766 7650 7852
rect 7310 7710 7382 7766
rect 7438 7710 7524 7766
rect 7580 7710 7650 7766
rect 7310 7624 7650 7710
rect 7310 7568 7382 7624
rect 7438 7568 7524 7624
rect 7580 7568 7650 7624
rect 7310 7482 7650 7568
rect 7310 7426 7382 7482
rect 7438 7426 7524 7482
rect 7580 7426 7650 7482
rect 7310 7340 7650 7426
rect 7310 7284 7382 7340
rect 7438 7284 7524 7340
rect 7580 7284 7650 7340
rect 7310 7198 7650 7284
rect 7310 7142 7382 7198
rect 7438 7142 7524 7198
rect 7580 7142 7650 7198
rect 7310 7056 7650 7142
rect 7310 7000 7382 7056
rect 7438 7000 7524 7056
rect 7580 7000 7650 7056
rect 7310 6914 7650 7000
rect 7310 6858 7382 6914
rect 7438 6858 7524 6914
rect 7580 6858 7650 6914
rect 7310 6772 7650 6858
rect 7310 6716 7382 6772
rect 7438 6716 7524 6772
rect 7580 6716 7650 6772
rect 7310 6630 7650 6716
rect 7310 6574 7382 6630
rect 7438 6574 7524 6630
rect 7580 6574 7650 6630
rect 7310 6488 7650 6574
rect 7310 6432 7382 6488
rect 7438 6432 7524 6488
rect 7580 6432 7650 6488
rect 7310 6346 7650 6432
rect 7310 6290 7382 6346
rect 7438 6290 7524 6346
rect 7580 6290 7650 6346
rect 7310 6204 7650 6290
rect 7310 6148 7382 6204
rect 7438 6148 7524 6204
rect 7580 6148 7650 6204
rect 7310 6062 7650 6148
rect 7310 6006 7382 6062
rect 7438 6006 7524 6062
rect 7580 6006 7650 6062
rect 7310 5920 7650 6006
rect 7310 5864 7382 5920
rect 7438 5864 7524 5920
rect 7580 5864 7650 5920
rect 7310 5778 7650 5864
rect 7310 5722 7382 5778
rect 7438 5722 7524 5778
rect 7580 5722 7650 5778
rect 7310 5636 7650 5722
rect 7310 5580 7382 5636
rect 7438 5580 7524 5636
rect 7580 5580 7650 5636
rect 7310 5494 7650 5580
rect 7310 5438 7382 5494
rect 7438 5438 7524 5494
rect 7580 5438 7650 5494
rect 7310 5352 7650 5438
rect 7310 5296 7382 5352
rect 7438 5296 7524 5352
rect 7580 5296 7650 5352
rect 7310 5210 7650 5296
rect 7310 5154 7382 5210
rect 7438 5154 7524 5210
rect 7580 5154 7650 5210
rect 7310 5068 7650 5154
rect 7310 5012 7382 5068
rect 7438 5012 7524 5068
rect 7580 5012 7650 5068
rect 7310 4926 7650 5012
rect 7310 4870 7382 4926
rect 7438 4870 7524 4926
rect 7580 4870 7650 4926
rect 7310 4784 7650 4870
rect 7310 4728 7382 4784
rect 7438 4728 7524 4784
rect 7580 4728 7650 4784
rect 7310 4642 7650 4728
rect 7310 4586 7382 4642
rect 7438 4586 7524 4642
rect 7580 4586 7650 4642
rect 7310 4500 7650 4586
rect 7310 4444 7382 4500
rect 7438 4444 7524 4500
rect 7580 4444 7650 4500
rect 7310 4358 7650 4444
rect 7310 4302 7382 4358
rect 7438 4302 7524 4358
rect 7580 4302 7650 4358
rect 7310 4216 7650 4302
rect 7310 4160 7382 4216
rect 7438 4160 7524 4216
rect 7580 4160 7650 4216
rect 7310 4074 7650 4160
rect 7310 4018 7382 4074
rect 7438 4018 7524 4074
rect 7580 4018 7650 4074
rect 7310 3932 7650 4018
rect 7310 3876 7382 3932
rect 7438 3876 7524 3932
rect 7580 3876 7650 3932
rect 7310 3790 7650 3876
rect 7310 3734 7382 3790
rect 7438 3734 7524 3790
rect 7580 3734 7650 3790
rect 7310 3648 7650 3734
rect 7310 3592 7382 3648
rect 7438 3592 7524 3648
rect 7580 3592 7650 3648
rect 7310 3506 7650 3592
rect 7310 3450 7382 3506
rect 7438 3450 7524 3506
rect 7580 3450 7650 3506
rect 7310 3364 7650 3450
rect 7310 3308 7382 3364
rect 7438 3308 7524 3364
rect 7580 3308 7650 3364
rect 7310 3222 7650 3308
rect 7310 3166 7382 3222
rect 7438 3166 7524 3222
rect 7580 3166 7650 3222
rect 7310 3080 7650 3166
rect 7310 3024 7382 3080
rect 7438 3024 7524 3080
rect 7580 3024 7650 3080
rect 7310 2938 7650 3024
rect 7310 2882 7382 2938
rect 7438 2882 7524 2938
rect 7580 2882 7650 2938
rect 7310 2796 7650 2882
rect 7310 2740 7382 2796
rect 7438 2740 7524 2796
rect 7580 2740 7650 2796
rect 7310 2654 7650 2740
rect 7310 2598 7382 2654
rect 7438 2598 7524 2654
rect 7580 2598 7650 2654
rect 7310 2512 7650 2598
rect 7310 2456 7382 2512
rect 7438 2456 7524 2512
rect 7580 2456 7650 2512
rect 7310 2370 7650 2456
rect 7310 2314 7382 2370
rect 7438 2314 7524 2370
rect 7580 2314 7650 2370
rect 7310 2228 7650 2314
rect 7310 2172 7382 2228
rect 7438 2172 7524 2228
rect 7580 2172 7650 2228
rect 7310 2086 7650 2172
rect 7310 2030 7382 2086
rect 7438 2030 7524 2086
rect 7580 2030 7650 2086
rect 7310 1944 7650 2030
rect 7310 1888 7382 1944
rect 7438 1888 7524 1944
rect 7580 1888 7650 1944
rect 7310 1802 7650 1888
rect 7310 1746 7382 1802
rect 7438 1746 7524 1802
rect 7580 1746 7650 1802
rect 7310 1660 7650 1746
rect 7310 1604 7382 1660
rect 7438 1604 7524 1660
rect 7580 1604 7650 1660
rect 7310 1518 7650 1604
rect 7310 1462 7382 1518
rect 7438 1462 7524 1518
rect 7580 1462 7650 1518
rect 7310 1376 7650 1462
rect 7310 1320 7382 1376
rect 7438 1320 7524 1376
rect 7580 1320 7650 1376
rect 7310 1234 7650 1320
rect 7310 1178 7382 1234
rect 7438 1178 7524 1234
rect 7580 1178 7650 1234
rect 7310 1092 7650 1178
rect 7310 1036 7382 1092
rect 7438 1036 7524 1092
rect 7580 1036 7650 1092
rect 7310 950 7650 1036
rect 7310 894 7382 950
rect 7438 894 7524 950
rect 7580 894 7650 950
rect 7310 808 7650 894
rect 7310 752 7382 808
rect 7438 752 7524 808
rect 7580 752 7650 808
rect 7310 666 7650 752
rect 7310 610 7382 666
rect 7438 610 7524 666
rect 7580 610 7650 666
rect 7310 524 7650 610
rect 7310 468 7382 524
rect 7438 468 7524 524
rect 7580 468 7650 524
rect 7310 400 7650 468
rect 7850 12310 8190 12400
rect 7850 12254 7919 12310
rect 7975 12254 8061 12310
rect 8117 12254 8190 12310
rect 7850 12168 8190 12254
rect 7850 12112 7919 12168
rect 7975 12112 8061 12168
rect 8117 12112 8190 12168
rect 7850 12026 8190 12112
rect 7850 11970 7919 12026
rect 7975 11970 8061 12026
rect 8117 11970 8190 12026
rect 7850 11884 8190 11970
rect 7850 11828 7919 11884
rect 7975 11828 8061 11884
rect 8117 11828 8190 11884
rect 7850 11742 8190 11828
rect 7850 11686 7919 11742
rect 7975 11686 8061 11742
rect 8117 11686 8190 11742
rect 7850 11600 8190 11686
rect 7850 11544 7919 11600
rect 7975 11544 8061 11600
rect 8117 11544 8190 11600
rect 7850 11458 8190 11544
rect 7850 11402 7919 11458
rect 7975 11402 8061 11458
rect 8117 11402 8190 11458
rect 7850 11316 8190 11402
rect 7850 11260 7919 11316
rect 7975 11260 8061 11316
rect 8117 11260 8190 11316
rect 7850 11174 8190 11260
rect 7850 11118 7919 11174
rect 7975 11118 8061 11174
rect 8117 11118 8190 11174
rect 7850 11032 8190 11118
rect 7850 10976 7919 11032
rect 7975 10976 8061 11032
rect 8117 10976 8190 11032
rect 7850 10890 8190 10976
rect 7850 10834 7919 10890
rect 7975 10834 8061 10890
rect 8117 10834 8190 10890
rect 7850 10748 8190 10834
rect 7850 10692 7919 10748
rect 7975 10692 8061 10748
rect 8117 10692 8190 10748
rect 7850 10606 8190 10692
rect 7850 10550 7919 10606
rect 7975 10550 8061 10606
rect 8117 10550 8190 10606
rect 7850 10464 8190 10550
rect 7850 10408 7919 10464
rect 7975 10408 8061 10464
rect 8117 10408 8190 10464
rect 7850 10322 8190 10408
rect 7850 10266 7919 10322
rect 7975 10266 8061 10322
rect 8117 10266 8190 10322
rect 7850 10180 8190 10266
rect 7850 10124 7919 10180
rect 7975 10124 8061 10180
rect 8117 10124 8190 10180
rect 7850 10038 8190 10124
rect 7850 9982 7919 10038
rect 7975 9982 8061 10038
rect 8117 9982 8190 10038
rect 7850 9896 8190 9982
rect 7850 9840 7919 9896
rect 7975 9840 8061 9896
rect 8117 9840 8190 9896
rect 7850 9754 8190 9840
rect 7850 9698 7919 9754
rect 7975 9698 8061 9754
rect 8117 9698 8190 9754
rect 7850 9612 8190 9698
rect 7850 9556 7919 9612
rect 7975 9556 8061 9612
rect 8117 9556 8190 9612
rect 7850 9470 8190 9556
rect 7850 9414 7919 9470
rect 7975 9414 8061 9470
rect 8117 9414 8190 9470
rect 7850 9328 8190 9414
rect 7850 9272 7919 9328
rect 7975 9272 8061 9328
rect 8117 9272 8190 9328
rect 7850 9186 8190 9272
rect 7850 9130 7919 9186
rect 7975 9130 8061 9186
rect 8117 9130 8190 9186
rect 7850 9044 8190 9130
rect 7850 8988 7919 9044
rect 7975 8988 8061 9044
rect 8117 8988 8190 9044
rect 7850 8902 8190 8988
rect 7850 8846 7919 8902
rect 7975 8846 8061 8902
rect 8117 8846 8190 8902
rect 7850 8760 8190 8846
rect 7850 8704 7919 8760
rect 7975 8704 8061 8760
rect 8117 8704 8190 8760
rect 7850 8618 8190 8704
rect 7850 8562 7919 8618
rect 7975 8562 8061 8618
rect 8117 8562 8190 8618
rect 7850 8476 8190 8562
rect 7850 8420 7919 8476
rect 7975 8420 8061 8476
rect 8117 8420 8190 8476
rect 7850 8334 8190 8420
rect 7850 8278 7919 8334
rect 7975 8278 8061 8334
rect 8117 8278 8190 8334
rect 7850 8192 8190 8278
rect 7850 8136 7919 8192
rect 7975 8136 8061 8192
rect 8117 8136 8190 8192
rect 7850 8050 8190 8136
rect 7850 7994 7919 8050
rect 7975 7994 8061 8050
rect 8117 7994 8190 8050
rect 7850 7908 8190 7994
rect 7850 7852 7919 7908
rect 7975 7852 8061 7908
rect 8117 7852 8190 7908
rect 7850 7766 8190 7852
rect 7850 7710 7919 7766
rect 7975 7710 8061 7766
rect 8117 7710 8190 7766
rect 7850 7624 8190 7710
rect 7850 7568 7919 7624
rect 7975 7568 8061 7624
rect 8117 7568 8190 7624
rect 7850 7482 8190 7568
rect 7850 7426 7919 7482
rect 7975 7426 8061 7482
rect 8117 7426 8190 7482
rect 7850 7340 8190 7426
rect 7850 7284 7919 7340
rect 7975 7284 8061 7340
rect 8117 7284 8190 7340
rect 7850 7198 8190 7284
rect 7850 7142 7919 7198
rect 7975 7142 8061 7198
rect 8117 7142 8190 7198
rect 7850 7056 8190 7142
rect 7850 7000 7919 7056
rect 7975 7000 8061 7056
rect 8117 7000 8190 7056
rect 7850 6914 8190 7000
rect 7850 6858 7919 6914
rect 7975 6858 8061 6914
rect 8117 6858 8190 6914
rect 7850 6772 8190 6858
rect 7850 6716 7919 6772
rect 7975 6716 8061 6772
rect 8117 6716 8190 6772
rect 7850 6630 8190 6716
rect 7850 6574 7919 6630
rect 7975 6574 8061 6630
rect 8117 6574 8190 6630
rect 7850 6488 8190 6574
rect 7850 6432 7919 6488
rect 7975 6432 8061 6488
rect 8117 6432 8190 6488
rect 7850 6346 8190 6432
rect 7850 6290 7919 6346
rect 7975 6290 8061 6346
rect 8117 6290 8190 6346
rect 7850 6204 8190 6290
rect 7850 6148 7919 6204
rect 7975 6148 8061 6204
rect 8117 6148 8190 6204
rect 7850 6062 8190 6148
rect 7850 6006 7919 6062
rect 7975 6006 8061 6062
rect 8117 6006 8190 6062
rect 7850 5920 8190 6006
rect 7850 5864 7919 5920
rect 7975 5864 8061 5920
rect 8117 5864 8190 5920
rect 7850 5778 8190 5864
rect 7850 5722 7919 5778
rect 7975 5722 8061 5778
rect 8117 5722 8190 5778
rect 7850 5636 8190 5722
rect 7850 5580 7919 5636
rect 7975 5580 8061 5636
rect 8117 5580 8190 5636
rect 7850 5494 8190 5580
rect 7850 5438 7919 5494
rect 7975 5438 8061 5494
rect 8117 5438 8190 5494
rect 7850 5352 8190 5438
rect 7850 5296 7919 5352
rect 7975 5296 8061 5352
rect 8117 5296 8190 5352
rect 7850 5210 8190 5296
rect 7850 5154 7919 5210
rect 7975 5154 8061 5210
rect 8117 5154 8190 5210
rect 7850 5068 8190 5154
rect 7850 5012 7919 5068
rect 7975 5012 8061 5068
rect 8117 5012 8190 5068
rect 7850 4926 8190 5012
rect 7850 4870 7919 4926
rect 7975 4870 8061 4926
rect 8117 4870 8190 4926
rect 7850 4784 8190 4870
rect 7850 4728 7919 4784
rect 7975 4728 8061 4784
rect 8117 4728 8190 4784
rect 7850 4642 8190 4728
rect 7850 4586 7919 4642
rect 7975 4586 8061 4642
rect 8117 4586 8190 4642
rect 7850 4500 8190 4586
rect 7850 4444 7919 4500
rect 7975 4444 8061 4500
rect 8117 4444 8190 4500
rect 7850 4358 8190 4444
rect 7850 4302 7919 4358
rect 7975 4302 8061 4358
rect 8117 4302 8190 4358
rect 7850 4216 8190 4302
rect 7850 4160 7919 4216
rect 7975 4160 8061 4216
rect 8117 4160 8190 4216
rect 7850 4074 8190 4160
rect 7850 4018 7919 4074
rect 7975 4018 8061 4074
rect 8117 4018 8190 4074
rect 7850 3932 8190 4018
rect 7850 3876 7919 3932
rect 7975 3876 8061 3932
rect 8117 3876 8190 3932
rect 7850 3790 8190 3876
rect 7850 3734 7919 3790
rect 7975 3734 8061 3790
rect 8117 3734 8190 3790
rect 7850 3648 8190 3734
rect 7850 3592 7919 3648
rect 7975 3592 8061 3648
rect 8117 3592 8190 3648
rect 7850 3506 8190 3592
rect 7850 3450 7919 3506
rect 7975 3450 8061 3506
rect 8117 3450 8190 3506
rect 7850 3364 8190 3450
rect 7850 3308 7919 3364
rect 7975 3308 8061 3364
rect 8117 3308 8190 3364
rect 7850 3222 8190 3308
rect 7850 3166 7919 3222
rect 7975 3166 8061 3222
rect 8117 3166 8190 3222
rect 7850 3080 8190 3166
rect 7850 3024 7919 3080
rect 7975 3024 8061 3080
rect 8117 3024 8190 3080
rect 7850 2938 8190 3024
rect 7850 2882 7919 2938
rect 7975 2882 8061 2938
rect 8117 2882 8190 2938
rect 7850 2796 8190 2882
rect 7850 2740 7919 2796
rect 7975 2740 8061 2796
rect 8117 2740 8190 2796
rect 7850 2654 8190 2740
rect 7850 2598 7919 2654
rect 7975 2598 8061 2654
rect 8117 2598 8190 2654
rect 7850 2512 8190 2598
rect 7850 2456 7919 2512
rect 7975 2456 8061 2512
rect 8117 2456 8190 2512
rect 7850 2370 8190 2456
rect 7850 2314 7919 2370
rect 7975 2314 8061 2370
rect 8117 2314 8190 2370
rect 7850 2228 8190 2314
rect 7850 2172 7919 2228
rect 7975 2172 8061 2228
rect 8117 2172 8190 2228
rect 7850 2086 8190 2172
rect 7850 2030 7919 2086
rect 7975 2030 8061 2086
rect 8117 2030 8190 2086
rect 7850 1944 8190 2030
rect 7850 1888 7919 1944
rect 7975 1888 8061 1944
rect 8117 1888 8190 1944
rect 7850 1802 8190 1888
rect 7850 1746 7919 1802
rect 7975 1746 8061 1802
rect 8117 1746 8190 1802
rect 7850 1660 8190 1746
rect 7850 1604 7919 1660
rect 7975 1604 8061 1660
rect 8117 1604 8190 1660
rect 7850 1518 8190 1604
rect 7850 1462 7919 1518
rect 7975 1462 8061 1518
rect 8117 1462 8190 1518
rect 7850 1376 8190 1462
rect 7850 1320 7919 1376
rect 7975 1320 8061 1376
rect 8117 1320 8190 1376
rect 7850 1234 8190 1320
rect 7850 1178 7919 1234
rect 7975 1178 8061 1234
rect 8117 1178 8190 1234
rect 7850 1092 8190 1178
rect 7850 1036 7919 1092
rect 7975 1036 8061 1092
rect 8117 1036 8190 1092
rect 7850 950 8190 1036
rect 7850 894 7919 950
rect 7975 894 8061 950
rect 8117 894 8190 950
rect 7850 808 8190 894
rect 7850 752 7919 808
rect 7975 752 8061 808
rect 8117 752 8190 808
rect 7850 666 8190 752
rect 7850 610 7919 666
rect 7975 610 8061 666
rect 8117 610 8190 666
rect 7850 524 8190 610
rect 7850 468 7919 524
rect 7975 468 8061 524
rect 8117 468 8190 524
rect 7850 400 8190 468
rect 8390 12310 8730 12400
rect 8390 12254 8462 12310
rect 8518 12254 8604 12310
rect 8660 12254 8730 12310
rect 8390 12168 8730 12254
rect 8390 12112 8462 12168
rect 8518 12112 8604 12168
rect 8660 12112 8730 12168
rect 8390 12026 8730 12112
rect 8390 11970 8462 12026
rect 8518 11970 8604 12026
rect 8660 11970 8730 12026
rect 8390 11884 8730 11970
rect 8390 11828 8462 11884
rect 8518 11828 8604 11884
rect 8660 11828 8730 11884
rect 8390 11742 8730 11828
rect 8390 11686 8462 11742
rect 8518 11686 8604 11742
rect 8660 11686 8730 11742
rect 8390 11600 8730 11686
rect 8390 11544 8462 11600
rect 8518 11544 8604 11600
rect 8660 11544 8730 11600
rect 8390 11458 8730 11544
rect 8390 11402 8462 11458
rect 8518 11402 8604 11458
rect 8660 11402 8730 11458
rect 8390 11316 8730 11402
rect 8390 11260 8462 11316
rect 8518 11260 8604 11316
rect 8660 11260 8730 11316
rect 8390 11174 8730 11260
rect 8390 11118 8462 11174
rect 8518 11118 8604 11174
rect 8660 11118 8730 11174
rect 8390 11032 8730 11118
rect 8390 10976 8462 11032
rect 8518 10976 8604 11032
rect 8660 10976 8730 11032
rect 8390 10890 8730 10976
rect 8390 10834 8462 10890
rect 8518 10834 8604 10890
rect 8660 10834 8730 10890
rect 8390 10748 8730 10834
rect 8390 10692 8462 10748
rect 8518 10692 8604 10748
rect 8660 10692 8730 10748
rect 8390 10606 8730 10692
rect 8390 10550 8462 10606
rect 8518 10550 8604 10606
rect 8660 10550 8730 10606
rect 8390 10464 8730 10550
rect 8390 10408 8462 10464
rect 8518 10408 8604 10464
rect 8660 10408 8730 10464
rect 8390 10322 8730 10408
rect 8390 10266 8462 10322
rect 8518 10266 8604 10322
rect 8660 10266 8730 10322
rect 8390 10180 8730 10266
rect 8390 10124 8462 10180
rect 8518 10124 8604 10180
rect 8660 10124 8730 10180
rect 8390 10038 8730 10124
rect 8390 9982 8462 10038
rect 8518 9982 8604 10038
rect 8660 9982 8730 10038
rect 8390 9896 8730 9982
rect 8390 9840 8462 9896
rect 8518 9840 8604 9896
rect 8660 9840 8730 9896
rect 8390 9754 8730 9840
rect 8390 9698 8462 9754
rect 8518 9698 8604 9754
rect 8660 9698 8730 9754
rect 8390 9612 8730 9698
rect 8390 9556 8462 9612
rect 8518 9556 8604 9612
rect 8660 9556 8730 9612
rect 8390 9470 8730 9556
rect 8390 9414 8462 9470
rect 8518 9414 8604 9470
rect 8660 9414 8730 9470
rect 8390 9328 8730 9414
rect 8390 9272 8462 9328
rect 8518 9272 8604 9328
rect 8660 9272 8730 9328
rect 8390 9186 8730 9272
rect 8390 9130 8462 9186
rect 8518 9130 8604 9186
rect 8660 9130 8730 9186
rect 8390 9044 8730 9130
rect 8390 8988 8462 9044
rect 8518 8988 8604 9044
rect 8660 8988 8730 9044
rect 8390 8902 8730 8988
rect 8390 8846 8462 8902
rect 8518 8846 8604 8902
rect 8660 8846 8730 8902
rect 8390 8760 8730 8846
rect 8390 8704 8462 8760
rect 8518 8704 8604 8760
rect 8660 8704 8730 8760
rect 8390 8618 8730 8704
rect 8390 8562 8462 8618
rect 8518 8562 8604 8618
rect 8660 8562 8730 8618
rect 8390 8476 8730 8562
rect 8390 8420 8462 8476
rect 8518 8420 8604 8476
rect 8660 8420 8730 8476
rect 8390 8334 8730 8420
rect 8390 8278 8462 8334
rect 8518 8278 8604 8334
rect 8660 8278 8730 8334
rect 8390 8192 8730 8278
rect 8390 8136 8462 8192
rect 8518 8136 8604 8192
rect 8660 8136 8730 8192
rect 8390 8050 8730 8136
rect 8390 7994 8462 8050
rect 8518 7994 8604 8050
rect 8660 7994 8730 8050
rect 8390 7908 8730 7994
rect 8390 7852 8462 7908
rect 8518 7852 8604 7908
rect 8660 7852 8730 7908
rect 8390 7766 8730 7852
rect 8390 7710 8462 7766
rect 8518 7710 8604 7766
rect 8660 7710 8730 7766
rect 8390 7624 8730 7710
rect 8390 7568 8462 7624
rect 8518 7568 8604 7624
rect 8660 7568 8730 7624
rect 8390 7482 8730 7568
rect 8390 7426 8462 7482
rect 8518 7426 8604 7482
rect 8660 7426 8730 7482
rect 8390 7340 8730 7426
rect 8390 7284 8462 7340
rect 8518 7284 8604 7340
rect 8660 7284 8730 7340
rect 8390 7198 8730 7284
rect 8390 7142 8462 7198
rect 8518 7142 8604 7198
rect 8660 7142 8730 7198
rect 8390 7056 8730 7142
rect 8390 7000 8462 7056
rect 8518 7000 8604 7056
rect 8660 7000 8730 7056
rect 8390 6914 8730 7000
rect 8390 6858 8462 6914
rect 8518 6858 8604 6914
rect 8660 6858 8730 6914
rect 8390 6772 8730 6858
rect 8390 6716 8462 6772
rect 8518 6716 8604 6772
rect 8660 6716 8730 6772
rect 8390 6630 8730 6716
rect 8390 6574 8462 6630
rect 8518 6574 8604 6630
rect 8660 6574 8730 6630
rect 8390 6488 8730 6574
rect 8390 6432 8462 6488
rect 8518 6432 8604 6488
rect 8660 6432 8730 6488
rect 8390 6346 8730 6432
rect 8390 6290 8462 6346
rect 8518 6290 8604 6346
rect 8660 6290 8730 6346
rect 8390 6204 8730 6290
rect 8390 6148 8462 6204
rect 8518 6148 8604 6204
rect 8660 6148 8730 6204
rect 8390 6062 8730 6148
rect 8390 6006 8462 6062
rect 8518 6006 8604 6062
rect 8660 6006 8730 6062
rect 8390 5920 8730 6006
rect 8390 5864 8462 5920
rect 8518 5864 8604 5920
rect 8660 5864 8730 5920
rect 8390 5778 8730 5864
rect 8390 5722 8462 5778
rect 8518 5722 8604 5778
rect 8660 5722 8730 5778
rect 8390 5636 8730 5722
rect 8390 5580 8462 5636
rect 8518 5580 8604 5636
rect 8660 5580 8730 5636
rect 8390 5494 8730 5580
rect 8390 5438 8462 5494
rect 8518 5438 8604 5494
rect 8660 5438 8730 5494
rect 8390 5352 8730 5438
rect 8390 5296 8462 5352
rect 8518 5296 8604 5352
rect 8660 5296 8730 5352
rect 8390 5210 8730 5296
rect 8390 5154 8462 5210
rect 8518 5154 8604 5210
rect 8660 5154 8730 5210
rect 8390 5068 8730 5154
rect 8390 5012 8462 5068
rect 8518 5012 8604 5068
rect 8660 5012 8730 5068
rect 8390 4926 8730 5012
rect 8390 4870 8462 4926
rect 8518 4870 8604 4926
rect 8660 4870 8730 4926
rect 8390 4784 8730 4870
rect 8390 4728 8462 4784
rect 8518 4728 8604 4784
rect 8660 4728 8730 4784
rect 8390 4642 8730 4728
rect 8390 4586 8462 4642
rect 8518 4586 8604 4642
rect 8660 4586 8730 4642
rect 8390 4500 8730 4586
rect 8390 4444 8462 4500
rect 8518 4444 8604 4500
rect 8660 4444 8730 4500
rect 8390 4358 8730 4444
rect 8390 4302 8462 4358
rect 8518 4302 8604 4358
rect 8660 4302 8730 4358
rect 8390 4216 8730 4302
rect 8390 4160 8462 4216
rect 8518 4160 8604 4216
rect 8660 4160 8730 4216
rect 8390 4074 8730 4160
rect 8390 4018 8462 4074
rect 8518 4018 8604 4074
rect 8660 4018 8730 4074
rect 8390 3932 8730 4018
rect 8390 3876 8462 3932
rect 8518 3876 8604 3932
rect 8660 3876 8730 3932
rect 8390 3790 8730 3876
rect 8390 3734 8462 3790
rect 8518 3734 8604 3790
rect 8660 3734 8730 3790
rect 8390 3648 8730 3734
rect 8390 3592 8462 3648
rect 8518 3592 8604 3648
rect 8660 3592 8730 3648
rect 8390 3506 8730 3592
rect 8390 3450 8462 3506
rect 8518 3450 8604 3506
rect 8660 3450 8730 3506
rect 8390 3364 8730 3450
rect 8390 3308 8462 3364
rect 8518 3308 8604 3364
rect 8660 3308 8730 3364
rect 8390 3222 8730 3308
rect 8390 3166 8462 3222
rect 8518 3166 8604 3222
rect 8660 3166 8730 3222
rect 8390 3080 8730 3166
rect 8390 3024 8462 3080
rect 8518 3024 8604 3080
rect 8660 3024 8730 3080
rect 8390 2938 8730 3024
rect 8390 2882 8462 2938
rect 8518 2882 8604 2938
rect 8660 2882 8730 2938
rect 8390 2796 8730 2882
rect 8390 2740 8462 2796
rect 8518 2740 8604 2796
rect 8660 2740 8730 2796
rect 8390 2654 8730 2740
rect 8390 2598 8462 2654
rect 8518 2598 8604 2654
rect 8660 2598 8730 2654
rect 8390 2512 8730 2598
rect 8390 2456 8462 2512
rect 8518 2456 8604 2512
rect 8660 2456 8730 2512
rect 8390 2370 8730 2456
rect 8390 2314 8462 2370
rect 8518 2314 8604 2370
rect 8660 2314 8730 2370
rect 8390 2228 8730 2314
rect 8390 2172 8462 2228
rect 8518 2172 8604 2228
rect 8660 2172 8730 2228
rect 8390 2086 8730 2172
rect 8390 2030 8462 2086
rect 8518 2030 8604 2086
rect 8660 2030 8730 2086
rect 8390 1944 8730 2030
rect 8390 1888 8462 1944
rect 8518 1888 8604 1944
rect 8660 1888 8730 1944
rect 8390 1802 8730 1888
rect 8390 1746 8462 1802
rect 8518 1746 8604 1802
rect 8660 1746 8730 1802
rect 8390 1660 8730 1746
rect 8390 1604 8462 1660
rect 8518 1604 8604 1660
rect 8660 1604 8730 1660
rect 8390 1518 8730 1604
rect 8390 1462 8462 1518
rect 8518 1462 8604 1518
rect 8660 1462 8730 1518
rect 8390 1376 8730 1462
rect 8390 1320 8462 1376
rect 8518 1320 8604 1376
rect 8660 1320 8730 1376
rect 8390 1234 8730 1320
rect 8390 1178 8462 1234
rect 8518 1178 8604 1234
rect 8660 1178 8730 1234
rect 8390 1092 8730 1178
rect 8390 1036 8462 1092
rect 8518 1036 8604 1092
rect 8660 1036 8730 1092
rect 8390 950 8730 1036
rect 8390 894 8462 950
rect 8518 894 8604 950
rect 8660 894 8730 950
rect 8390 808 8730 894
rect 8390 752 8462 808
rect 8518 752 8604 808
rect 8660 752 8730 808
rect 8390 666 8730 752
rect 8390 610 8462 666
rect 8518 610 8604 666
rect 8660 610 8730 666
rect 8390 524 8730 610
rect 8390 468 8462 524
rect 8518 468 8604 524
rect 8660 468 8730 524
rect 8390 400 8730 468
rect 8930 12310 9270 12400
rect 8930 12254 9004 12310
rect 9060 12254 9146 12310
rect 9202 12254 9270 12310
rect 8930 12168 9270 12254
rect 8930 12112 9004 12168
rect 9060 12112 9146 12168
rect 9202 12112 9270 12168
rect 8930 12026 9270 12112
rect 8930 11970 9004 12026
rect 9060 11970 9146 12026
rect 9202 11970 9270 12026
rect 8930 11884 9270 11970
rect 8930 11828 9004 11884
rect 9060 11828 9146 11884
rect 9202 11828 9270 11884
rect 8930 11742 9270 11828
rect 8930 11686 9004 11742
rect 9060 11686 9146 11742
rect 9202 11686 9270 11742
rect 8930 11600 9270 11686
rect 8930 11544 9004 11600
rect 9060 11544 9146 11600
rect 9202 11544 9270 11600
rect 8930 11458 9270 11544
rect 8930 11402 9004 11458
rect 9060 11402 9146 11458
rect 9202 11402 9270 11458
rect 8930 11316 9270 11402
rect 8930 11260 9004 11316
rect 9060 11260 9146 11316
rect 9202 11260 9270 11316
rect 8930 11174 9270 11260
rect 8930 11118 9004 11174
rect 9060 11118 9146 11174
rect 9202 11118 9270 11174
rect 8930 11032 9270 11118
rect 8930 10976 9004 11032
rect 9060 10976 9146 11032
rect 9202 10976 9270 11032
rect 8930 10890 9270 10976
rect 8930 10834 9004 10890
rect 9060 10834 9146 10890
rect 9202 10834 9270 10890
rect 8930 10748 9270 10834
rect 8930 10692 9004 10748
rect 9060 10692 9146 10748
rect 9202 10692 9270 10748
rect 8930 10606 9270 10692
rect 8930 10550 9004 10606
rect 9060 10550 9146 10606
rect 9202 10550 9270 10606
rect 8930 10464 9270 10550
rect 8930 10408 9004 10464
rect 9060 10408 9146 10464
rect 9202 10408 9270 10464
rect 8930 10322 9270 10408
rect 8930 10266 9004 10322
rect 9060 10266 9146 10322
rect 9202 10266 9270 10322
rect 8930 10180 9270 10266
rect 8930 10124 9004 10180
rect 9060 10124 9146 10180
rect 9202 10124 9270 10180
rect 8930 10038 9270 10124
rect 8930 9982 9004 10038
rect 9060 9982 9146 10038
rect 9202 9982 9270 10038
rect 8930 9896 9270 9982
rect 8930 9840 9004 9896
rect 9060 9840 9146 9896
rect 9202 9840 9270 9896
rect 8930 9754 9270 9840
rect 8930 9698 9004 9754
rect 9060 9698 9146 9754
rect 9202 9698 9270 9754
rect 8930 9612 9270 9698
rect 8930 9556 9004 9612
rect 9060 9556 9146 9612
rect 9202 9556 9270 9612
rect 8930 9470 9270 9556
rect 8930 9414 9004 9470
rect 9060 9414 9146 9470
rect 9202 9414 9270 9470
rect 8930 9328 9270 9414
rect 8930 9272 9004 9328
rect 9060 9272 9146 9328
rect 9202 9272 9270 9328
rect 8930 9186 9270 9272
rect 8930 9130 9004 9186
rect 9060 9130 9146 9186
rect 9202 9130 9270 9186
rect 8930 9044 9270 9130
rect 8930 8988 9004 9044
rect 9060 8988 9146 9044
rect 9202 8988 9270 9044
rect 8930 8902 9270 8988
rect 8930 8846 9004 8902
rect 9060 8846 9146 8902
rect 9202 8846 9270 8902
rect 8930 8760 9270 8846
rect 8930 8704 9004 8760
rect 9060 8704 9146 8760
rect 9202 8704 9270 8760
rect 8930 8618 9270 8704
rect 8930 8562 9004 8618
rect 9060 8562 9146 8618
rect 9202 8562 9270 8618
rect 8930 8476 9270 8562
rect 8930 8420 9004 8476
rect 9060 8420 9146 8476
rect 9202 8420 9270 8476
rect 8930 8334 9270 8420
rect 8930 8278 9004 8334
rect 9060 8278 9146 8334
rect 9202 8278 9270 8334
rect 8930 8192 9270 8278
rect 8930 8136 9004 8192
rect 9060 8136 9146 8192
rect 9202 8136 9270 8192
rect 8930 8050 9270 8136
rect 8930 7994 9004 8050
rect 9060 7994 9146 8050
rect 9202 7994 9270 8050
rect 8930 7908 9270 7994
rect 8930 7852 9004 7908
rect 9060 7852 9146 7908
rect 9202 7852 9270 7908
rect 8930 7766 9270 7852
rect 8930 7710 9004 7766
rect 9060 7710 9146 7766
rect 9202 7710 9270 7766
rect 8930 7624 9270 7710
rect 8930 7568 9004 7624
rect 9060 7568 9146 7624
rect 9202 7568 9270 7624
rect 8930 7482 9270 7568
rect 8930 7426 9004 7482
rect 9060 7426 9146 7482
rect 9202 7426 9270 7482
rect 8930 7340 9270 7426
rect 8930 7284 9004 7340
rect 9060 7284 9146 7340
rect 9202 7284 9270 7340
rect 8930 7198 9270 7284
rect 8930 7142 9004 7198
rect 9060 7142 9146 7198
rect 9202 7142 9270 7198
rect 8930 7056 9270 7142
rect 8930 7000 9004 7056
rect 9060 7000 9146 7056
rect 9202 7000 9270 7056
rect 8930 6914 9270 7000
rect 8930 6858 9004 6914
rect 9060 6858 9146 6914
rect 9202 6858 9270 6914
rect 8930 6772 9270 6858
rect 8930 6716 9004 6772
rect 9060 6716 9146 6772
rect 9202 6716 9270 6772
rect 8930 6630 9270 6716
rect 8930 6574 9004 6630
rect 9060 6574 9146 6630
rect 9202 6574 9270 6630
rect 8930 6488 9270 6574
rect 8930 6432 9004 6488
rect 9060 6432 9146 6488
rect 9202 6432 9270 6488
rect 8930 6346 9270 6432
rect 8930 6290 9004 6346
rect 9060 6290 9146 6346
rect 9202 6290 9270 6346
rect 8930 6204 9270 6290
rect 8930 6148 9004 6204
rect 9060 6148 9146 6204
rect 9202 6148 9270 6204
rect 8930 6062 9270 6148
rect 8930 6006 9004 6062
rect 9060 6006 9146 6062
rect 9202 6006 9270 6062
rect 8930 5920 9270 6006
rect 8930 5864 9004 5920
rect 9060 5864 9146 5920
rect 9202 5864 9270 5920
rect 8930 5778 9270 5864
rect 8930 5722 9004 5778
rect 9060 5722 9146 5778
rect 9202 5722 9270 5778
rect 8930 5636 9270 5722
rect 8930 5580 9004 5636
rect 9060 5580 9146 5636
rect 9202 5580 9270 5636
rect 8930 5494 9270 5580
rect 8930 5438 9004 5494
rect 9060 5438 9146 5494
rect 9202 5438 9270 5494
rect 8930 5352 9270 5438
rect 8930 5296 9004 5352
rect 9060 5296 9146 5352
rect 9202 5296 9270 5352
rect 8930 5210 9270 5296
rect 8930 5154 9004 5210
rect 9060 5154 9146 5210
rect 9202 5154 9270 5210
rect 8930 5068 9270 5154
rect 8930 5012 9004 5068
rect 9060 5012 9146 5068
rect 9202 5012 9270 5068
rect 8930 4926 9270 5012
rect 8930 4870 9004 4926
rect 9060 4870 9146 4926
rect 9202 4870 9270 4926
rect 8930 4784 9270 4870
rect 8930 4728 9004 4784
rect 9060 4728 9146 4784
rect 9202 4728 9270 4784
rect 8930 4642 9270 4728
rect 8930 4586 9004 4642
rect 9060 4586 9146 4642
rect 9202 4586 9270 4642
rect 8930 4500 9270 4586
rect 8930 4444 9004 4500
rect 9060 4444 9146 4500
rect 9202 4444 9270 4500
rect 8930 4358 9270 4444
rect 8930 4302 9004 4358
rect 9060 4302 9146 4358
rect 9202 4302 9270 4358
rect 8930 4216 9270 4302
rect 8930 4160 9004 4216
rect 9060 4160 9146 4216
rect 9202 4160 9270 4216
rect 8930 4074 9270 4160
rect 8930 4018 9004 4074
rect 9060 4018 9146 4074
rect 9202 4018 9270 4074
rect 8930 3932 9270 4018
rect 8930 3876 9004 3932
rect 9060 3876 9146 3932
rect 9202 3876 9270 3932
rect 8930 3790 9270 3876
rect 8930 3734 9004 3790
rect 9060 3734 9146 3790
rect 9202 3734 9270 3790
rect 8930 3648 9270 3734
rect 8930 3592 9004 3648
rect 9060 3592 9146 3648
rect 9202 3592 9270 3648
rect 8930 3506 9270 3592
rect 8930 3450 9004 3506
rect 9060 3450 9146 3506
rect 9202 3450 9270 3506
rect 8930 3364 9270 3450
rect 8930 3308 9004 3364
rect 9060 3308 9146 3364
rect 9202 3308 9270 3364
rect 8930 3222 9270 3308
rect 8930 3166 9004 3222
rect 9060 3166 9146 3222
rect 9202 3166 9270 3222
rect 8930 3080 9270 3166
rect 8930 3024 9004 3080
rect 9060 3024 9146 3080
rect 9202 3024 9270 3080
rect 8930 2938 9270 3024
rect 8930 2882 9004 2938
rect 9060 2882 9146 2938
rect 9202 2882 9270 2938
rect 8930 2796 9270 2882
rect 8930 2740 9004 2796
rect 9060 2740 9146 2796
rect 9202 2740 9270 2796
rect 8930 2654 9270 2740
rect 8930 2598 9004 2654
rect 9060 2598 9146 2654
rect 9202 2598 9270 2654
rect 8930 2512 9270 2598
rect 8930 2456 9004 2512
rect 9060 2456 9146 2512
rect 9202 2456 9270 2512
rect 8930 2370 9270 2456
rect 8930 2314 9004 2370
rect 9060 2314 9146 2370
rect 9202 2314 9270 2370
rect 8930 2228 9270 2314
rect 8930 2172 9004 2228
rect 9060 2172 9146 2228
rect 9202 2172 9270 2228
rect 8930 2086 9270 2172
rect 8930 2030 9004 2086
rect 9060 2030 9146 2086
rect 9202 2030 9270 2086
rect 8930 1944 9270 2030
rect 8930 1888 9004 1944
rect 9060 1888 9146 1944
rect 9202 1888 9270 1944
rect 8930 1802 9270 1888
rect 8930 1746 9004 1802
rect 9060 1746 9146 1802
rect 9202 1746 9270 1802
rect 8930 1660 9270 1746
rect 8930 1604 9004 1660
rect 9060 1604 9146 1660
rect 9202 1604 9270 1660
rect 8930 1518 9270 1604
rect 8930 1462 9004 1518
rect 9060 1462 9146 1518
rect 9202 1462 9270 1518
rect 8930 1376 9270 1462
rect 8930 1320 9004 1376
rect 9060 1320 9146 1376
rect 9202 1320 9270 1376
rect 8930 1234 9270 1320
rect 8930 1178 9004 1234
rect 9060 1178 9146 1234
rect 9202 1178 9270 1234
rect 8930 1092 9270 1178
rect 8930 1036 9004 1092
rect 9060 1036 9146 1092
rect 9202 1036 9270 1092
rect 8930 950 9270 1036
rect 8930 894 9004 950
rect 9060 894 9146 950
rect 9202 894 9270 950
rect 8930 808 9270 894
rect 8930 752 9004 808
rect 9060 752 9146 808
rect 9202 752 9270 808
rect 8930 666 9270 752
rect 8930 610 9004 666
rect 9060 610 9146 666
rect 9202 610 9270 666
rect 8930 524 9270 610
rect 8930 468 9004 524
rect 9060 468 9146 524
rect 9202 468 9270 524
rect 8930 400 9270 468
rect 9470 12310 9810 12400
rect 9470 12254 9547 12310
rect 9603 12254 9689 12310
rect 9745 12254 9810 12310
rect 9470 12168 9810 12254
rect 9470 12112 9547 12168
rect 9603 12112 9689 12168
rect 9745 12112 9810 12168
rect 9470 12026 9810 12112
rect 9470 11970 9547 12026
rect 9603 11970 9689 12026
rect 9745 11970 9810 12026
rect 9470 11884 9810 11970
rect 9470 11828 9547 11884
rect 9603 11828 9689 11884
rect 9745 11828 9810 11884
rect 9470 11742 9810 11828
rect 9470 11686 9547 11742
rect 9603 11686 9689 11742
rect 9745 11686 9810 11742
rect 9470 11600 9810 11686
rect 9470 11544 9547 11600
rect 9603 11544 9689 11600
rect 9745 11544 9810 11600
rect 9470 11458 9810 11544
rect 9470 11402 9547 11458
rect 9603 11402 9689 11458
rect 9745 11402 9810 11458
rect 9470 11316 9810 11402
rect 9470 11260 9547 11316
rect 9603 11260 9689 11316
rect 9745 11260 9810 11316
rect 9470 11174 9810 11260
rect 9470 11118 9547 11174
rect 9603 11118 9689 11174
rect 9745 11118 9810 11174
rect 9470 11032 9810 11118
rect 9470 10976 9547 11032
rect 9603 10976 9689 11032
rect 9745 10976 9810 11032
rect 9470 10890 9810 10976
rect 9470 10834 9547 10890
rect 9603 10834 9689 10890
rect 9745 10834 9810 10890
rect 9470 10748 9810 10834
rect 9470 10692 9547 10748
rect 9603 10692 9689 10748
rect 9745 10692 9810 10748
rect 9470 10606 9810 10692
rect 9470 10550 9547 10606
rect 9603 10550 9689 10606
rect 9745 10550 9810 10606
rect 9470 10464 9810 10550
rect 9470 10408 9547 10464
rect 9603 10408 9689 10464
rect 9745 10408 9810 10464
rect 9470 10322 9810 10408
rect 9470 10266 9547 10322
rect 9603 10266 9689 10322
rect 9745 10266 9810 10322
rect 9470 10180 9810 10266
rect 9470 10124 9547 10180
rect 9603 10124 9689 10180
rect 9745 10124 9810 10180
rect 9470 10038 9810 10124
rect 9470 9982 9547 10038
rect 9603 9982 9689 10038
rect 9745 9982 9810 10038
rect 9470 9896 9810 9982
rect 9470 9840 9547 9896
rect 9603 9840 9689 9896
rect 9745 9840 9810 9896
rect 9470 9754 9810 9840
rect 9470 9698 9547 9754
rect 9603 9698 9689 9754
rect 9745 9698 9810 9754
rect 9470 9612 9810 9698
rect 9470 9556 9547 9612
rect 9603 9556 9689 9612
rect 9745 9556 9810 9612
rect 9470 9470 9810 9556
rect 9470 9414 9547 9470
rect 9603 9414 9689 9470
rect 9745 9414 9810 9470
rect 9470 9328 9810 9414
rect 9470 9272 9547 9328
rect 9603 9272 9689 9328
rect 9745 9272 9810 9328
rect 9470 9186 9810 9272
rect 9470 9130 9547 9186
rect 9603 9130 9689 9186
rect 9745 9130 9810 9186
rect 9470 9044 9810 9130
rect 9470 8988 9547 9044
rect 9603 8988 9689 9044
rect 9745 8988 9810 9044
rect 9470 8902 9810 8988
rect 9470 8846 9547 8902
rect 9603 8846 9689 8902
rect 9745 8846 9810 8902
rect 9470 8760 9810 8846
rect 9470 8704 9547 8760
rect 9603 8704 9689 8760
rect 9745 8704 9810 8760
rect 9470 8618 9810 8704
rect 9470 8562 9547 8618
rect 9603 8562 9689 8618
rect 9745 8562 9810 8618
rect 9470 8476 9810 8562
rect 9470 8420 9547 8476
rect 9603 8420 9689 8476
rect 9745 8420 9810 8476
rect 9470 8334 9810 8420
rect 9470 8278 9547 8334
rect 9603 8278 9689 8334
rect 9745 8278 9810 8334
rect 9470 8192 9810 8278
rect 9470 8136 9547 8192
rect 9603 8136 9689 8192
rect 9745 8136 9810 8192
rect 9470 8050 9810 8136
rect 9470 7994 9547 8050
rect 9603 7994 9689 8050
rect 9745 7994 9810 8050
rect 9470 7908 9810 7994
rect 9470 7852 9547 7908
rect 9603 7852 9689 7908
rect 9745 7852 9810 7908
rect 9470 7766 9810 7852
rect 9470 7710 9547 7766
rect 9603 7710 9689 7766
rect 9745 7710 9810 7766
rect 9470 7624 9810 7710
rect 9470 7568 9547 7624
rect 9603 7568 9689 7624
rect 9745 7568 9810 7624
rect 9470 7482 9810 7568
rect 9470 7426 9547 7482
rect 9603 7426 9689 7482
rect 9745 7426 9810 7482
rect 9470 7340 9810 7426
rect 9470 7284 9547 7340
rect 9603 7284 9689 7340
rect 9745 7284 9810 7340
rect 9470 7198 9810 7284
rect 9470 7142 9547 7198
rect 9603 7142 9689 7198
rect 9745 7142 9810 7198
rect 9470 7056 9810 7142
rect 9470 7000 9547 7056
rect 9603 7000 9689 7056
rect 9745 7000 9810 7056
rect 9470 6914 9810 7000
rect 9470 6858 9547 6914
rect 9603 6858 9689 6914
rect 9745 6858 9810 6914
rect 9470 6772 9810 6858
rect 9470 6716 9547 6772
rect 9603 6716 9689 6772
rect 9745 6716 9810 6772
rect 9470 6630 9810 6716
rect 9470 6574 9547 6630
rect 9603 6574 9689 6630
rect 9745 6574 9810 6630
rect 9470 6488 9810 6574
rect 9470 6432 9547 6488
rect 9603 6432 9689 6488
rect 9745 6432 9810 6488
rect 9470 6346 9810 6432
rect 9470 6290 9547 6346
rect 9603 6290 9689 6346
rect 9745 6290 9810 6346
rect 9470 6204 9810 6290
rect 9470 6148 9547 6204
rect 9603 6148 9689 6204
rect 9745 6148 9810 6204
rect 9470 6062 9810 6148
rect 9470 6006 9547 6062
rect 9603 6006 9689 6062
rect 9745 6006 9810 6062
rect 9470 5920 9810 6006
rect 9470 5864 9547 5920
rect 9603 5864 9689 5920
rect 9745 5864 9810 5920
rect 9470 5778 9810 5864
rect 9470 5722 9547 5778
rect 9603 5722 9689 5778
rect 9745 5722 9810 5778
rect 9470 5636 9810 5722
rect 9470 5580 9547 5636
rect 9603 5580 9689 5636
rect 9745 5580 9810 5636
rect 9470 5494 9810 5580
rect 9470 5438 9547 5494
rect 9603 5438 9689 5494
rect 9745 5438 9810 5494
rect 9470 5352 9810 5438
rect 9470 5296 9547 5352
rect 9603 5296 9689 5352
rect 9745 5296 9810 5352
rect 9470 5210 9810 5296
rect 9470 5154 9547 5210
rect 9603 5154 9689 5210
rect 9745 5154 9810 5210
rect 9470 5068 9810 5154
rect 9470 5012 9547 5068
rect 9603 5012 9689 5068
rect 9745 5012 9810 5068
rect 9470 4926 9810 5012
rect 9470 4870 9547 4926
rect 9603 4870 9689 4926
rect 9745 4870 9810 4926
rect 9470 4784 9810 4870
rect 9470 4728 9547 4784
rect 9603 4728 9689 4784
rect 9745 4728 9810 4784
rect 9470 4642 9810 4728
rect 9470 4586 9547 4642
rect 9603 4586 9689 4642
rect 9745 4586 9810 4642
rect 9470 4500 9810 4586
rect 9470 4444 9547 4500
rect 9603 4444 9689 4500
rect 9745 4444 9810 4500
rect 9470 4358 9810 4444
rect 9470 4302 9547 4358
rect 9603 4302 9689 4358
rect 9745 4302 9810 4358
rect 9470 4216 9810 4302
rect 9470 4160 9547 4216
rect 9603 4160 9689 4216
rect 9745 4160 9810 4216
rect 9470 4074 9810 4160
rect 9470 4018 9547 4074
rect 9603 4018 9689 4074
rect 9745 4018 9810 4074
rect 9470 3932 9810 4018
rect 9470 3876 9547 3932
rect 9603 3876 9689 3932
rect 9745 3876 9810 3932
rect 9470 3790 9810 3876
rect 9470 3734 9547 3790
rect 9603 3734 9689 3790
rect 9745 3734 9810 3790
rect 9470 3648 9810 3734
rect 9470 3592 9547 3648
rect 9603 3592 9689 3648
rect 9745 3592 9810 3648
rect 9470 3506 9810 3592
rect 9470 3450 9547 3506
rect 9603 3450 9689 3506
rect 9745 3450 9810 3506
rect 9470 3364 9810 3450
rect 9470 3308 9547 3364
rect 9603 3308 9689 3364
rect 9745 3308 9810 3364
rect 9470 3222 9810 3308
rect 9470 3166 9547 3222
rect 9603 3166 9689 3222
rect 9745 3166 9810 3222
rect 9470 3080 9810 3166
rect 9470 3024 9547 3080
rect 9603 3024 9689 3080
rect 9745 3024 9810 3080
rect 9470 2938 9810 3024
rect 9470 2882 9547 2938
rect 9603 2882 9689 2938
rect 9745 2882 9810 2938
rect 9470 2796 9810 2882
rect 9470 2740 9547 2796
rect 9603 2740 9689 2796
rect 9745 2740 9810 2796
rect 9470 2654 9810 2740
rect 9470 2598 9547 2654
rect 9603 2598 9689 2654
rect 9745 2598 9810 2654
rect 9470 2512 9810 2598
rect 9470 2456 9547 2512
rect 9603 2456 9689 2512
rect 9745 2456 9810 2512
rect 9470 2370 9810 2456
rect 9470 2314 9547 2370
rect 9603 2314 9689 2370
rect 9745 2314 9810 2370
rect 9470 2228 9810 2314
rect 9470 2172 9547 2228
rect 9603 2172 9689 2228
rect 9745 2172 9810 2228
rect 9470 2086 9810 2172
rect 9470 2030 9547 2086
rect 9603 2030 9689 2086
rect 9745 2030 9810 2086
rect 9470 1944 9810 2030
rect 9470 1888 9547 1944
rect 9603 1888 9689 1944
rect 9745 1888 9810 1944
rect 9470 1802 9810 1888
rect 9470 1746 9547 1802
rect 9603 1746 9689 1802
rect 9745 1746 9810 1802
rect 9470 1660 9810 1746
rect 9470 1604 9547 1660
rect 9603 1604 9689 1660
rect 9745 1604 9810 1660
rect 9470 1518 9810 1604
rect 9470 1462 9547 1518
rect 9603 1462 9689 1518
rect 9745 1462 9810 1518
rect 9470 1376 9810 1462
rect 9470 1320 9547 1376
rect 9603 1320 9689 1376
rect 9745 1320 9810 1376
rect 9470 1234 9810 1320
rect 9470 1178 9547 1234
rect 9603 1178 9689 1234
rect 9745 1178 9810 1234
rect 9470 1092 9810 1178
rect 9470 1036 9547 1092
rect 9603 1036 9689 1092
rect 9745 1036 9810 1092
rect 9470 950 9810 1036
rect 9470 894 9547 950
rect 9603 894 9689 950
rect 9745 894 9810 950
rect 9470 808 9810 894
rect 9470 752 9547 808
rect 9603 752 9689 808
rect 9745 752 9810 808
rect 9470 666 9810 752
rect 9470 610 9547 666
rect 9603 610 9689 666
rect 9745 610 9810 666
rect 9470 524 9810 610
rect 9470 468 9547 524
rect 9603 468 9689 524
rect 9745 468 9810 524
rect 9470 400 9810 468
rect 10010 12310 10350 12400
rect 10010 12254 10081 12310
rect 10137 12254 10223 12310
rect 10279 12254 10350 12310
rect 10010 12168 10350 12254
rect 10010 12112 10081 12168
rect 10137 12112 10223 12168
rect 10279 12112 10350 12168
rect 10010 12026 10350 12112
rect 10010 11970 10081 12026
rect 10137 11970 10223 12026
rect 10279 11970 10350 12026
rect 10010 11884 10350 11970
rect 10010 11828 10081 11884
rect 10137 11828 10223 11884
rect 10279 11828 10350 11884
rect 10010 11742 10350 11828
rect 10010 11686 10081 11742
rect 10137 11686 10223 11742
rect 10279 11686 10350 11742
rect 10010 11600 10350 11686
rect 10010 11544 10081 11600
rect 10137 11544 10223 11600
rect 10279 11544 10350 11600
rect 10010 11458 10350 11544
rect 10010 11402 10081 11458
rect 10137 11402 10223 11458
rect 10279 11402 10350 11458
rect 10010 11316 10350 11402
rect 10010 11260 10081 11316
rect 10137 11260 10223 11316
rect 10279 11260 10350 11316
rect 10010 11174 10350 11260
rect 10010 11118 10081 11174
rect 10137 11118 10223 11174
rect 10279 11118 10350 11174
rect 10010 11032 10350 11118
rect 10010 10976 10081 11032
rect 10137 10976 10223 11032
rect 10279 10976 10350 11032
rect 10010 10890 10350 10976
rect 10010 10834 10081 10890
rect 10137 10834 10223 10890
rect 10279 10834 10350 10890
rect 10010 10748 10350 10834
rect 10010 10692 10081 10748
rect 10137 10692 10223 10748
rect 10279 10692 10350 10748
rect 10010 10606 10350 10692
rect 10010 10550 10081 10606
rect 10137 10550 10223 10606
rect 10279 10550 10350 10606
rect 10010 10464 10350 10550
rect 10010 10408 10081 10464
rect 10137 10408 10223 10464
rect 10279 10408 10350 10464
rect 10010 10322 10350 10408
rect 10010 10266 10081 10322
rect 10137 10266 10223 10322
rect 10279 10266 10350 10322
rect 10010 10180 10350 10266
rect 10010 10124 10081 10180
rect 10137 10124 10223 10180
rect 10279 10124 10350 10180
rect 10010 10038 10350 10124
rect 10010 9982 10081 10038
rect 10137 9982 10223 10038
rect 10279 9982 10350 10038
rect 10010 9896 10350 9982
rect 10010 9840 10081 9896
rect 10137 9840 10223 9896
rect 10279 9840 10350 9896
rect 10010 9754 10350 9840
rect 10010 9698 10081 9754
rect 10137 9698 10223 9754
rect 10279 9698 10350 9754
rect 10010 9612 10350 9698
rect 10010 9556 10081 9612
rect 10137 9556 10223 9612
rect 10279 9556 10350 9612
rect 10010 9470 10350 9556
rect 10010 9414 10081 9470
rect 10137 9414 10223 9470
rect 10279 9414 10350 9470
rect 10010 9328 10350 9414
rect 10010 9272 10081 9328
rect 10137 9272 10223 9328
rect 10279 9272 10350 9328
rect 10010 9186 10350 9272
rect 10010 9130 10081 9186
rect 10137 9130 10223 9186
rect 10279 9130 10350 9186
rect 10010 9044 10350 9130
rect 10010 8988 10081 9044
rect 10137 8988 10223 9044
rect 10279 8988 10350 9044
rect 10010 8902 10350 8988
rect 10010 8846 10081 8902
rect 10137 8846 10223 8902
rect 10279 8846 10350 8902
rect 10010 8760 10350 8846
rect 10010 8704 10081 8760
rect 10137 8704 10223 8760
rect 10279 8704 10350 8760
rect 10010 8618 10350 8704
rect 10010 8562 10081 8618
rect 10137 8562 10223 8618
rect 10279 8562 10350 8618
rect 10010 8476 10350 8562
rect 10010 8420 10081 8476
rect 10137 8420 10223 8476
rect 10279 8420 10350 8476
rect 10010 8334 10350 8420
rect 10010 8278 10081 8334
rect 10137 8278 10223 8334
rect 10279 8278 10350 8334
rect 10010 8192 10350 8278
rect 10010 8136 10081 8192
rect 10137 8136 10223 8192
rect 10279 8136 10350 8192
rect 10010 8050 10350 8136
rect 10010 7994 10081 8050
rect 10137 7994 10223 8050
rect 10279 7994 10350 8050
rect 10010 7908 10350 7994
rect 10010 7852 10081 7908
rect 10137 7852 10223 7908
rect 10279 7852 10350 7908
rect 10010 7766 10350 7852
rect 10010 7710 10081 7766
rect 10137 7710 10223 7766
rect 10279 7710 10350 7766
rect 10010 7624 10350 7710
rect 10010 7568 10081 7624
rect 10137 7568 10223 7624
rect 10279 7568 10350 7624
rect 10010 7482 10350 7568
rect 10010 7426 10081 7482
rect 10137 7426 10223 7482
rect 10279 7426 10350 7482
rect 10010 7340 10350 7426
rect 10010 7284 10081 7340
rect 10137 7284 10223 7340
rect 10279 7284 10350 7340
rect 10010 7198 10350 7284
rect 10010 7142 10081 7198
rect 10137 7142 10223 7198
rect 10279 7142 10350 7198
rect 10010 7056 10350 7142
rect 10010 7000 10081 7056
rect 10137 7000 10223 7056
rect 10279 7000 10350 7056
rect 10010 6914 10350 7000
rect 10010 6858 10081 6914
rect 10137 6858 10223 6914
rect 10279 6858 10350 6914
rect 10010 6772 10350 6858
rect 10010 6716 10081 6772
rect 10137 6716 10223 6772
rect 10279 6716 10350 6772
rect 10010 6630 10350 6716
rect 10010 6574 10081 6630
rect 10137 6574 10223 6630
rect 10279 6574 10350 6630
rect 10010 6488 10350 6574
rect 10010 6432 10081 6488
rect 10137 6432 10223 6488
rect 10279 6432 10350 6488
rect 10010 6346 10350 6432
rect 10010 6290 10081 6346
rect 10137 6290 10223 6346
rect 10279 6290 10350 6346
rect 10010 6204 10350 6290
rect 10010 6148 10081 6204
rect 10137 6148 10223 6204
rect 10279 6148 10350 6204
rect 10010 6062 10350 6148
rect 10010 6006 10081 6062
rect 10137 6006 10223 6062
rect 10279 6006 10350 6062
rect 10010 5920 10350 6006
rect 10010 5864 10081 5920
rect 10137 5864 10223 5920
rect 10279 5864 10350 5920
rect 10010 5778 10350 5864
rect 10010 5722 10081 5778
rect 10137 5722 10223 5778
rect 10279 5722 10350 5778
rect 10010 5636 10350 5722
rect 10010 5580 10081 5636
rect 10137 5580 10223 5636
rect 10279 5580 10350 5636
rect 10010 5494 10350 5580
rect 10010 5438 10081 5494
rect 10137 5438 10223 5494
rect 10279 5438 10350 5494
rect 10010 5352 10350 5438
rect 10010 5296 10081 5352
rect 10137 5296 10223 5352
rect 10279 5296 10350 5352
rect 10010 5210 10350 5296
rect 10010 5154 10081 5210
rect 10137 5154 10223 5210
rect 10279 5154 10350 5210
rect 10010 5068 10350 5154
rect 10010 5012 10081 5068
rect 10137 5012 10223 5068
rect 10279 5012 10350 5068
rect 10010 4926 10350 5012
rect 10010 4870 10081 4926
rect 10137 4870 10223 4926
rect 10279 4870 10350 4926
rect 10010 4784 10350 4870
rect 10010 4728 10081 4784
rect 10137 4728 10223 4784
rect 10279 4728 10350 4784
rect 10010 4642 10350 4728
rect 10010 4586 10081 4642
rect 10137 4586 10223 4642
rect 10279 4586 10350 4642
rect 10010 4500 10350 4586
rect 10010 4444 10081 4500
rect 10137 4444 10223 4500
rect 10279 4444 10350 4500
rect 10010 4358 10350 4444
rect 10010 4302 10081 4358
rect 10137 4302 10223 4358
rect 10279 4302 10350 4358
rect 10010 4216 10350 4302
rect 10010 4160 10081 4216
rect 10137 4160 10223 4216
rect 10279 4160 10350 4216
rect 10010 4074 10350 4160
rect 10010 4018 10081 4074
rect 10137 4018 10223 4074
rect 10279 4018 10350 4074
rect 10010 3932 10350 4018
rect 10010 3876 10081 3932
rect 10137 3876 10223 3932
rect 10279 3876 10350 3932
rect 10010 3790 10350 3876
rect 10010 3734 10081 3790
rect 10137 3734 10223 3790
rect 10279 3734 10350 3790
rect 10010 3648 10350 3734
rect 10010 3592 10081 3648
rect 10137 3592 10223 3648
rect 10279 3592 10350 3648
rect 10010 3506 10350 3592
rect 10010 3450 10081 3506
rect 10137 3450 10223 3506
rect 10279 3450 10350 3506
rect 10010 3364 10350 3450
rect 10010 3308 10081 3364
rect 10137 3308 10223 3364
rect 10279 3308 10350 3364
rect 10010 3222 10350 3308
rect 10010 3166 10081 3222
rect 10137 3166 10223 3222
rect 10279 3166 10350 3222
rect 10010 3080 10350 3166
rect 10010 3024 10081 3080
rect 10137 3024 10223 3080
rect 10279 3024 10350 3080
rect 10010 2938 10350 3024
rect 10010 2882 10081 2938
rect 10137 2882 10223 2938
rect 10279 2882 10350 2938
rect 10010 2796 10350 2882
rect 10010 2740 10081 2796
rect 10137 2740 10223 2796
rect 10279 2740 10350 2796
rect 10010 2654 10350 2740
rect 10010 2598 10081 2654
rect 10137 2598 10223 2654
rect 10279 2598 10350 2654
rect 10010 2512 10350 2598
rect 10010 2456 10081 2512
rect 10137 2456 10223 2512
rect 10279 2456 10350 2512
rect 10010 2370 10350 2456
rect 10010 2314 10081 2370
rect 10137 2314 10223 2370
rect 10279 2314 10350 2370
rect 10010 2228 10350 2314
rect 10010 2172 10081 2228
rect 10137 2172 10223 2228
rect 10279 2172 10350 2228
rect 10010 2086 10350 2172
rect 10010 2030 10081 2086
rect 10137 2030 10223 2086
rect 10279 2030 10350 2086
rect 10010 1944 10350 2030
rect 10010 1888 10081 1944
rect 10137 1888 10223 1944
rect 10279 1888 10350 1944
rect 10010 1802 10350 1888
rect 10010 1746 10081 1802
rect 10137 1746 10223 1802
rect 10279 1746 10350 1802
rect 10010 1660 10350 1746
rect 10010 1604 10081 1660
rect 10137 1604 10223 1660
rect 10279 1604 10350 1660
rect 10010 1518 10350 1604
rect 10010 1462 10081 1518
rect 10137 1462 10223 1518
rect 10279 1462 10350 1518
rect 10010 1376 10350 1462
rect 10010 1320 10081 1376
rect 10137 1320 10223 1376
rect 10279 1320 10350 1376
rect 10010 1234 10350 1320
rect 10010 1178 10081 1234
rect 10137 1178 10223 1234
rect 10279 1178 10350 1234
rect 10010 1092 10350 1178
rect 10010 1036 10081 1092
rect 10137 1036 10223 1092
rect 10279 1036 10350 1092
rect 10010 950 10350 1036
rect 10010 894 10081 950
rect 10137 894 10223 950
rect 10279 894 10350 950
rect 10010 808 10350 894
rect 10010 752 10081 808
rect 10137 752 10223 808
rect 10279 752 10350 808
rect 10010 666 10350 752
rect 10010 610 10081 666
rect 10137 610 10223 666
rect 10279 610 10350 666
rect 10010 524 10350 610
rect 10010 468 10081 524
rect 10137 468 10223 524
rect 10279 468 10350 524
rect 10010 400 10350 468
rect 10550 12310 10890 12400
rect 10550 12254 10622 12310
rect 10678 12254 10764 12310
rect 10820 12254 10890 12310
rect 10550 12168 10890 12254
rect 10550 12112 10622 12168
rect 10678 12112 10764 12168
rect 10820 12112 10890 12168
rect 10550 12026 10890 12112
rect 10550 11970 10622 12026
rect 10678 11970 10764 12026
rect 10820 11970 10890 12026
rect 10550 11884 10890 11970
rect 10550 11828 10622 11884
rect 10678 11828 10764 11884
rect 10820 11828 10890 11884
rect 10550 11742 10890 11828
rect 10550 11686 10622 11742
rect 10678 11686 10764 11742
rect 10820 11686 10890 11742
rect 10550 11600 10890 11686
rect 10550 11544 10622 11600
rect 10678 11544 10764 11600
rect 10820 11544 10890 11600
rect 10550 11458 10890 11544
rect 10550 11402 10622 11458
rect 10678 11402 10764 11458
rect 10820 11402 10890 11458
rect 10550 11316 10890 11402
rect 10550 11260 10622 11316
rect 10678 11260 10764 11316
rect 10820 11260 10890 11316
rect 10550 11174 10890 11260
rect 10550 11118 10622 11174
rect 10678 11118 10764 11174
rect 10820 11118 10890 11174
rect 10550 11032 10890 11118
rect 10550 10976 10622 11032
rect 10678 10976 10764 11032
rect 10820 10976 10890 11032
rect 10550 10890 10890 10976
rect 10550 10834 10622 10890
rect 10678 10834 10764 10890
rect 10820 10834 10890 10890
rect 10550 10748 10890 10834
rect 10550 10692 10622 10748
rect 10678 10692 10764 10748
rect 10820 10692 10890 10748
rect 10550 10606 10890 10692
rect 10550 10550 10622 10606
rect 10678 10550 10764 10606
rect 10820 10550 10890 10606
rect 10550 10464 10890 10550
rect 10550 10408 10622 10464
rect 10678 10408 10764 10464
rect 10820 10408 10890 10464
rect 10550 10322 10890 10408
rect 10550 10266 10622 10322
rect 10678 10266 10764 10322
rect 10820 10266 10890 10322
rect 10550 10180 10890 10266
rect 10550 10124 10622 10180
rect 10678 10124 10764 10180
rect 10820 10124 10890 10180
rect 10550 10038 10890 10124
rect 10550 9982 10622 10038
rect 10678 9982 10764 10038
rect 10820 9982 10890 10038
rect 10550 9896 10890 9982
rect 10550 9840 10622 9896
rect 10678 9840 10764 9896
rect 10820 9840 10890 9896
rect 10550 9754 10890 9840
rect 10550 9698 10622 9754
rect 10678 9698 10764 9754
rect 10820 9698 10890 9754
rect 10550 9612 10890 9698
rect 10550 9556 10622 9612
rect 10678 9556 10764 9612
rect 10820 9556 10890 9612
rect 10550 9470 10890 9556
rect 10550 9414 10622 9470
rect 10678 9414 10764 9470
rect 10820 9414 10890 9470
rect 10550 9328 10890 9414
rect 10550 9272 10622 9328
rect 10678 9272 10764 9328
rect 10820 9272 10890 9328
rect 10550 9186 10890 9272
rect 10550 9130 10622 9186
rect 10678 9130 10764 9186
rect 10820 9130 10890 9186
rect 10550 9044 10890 9130
rect 10550 8988 10622 9044
rect 10678 8988 10764 9044
rect 10820 8988 10890 9044
rect 10550 8902 10890 8988
rect 10550 8846 10622 8902
rect 10678 8846 10764 8902
rect 10820 8846 10890 8902
rect 10550 8760 10890 8846
rect 10550 8704 10622 8760
rect 10678 8704 10764 8760
rect 10820 8704 10890 8760
rect 10550 8618 10890 8704
rect 10550 8562 10622 8618
rect 10678 8562 10764 8618
rect 10820 8562 10890 8618
rect 10550 8476 10890 8562
rect 10550 8420 10622 8476
rect 10678 8420 10764 8476
rect 10820 8420 10890 8476
rect 10550 8334 10890 8420
rect 10550 8278 10622 8334
rect 10678 8278 10764 8334
rect 10820 8278 10890 8334
rect 10550 8192 10890 8278
rect 10550 8136 10622 8192
rect 10678 8136 10764 8192
rect 10820 8136 10890 8192
rect 10550 8050 10890 8136
rect 10550 7994 10622 8050
rect 10678 7994 10764 8050
rect 10820 7994 10890 8050
rect 10550 7908 10890 7994
rect 10550 7852 10622 7908
rect 10678 7852 10764 7908
rect 10820 7852 10890 7908
rect 10550 7766 10890 7852
rect 10550 7710 10622 7766
rect 10678 7710 10764 7766
rect 10820 7710 10890 7766
rect 10550 7624 10890 7710
rect 10550 7568 10622 7624
rect 10678 7568 10764 7624
rect 10820 7568 10890 7624
rect 10550 7482 10890 7568
rect 10550 7426 10622 7482
rect 10678 7426 10764 7482
rect 10820 7426 10890 7482
rect 10550 7340 10890 7426
rect 10550 7284 10622 7340
rect 10678 7284 10764 7340
rect 10820 7284 10890 7340
rect 10550 7198 10890 7284
rect 10550 7142 10622 7198
rect 10678 7142 10764 7198
rect 10820 7142 10890 7198
rect 10550 7056 10890 7142
rect 10550 7000 10622 7056
rect 10678 7000 10764 7056
rect 10820 7000 10890 7056
rect 10550 6914 10890 7000
rect 10550 6858 10622 6914
rect 10678 6858 10764 6914
rect 10820 6858 10890 6914
rect 10550 6772 10890 6858
rect 10550 6716 10622 6772
rect 10678 6716 10764 6772
rect 10820 6716 10890 6772
rect 10550 6630 10890 6716
rect 10550 6574 10622 6630
rect 10678 6574 10764 6630
rect 10820 6574 10890 6630
rect 10550 6488 10890 6574
rect 10550 6432 10622 6488
rect 10678 6432 10764 6488
rect 10820 6432 10890 6488
rect 10550 6346 10890 6432
rect 10550 6290 10622 6346
rect 10678 6290 10764 6346
rect 10820 6290 10890 6346
rect 10550 6204 10890 6290
rect 10550 6148 10622 6204
rect 10678 6148 10764 6204
rect 10820 6148 10890 6204
rect 10550 6062 10890 6148
rect 10550 6006 10622 6062
rect 10678 6006 10764 6062
rect 10820 6006 10890 6062
rect 10550 5920 10890 6006
rect 10550 5864 10622 5920
rect 10678 5864 10764 5920
rect 10820 5864 10890 5920
rect 10550 5778 10890 5864
rect 10550 5722 10622 5778
rect 10678 5722 10764 5778
rect 10820 5722 10890 5778
rect 10550 5636 10890 5722
rect 10550 5580 10622 5636
rect 10678 5580 10764 5636
rect 10820 5580 10890 5636
rect 10550 5494 10890 5580
rect 10550 5438 10622 5494
rect 10678 5438 10764 5494
rect 10820 5438 10890 5494
rect 10550 5352 10890 5438
rect 10550 5296 10622 5352
rect 10678 5296 10764 5352
rect 10820 5296 10890 5352
rect 10550 5210 10890 5296
rect 10550 5154 10622 5210
rect 10678 5154 10764 5210
rect 10820 5154 10890 5210
rect 10550 5068 10890 5154
rect 10550 5012 10622 5068
rect 10678 5012 10764 5068
rect 10820 5012 10890 5068
rect 10550 4926 10890 5012
rect 10550 4870 10622 4926
rect 10678 4870 10764 4926
rect 10820 4870 10890 4926
rect 10550 4784 10890 4870
rect 10550 4728 10622 4784
rect 10678 4728 10764 4784
rect 10820 4728 10890 4784
rect 10550 4642 10890 4728
rect 10550 4586 10622 4642
rect 10678 4586 10764 4642
rect 10820 4586 10890 4642
rect 10550 4500 10890 4586
rect 10550 4444 10622 4500
rect 10678 4444 10764 4500
rect 10820 4444 10890 4500
rect 10550 4358 10890 4444
rect 10550 4302 10622 4358
rect 10678 4302 10764 4358
rect 10820 4302 10890 4358
rect 10550 4216 10890 4302
rect 10550 4160 10622 4216
rect 10678 4160 10764 4216
rect 10820 4160 10890 4216
rect 10550 4074 10890 4160
rect 10550 4018 10622 4074
rect 10678 4018 10764 4074
rect 10820 4018 10890 4074
rect 10550 3932 10890 4018
rect 10550 3876 10622 3932
rect 10678 3876 10764 3932
rect 10820 3876 10890 3932
rect 10550 3790 10890 3876
rect 10550 3734 10622 3790
rect 10678 3734 10764 3790
rect 10820 3734 10890 3790
rect 10550 3648 10890 3734
rect 10550 3592 10622 3648
rect 10678 3592 10764 3648
rect 10820 3592 10890 3648
rect 10550 3506 10890 3592
rect 10550 3450 10622 3506
rect 10678 3450 10764 3506
rect 10820 3450 10890 3506
rect 10550 3364 10890 3450
rect 10550 3308 10622 3364
rect 10678 3308 10764 3364
rect 10820 3308 10890 3364
rect 10550 3222 10890 3308
rect 10550 3166 10622 3222
rect 10678 3166 10764 3222
rect 10820 3166 10890 3222
rect 10550 3080 10890 3166
rect 10550 3024 10622 3080
rect 10678 3024 10764 3080
rect 10820 3024 10890 3080
rect 10550 2938 10890 3024
rect 10550 2882 10622 2938
rect 10678 2882 10764 2938
rect 10820 2882 10890 2938
rect 10550 2796 10890 2882
rect 10550 2740 10622 2796
rect 10678 2740 10764 2796
rect 10820 2740 10890 2796
rect 10550 2654 10890 2740
rect 10550 2598 10622 2654
rect 10678 2598 10764 2654
rect 10820 2598 10890 2654
rect 10550 2512 10890 2598
rect 10550 2456 10622 2512
rect 10678 2456 10764 2512
rect 10820 2456 10890 2512
rect 10550 2370 10890 2456
rect 10550 2314 10622 2370
rect 10678 2314 10764 2370
rect 10820 2314 10890 2370
rect 10550 2228 10890 2314
rect 10550 2172 10622 2228
rect 10678 2172 10764 2228
rect 10820 2172 10890 2228
rect 10550 2086 10890 2172
rect 10550 2030 10622 2086
rect 10678 2030 10764 2086
rect 10820 2030 10890 2086
rect 10550 1944 10890 2030
rect 10550 1888 10622 1944
rect 10678 1888 10764 1944
rect 10820 1888 10890 1944
rect 10550 1802 10890 1888
rect 10550 1746 10622 1802
rect 10678 1746 10764 1802
rect 10820 1746 10890 1802
rect 10550 1660 10890 1746
rect 10550 1604 10622 1660
rect 10678 1604 10764 1660
rect 10820 1604 10890 1660
rect 10550 1518 10890 1604
rect 10550 1462 10622 1518
rect 10678 1462 10764 1518
rect 10820 1462 10890 1518
rect 10550 1376 10890 1462
rect 10550 1320 10622 1376
rect 10678 1320 10764 1376
rect 10820 1320 10890 1376
rect 10550 1234 10890 1320
rect 10550 1178 10622 1234
rect 10678 1178 10764 1234
rect 10820 1178 10890 1234
rect 10550 1092 10890 1178
rect 10550 1036 10622 1092
rect 10678 1036 10764 1092
rect 10820 1036 10890 1092
rect 10550 950 10890 1036
rect 10550 894 10622 950
rect 10678 894 10764 950
rect 10820 894 10890 950
rect 10550 808 10890 894
rect 10550 752 10622 808
rect 10678 752 10764 808
rect 10820 752 10890 808
rect 10550 666 10890 752
rect 10550 610 10622 666
rect 10678 610 10764 666
rect 10820 610 10890 666
rect 10550 524 10890 610
rect 10550 468 10622 524
rect 10678 468 10764 524
rect 10820 468 10890 524
rect 10550 400 10890 468
rect 11090 12310 11430 12400
rect 11090 12254 11162 12310
rect 11218 12254 11304 12310
rect 11360 12254 11430 12310
rect 11090 12168 11430 12254
rect 11090 12112 11162 12168
rect 11218 12112 11304 12168
rect 11360 12112 11430 12168
rect 11090 12026 11430 12112
rect 11090 11970 11162 12026
rect 11218 11970 11304 12026
rect 11360 11970 11430 12026
rect 11090 11884 11430 11970
rect 11090 11828 11162 11884
rect 11218 11828 11304 11884
rect 11360 11828 11430 11884
rect 11090 11742 11430 11828
rect 11090 11686 11162 11742
rect 11218 11686 11304 11742
rect 11360 11686 11430 11742
rect 11090 11600 11430 11686
rect 11090 11544 11162 11600
rect 11218 11544 11304 11600
rect 11360 11544 11430 11600
rect 11090 11458 11430 11544
rect 11090 11402 11162 11458
rect 11218 11402 11304 11458
rect 11360 11402 11430 11458
rect 11090 11316 11430 11402
rect 11090 11260 11162 11316
rect 11218 11260 11304 11316
rect 11360 11260 11430 11316
rect 11090 11174 11430 11260
rect 11090 11118 11162 11174
rect 11218 11118 11304 11174
rect 11360 11118 11430 11174
rect 11090 11032 11430 11118
rect 11090 10976 11162 11032
rect 11218 10976 11304 11032
rect 11360 10976 11430 11032
rect 11090 10890 11430 10976
rect 11090 10834 11162 10890
rect 11218 10834 11304 10890
rect 11360 10834 11430 10890
rect 11090 10748 11430 10834
rect 11090 10692 11162 10748
rect 11218 10692 11304 10748
rect 11360 10692 11430 10748
rect 11090 10606 11430 10692
rect 11090 10550 11162 10606
rect 11218 10550 11304 10606
rect 11360 10550 11430 10606
rect 11090 10464 11430 10550
rect 11090 10408 11162 10464
rect 11218 10408 11304 10464
rect 11360 10408 11430 10464
rect 11090 10322 11430 10408
rect 11090 10266 11162 10322
rect 11218 10266 11304 10322
rect 11360 10266 11430 10322
rect 11090 10180 11430 10266
rect 11090 10124 11162 10180
rect 11218 10124 11304 10180
rect 11360 10124 11430 10180
rect 11090 10038 11430 10124
rect 11090 9982 11162 10038
rect 11218 9982 11304 10038
rect 11360 9982 11430 10038
rect 11090 9896 11430 9982
rect 11090 9840 11162 9896
rect 11218 9840 11304 9896
rect 11360 9840 11430 9896
rect 11090 9754 11430 9840
rect 11090 9698 11162 9754
rect 11218 9698 11304 9754
rect 11360 9698 11430 9754
rect 11090 9612 11430 9698
rect 11090 9556 11162 9612
rect 11218 9556 11304 9612
rect 11360 9556 11430 9612
rect 11090 9470 11430 9556
rect 11090 9414 11162 9470
rect 11218 9414 11304 9470
rect 11360 9414 11430 9470
rect 11090 9328 11430 9414
rect 11090 9272 11162 9328
rect 11218 9272 11304 9328
rect 11360 9272 11430 9328
rect 11090 9186 11430 9272
rect 11090 9130 11162 9186
rect 11218 9130 11304 9186
rect 11360 9130 11430 9186
rect 11090 9044 11430 9130
rect 11090 8988 11162 9044
rect 11218 8988 11304 9044
rect 11360 8988 11430 9044
rect 11090 8902 11430 8988
rect 11090 8846 11162 8902
rect 11218 8846 11304 8902
rect 11360 8846 11430 8902
rect 11090 8760 11430 8846
rect 11090 8704 11162 8760
rect 11218 8704 11304 8760
rect 11360 8704 11430 8760
rect 11090 8618 11430 8704
rect 11090 8562 11162 8618
rect 11218 8562 11304 8618
rect 11360 8562 11430 8618
rect 11090 8476 11430 8562
rect 11090 8420 11162 8476
rect 11218 8420 11304 8476
rect 11360 8420 11430 8476
rect 11090 8334 11430 8420
rect 11090 8278 11162 8334
rect 11218 8278 11304 8334
rect 11360 8278 11430 8334
rect 11090 8192 11430 8278
rect 11090 8136 11162 8192
rect 11218 8136 11304 8192
rect 11360 8136 11430 8192
rect 11090 8050 11430 8136
rect 11090 7994 11162 8050
rect 11218 7994 11304 8050
rect 11360 7994 11430 8050
rect 11090 7908 11430 7994
rect 11090 7852 11162 7908
rect 11218 7852 11304 7908
rect 11360 7852 11430 7908
rect 11090 7766 11430 7852
rect 11090 7710 11162 7766
rect 11218 7710 11304 7766
rect 11360 7710 11430 7766
rect 11090 7624 11430 7710
rect 11090 7568 11162 7624
rect 11218 7568 11304 7624
rect 11360 7568 11430 7624
rect 11090 7482 11430 7568
rect 11090 7426 11162 7482
rect 11218 7426 11304 7482
rect 11360 7426 11430 7482
rect 11090 7340 11430 7426
rect 11090 7284 11162 7340
rect 11218 7284 11304 7340
rect 11360 7284 11430 7340
rect 11090 7198 11430 7284
rect 11090 7142 11162 7198
rect 11218 7142 11304 7198
rect 11360 7142 11430 7198
rect 11090 7056 11430 7142
rect 11090 7000 11162 7056
rect 11218 7000 11304 7056
rect 11360 7000 11430 7056
rect 11090 6914 11430 7000
rect 11090 6858 11162 6914
rect 11218 6858 11304 6914
rect 11360 6858 11430 6914
rect 11090 6772 11430 6858
rect 11090 6716 11162 6772
rect 11218 6716 11304 6772
rect 11360 6716 11430 6772
rect 11090 6630 11430 6716
rect 11090 6574 11162 6630
rect 11218 6574 11304 6630
rect 11360 6574 11430 6630
rect 11090 6488 11430 6574
rect 11090 6432 11162 6488
rect 11218 6432 11304 6488
rect 11360 6432 11430 6488
rect 11090 6346 11430 6432
rect 11090 6290 11162 6346
rect 11218 6290 11304 6346
rect 11360 6290 11430 6346
rect 11090 6204 11430 6290
rect 11090 6148 11162 6204
rect 11218 6148 11304 6204
rect 11360 6148 11430 6204
rect 11090 6062 11430 6148
rect 11090 6006 11162 6062
rect 11218 6006 11304 6062
rect 11360 6006 11430 6062
rect 11090 5920 11430 6006
rect 11090 5864 11162 5920
rect 11218 5864 11304 5920
rect 11360 5864 11430 5920
rect 11090 5778 11430 5864
rect 11090 5722 11162 5778
rect 11218 5722 11304 5778
rect 11360 5722 11430 5778
rect 11090 5636 11430 5722
rect 11090 5580 11162 5636
rect 11218 5580 11304 5636
rect 11360 5580 11430 5636
rect 11090 5494 11430 5580
rect 11090 5438 11162 5494
rect 11218 5438 11304 5494
rect 11360 5438 11430 5494
rect 11090 5352 11430 5438
rect 11090 5296 11162 5352
rect 11218 5296 11304 5352
rect 11360 5296 11430 5352
rect 11090 5210 11430 5296
rect 11090 5154 11162 5210
rect 11218 5154 11304 5210
rect 11360 5154 11430 5210
rect 11090 5068 11430 5154
rect 11090 5012 11162 5068
rect 11218 5012 11304 5068
rect 11360 5012 11430 5068
rect 11090 4926 11430 5012
rect 11090 4870 11162 4926
rect 11218 4870 11304 4926
rect 11360 4870 11430 4926
rect 11090 4784 11430 4870
rect 11090 4728 11162 4784
rect 11218 4728 11304 4784
rect 11360 4728 11430 4784
rect 11090 4642 11430 4728
rect 11090 4586 11162 4642
rect 11218 4586 11304 4642
rect 11360 4586 11430 4642
rect 11090 4500 11430 4586
rect 11090 4444 11162 4500
rect 11218 4444 11304 4500
rect 11360 4444 11430 4500
rect 11090 4358 11430 4444
rect 11090 4302 11162 4358
rect 11218 4302 11304 4358
rect 11360 4302 11430 4358
rect 11090 4216 11430 4302
rect 11090 4160 11162 4216
rect 11218 4160 11304 4216
rect 11360 4160 11430 4216
rect 11090 4074 11430 4160
rect 11090 4018 11162 4074
rect 11218 4018 11304 4074
rect 11360 4018 11430 4074
rect 11090 3932 11430 4018
rect 11090 3876 11162 3932
rect 11218 3876 11304 3932
rect 11360 3876 11430 3932
rect 11090 3790 11430 3876
rect 11090 3734 11162 3790
rect 11218 3734 11304 3790
rect 11360 3734 11430 3790
rect 11090 3648 11430 3734
rect 11090 3592 11162 3648
rect 11218 3592 11304 3648
rect 11360 3592 11430 3648
rect 11090 3506 11430 3592
rect 11090 3450 11162 3506
rect 11218 3450 11304 3506
rect 11360 3450 11430 3506
rect 11090 3364 11430 3450
rect 11090 3308 11162 3364
rect 11218 3308 11304 3364
rect 11360 3308 11430 3364
rect 11090 3222 11430 3308
rect 11090 3166 11162 3222
rect 11218 3166 11304 3222
rect 11360 3166 11430 3222
rect 11090 3080 11430 3166
rect 11090 3024 11162 3080
rect 11218 3024 11304 3080
rect 11360 3024 11430 3080
rect 11090 2938 11430 3024
rect 11090 2882 11162 2938
rect 11218 2882 11304 2938
rect 11360 2882 11430 2938
rect 11090 2796 11430 2882
rect 11090 2740 11162 2796
rect 11218 2740 11304 2796
rect 11360 2740 11430 2796
rect 11090 2654 11430 2740
rect 11090 2598 11162 2654
rect 11218 2598 11304 2654
rect 11360 2598 11430 2654
rect 11090 2512 11430 2598
rect 11090 2456 11162 2512
rect 11218 2456 11304 2512
rect 11360 2456 11430 2512
rect 11090 2370 11430 2456
rect 11090 2314 11162 2370
rect 11218 2314 11304 2370
rect 11360 2314 11430 2370
rect 11090 2228 11430 2314
rect 11090 2172 11162 2228
rect 11218 2172 11304 2228
rect 11360 2172 11430 2228
rect 11090 2086 11430 2172
rect 11090 2030 11162 2086
rect 11218 2030 11304 2086
rect 11360 2030 11430 2086
rect 11090 1944 11430 2030
rect 11090 1888 11162 1944
rect 11218 1888 11304 1944
rect 11360 1888 11430 1944
rect 11090 1802 11430 1888
rect 11090 1746 11162 1802
rect 11218 1746 11304 1802
rect 11360 1746 11430 1802
rect 11090 1660 11430 1746
rect 11090 1604 11162 1660
rect 11218 1604 11304 1660
rect 11360 1604 11430 1660
rect 11090 1518 11430 1604
rect 11090 1462 11162 1518
rect 11218 1462 11304 1518
rect 11360 1462 11430 1518
rect 11090 1376 11430 1462
rect 11090 1320 11162 1376
rect 11218 1320 11304 1376
rect 11360 1320 11430 1376
rect 11090 1234 11430 1320
rect 11090 1178 11162 1234
rect 11218 1178 11304 1234
rect 11360 1178 11430 1234
rect 11090 1092 11430 1178
rect 11090 1036 11162 1092
rect 11218 1036 11304 1092
rect 11360 1036 11430 1092
rect 11090 950 11430 1036
rect 11090 894 11162 950
rect 11218 894 11304 950
rect 11360 894 11430 950
rect 11090 808 11430 894
rect 11090 752 11162 808
rect 11218 752 11304 808
rect 11360 752 11430 808
rect 11090 666 11430 752
rect 11090 610 11162 666
rect 11218 610 11304 666
rect 11360 610 11430 666
rect 11090 524 11430 610
rect 11090 468 11162 524
rect 11218 468 11304 524
rect 11360 468 11430 524
rect 11090 400 11430 468
rect 11630 12310 11970 12400
rect 11630 12254 11702 12310
rect 11758 12254 11844 12310
rect 11900 12254 11970 12310
rect 11630 12168 11970 12254
rect 11630 12112 11702 12168
rect 11758 12112 11844 12168
rect 11900 12112 11970 12168
rect 11630 12026 11970 12112
rect 11630 11970 11702 12026
rect 11758 11970 11844 12026
rect 11900 11970 11970 12026
rect 11630 11884 11970 11970
rect 11630 11828 11702 11884
rect 11758 11828 11844 11884
rect 11900 11828 11970 11884
rect 11630 11742 11970 11828
rect 11630 11686 11702 11742
rect 11758 11686 11844 11742
rect 11900 11686 11970 11742
rect 11630 11600 11970 11686
rect 11630 11544 11702 11600
rect 11758 11544 11844 11600
rect 11900 11544 11970 11600
rect 11630 11458 11970 11544
rect 11630 11402 11702 11458
rect 11758 11402 11844 11458
rect 11900 11402 11970 11458
rect 11630 11316 11970 11402
rect 11630 11260 11702 11316
rect 11758 11260 11844 11316
rect 11900 11260 11970 11316
rect 11630 11174 11970 11260
rect 11630 11118 11702 11174
rect 11758 11118 11844 11174
rect 11900 11118 11970 11174
rect 11630 11032 11970 11118
rect 11630 10976 11702 11032
rect 11758 10976 11844 11032
rect 11900 10976 11970 11032
rect 11630 10890 11970 10976
rect 11630 10834 11702 10890
rect 11758 10834 11844 10890
rect 11900 10834 11970 10890
rect 11630 10748 11970 10834
rect 11630 10692 11702 10748
rect 11758 10692 11844 10748
rect 11900 10692 11970 10748
rect 11630 10606 11970 10692
rect 11630 10550 11702 10606
rect 11758 10550 11844 10606
rect 11900 10550 11970 10606
rect 11630 10464 11970 10550
rect 11630 10408 11702 10464
rect 11758 10408 11844 10464
rect 11900 10408 11970 10464
rect 11630 10322 11970 10408
rect 11630 10266 11702 10322
rect 11758 10266 11844 10322
rect 11900 10266 11970 10322
rect 11630 10180 11970 10266
rect 11630 10124 11702 10180
rect 11758 10124 11844 10180
rect 11900 10124 11970 10180
rect 11630 10038 11970 10124
rect 11630 9982 11702 10038
rect 11758 9982 11844 10038
rect 11900 9982 11970 10038
rect 11630 9896 11970 9982
rect 11630 9840 11702 9896
rect 11758 9840 11844 9896
rect 11900 9840 11970 9896
rect 11630 9754 11970 9840
rect 11630 9698 11702 9754
rect 11758 9698 11844 9754
rect 11900 9698 11970 9754
rect 11630 9612 11970 9698
rect 11630 9556 11702 9612
rect 11758 9556 11844 9612
rect 11900 9556 11970 9612
rect 11630 9470 11970 9556
rect 11630 9414 11702 9470
rect 11758 9414 11844 9470
rect 11900 9414 11970 9470
rect 11630 9328 11970 9414
rect 11630 9272 11702 9328
rect 11758 9272 11844 9328
rect 11900 9272 11970 9328
rect 11630 9186 11970 9272
rect 11630 9130 11702 9186
rect 11758 9130 11844 9186
rect 11900 9130 11970 9186
rect 11630 9044 11970 9130
rect 11630 8988 11702 9044
rect 11758 8988 11844 9044
rect 11900 8988 11970 9044
rect 11630 8902 11970 8988
rect 11630 8846 11702 8902
rect 11758 8846 11844 8902
rect 11900 8846 11970 8902
rect 11630 8760 11970 8846
rect 11630 8704 11702 8760
rect 11758 8704 11844 8760
rect 11900 8704 11970 8760
rect 11630 8618 11970 8704
rect 11630 8562 11702 8618
rect 11758 8562 11844 8618
rect 11900 8562 11970 8618
rect 11630 8476 11970 8562
rect 11630 8420 11702 8476
rect 11758 8420 11844 8476
rect 11900 8420 11970 8476
rect 11630 8334 11970 8420
rect 11630 8278 11702 8334
rect 11758 8278 11844 8334
rect 11900 8278 11970 8334
rect 11630 8192 11970 8278
rect 11630 8136 11702 8192
rect 11758 8136 11844 8192
rect 11900 8136 11970 8192
rect 11630 8050 11970 8136
rect 11630 7994 11702 8050
rect 11758 7994 11844 8050
rect 11900 7994 11970 8050
rect 11630 7908 11970 7994
rect 11630 7852 11702 7908
rect 11758 7852 11844 7908
rect 11900 7852 11970 7908
rect 11630 7766 11970 7852
rect 11630 7710 11702 7766
rect 11758 7710 11844 7766
rect 11900 7710 11970 7766
rect 11630 7624 11970 7710
rect 11630 7568 11702 7624
rect 11758 7568 11844 7624
rect 11900 7568 11970 7624
rect 11630 7482 11970 7568
rect 11630 7426 11702 7482
rect 11758 7426 11844 7482
rect 11900 7426 11970 7482
rect 11630 7340 11970 7426
rect 11630 7284 11702 7340
rect 11758 7284 11844 7340
rect 11900 7284 11970 7340
rect 11630 7198 11970 7284
rect 11630 7142 11702 7198
rect 11758 7142 11844 7198
rect 11900 7142 11970 7198
rect 11630 7056 11970 7142
rect 11630 7000 11702 7056
rect 11758 7000 11844 7056
rect 11900 7000 11970 7056
rect 11630 6914 11970 7000
rect 11630 6858 11702 6914
rect 11758 6858 11844 6914
rect 11900 6858 11970 6914
rect 11630 6772 11970 6858
rect 11630 6716 11702 6772
rect 11758 6716 11844 6772
rect 11900 6716 11970 6772
rect 11630 6630 11970 6716
rect 11630 6574 11702 6630
rect 11758 6574 11844 6630
rect 11900 6574 11970 6630
rect 11630 6488 11970 6574
rect 11630 6432 11702 6488
rect 11758 6432 11844 6488
rect 11900 6432 11970 6488
rect 11630 6346 11970 6432
rect 11630 6290 11702 6346
rect 11758 6290 11844 6346
rect 11900 6290 11970 6346
rect 11630 6204 11970 6290
rect 11630 6148 11702 6204
rect 11758 6148 11844 6204
rect 11900 6148 11970 6204
rect 11630 6062 11970 6148
rect 11630 6006 11702 6062
rect 11758 6006 11844 6062
rect 11900 6006 11970 6062
rect 11630 5920 11970 6006
rect 11630 5864 11702 5920
rect 11758 5864 11844 5920
rect 11900 5864 11970 5920
rect 11630 5778 11970 5864
rect 11630 5722 11702 5778
rect 11758 5722 11844 5778
rect 11900 5722 11970 5778
rect 11630 5636 11970 5722
rect 11630 5580 11702 5636
rect 11758 5580 11844 5636
rect 11900 5580 11970 5636
rect 11630 5494 11970 5580
rect 11630 5438 11702 5494
rect 11758 5438 11844 5494
rect 11900 5438 11970 5494
rect 11630 5352 11970 5438
rect 11630 5296 11702 5352
rect 11758 5296 11844 5352
rect 11900 5296 11970 5352
rect 11630 5210 11970 5296
rect 11630 5154 11702 5210
rect 11758 5154 11844 5210
rect 11900 5154 11970 5210
rect 11630 5068 11970 5154
rect 11630 5012 11702 5068
rect 11758 5012 11844 5068
rect 11900 5012 11970 5068
rect 11630 4926 11970 5012
rect 11630 4870 11702 4926
rect 11758 4870 11844 4926
rect 11900 4870 11970 4926
rect 11630 4784 11970 4870
rect 11630 4728 11702 4784
rect 11758 4728 11844 4784
rect 11900 4728 11970 4784
rect 11630 4642 11970 4728
rect 11630 4586 11702 4642
rect 11758 4586 11844 4642
rect 11900 4586 11970 4642
rect 11630 4500 11970 4586
rect 11630 4444 11702 4500
rect 11758 4444 11844 4500
rect 11900 4444 11970 4500
rect 11630 4358 11970 4444
rect 11630 4302 11702 4358
rect 11758 4302 11844 4358
rect 11900 4302 11970 4358
rect 11630 4216 11970 4302
rect 11630 4160 11702 4216
rect 11758 4160 11844 4216
rect 11900 4160 11970 4216
rect 11630 4074 11970 4160
rect 11630 4018 11702 4074
rect 11758 4018 11844 4074
rect 11900 4018 11970 4074
rect 11630 3932 11970 4018
rect 11630 3876 11702 3932
rect 11758 3876 11844 3932
rect 11900 3876 11970 3932
rect 11630 3790 11970 3876
rect 11630 3734 11702 3790
rect 11758 3734 11844 3790
rect 11900 3734 11970 3790
rect 11630 3648 11970 3734
rect 11630 3592 11702 3648
rect 11758 3592 11844 3648
rect 11900 3592 11970 3648
rect 11630 3506 11970 3592
rect 11630 3450 11702 3506
rect 11758 3450 11844 3506
rect 11900 3450 11970 3506
rect 11630 3364 11970 3450
rect 11630 3308 11702 3364
rect 11758 3308 11844 3364
rect 11900 3308 11970 3364
rect 11630 3222 11970 3308
rect 11630 3166 11702 3222
rect 11758 3166 11844 3222
rect 11900 3166 11970 3222
rect 11630 3080 11970 3166
rect 11630 3024 11702 3080
rect 11758 3024 11844 3080
rect 11900 3024 11970 3080
rect 11630 2938 11970 3024
rect 11630 2882 11702 2938
rect 11758 2882 11844 2938
rect 11900 2882 11970 2938
rect 11630 2796 11970 2882
rect 11630 2740 11702 2796
rect 11758 2740 11844 2796
rect 11900 2740 11970 2796
rect 11630 2654 11970 2740
rect 11630 2598 11702 2654
rect 11758 2598 11844 2654
rect 11900 2598 11970 2654
rect 11630 2512 11970 2598
rect 11630 2456 11702 2512
rect 11758 2456 11844 2512
rect 11900 2456 11970 2512
rect 11630 2370 11970 2456
rect 11630 2314 11702 2370
rect 11758 2314 11844 2370
rect 11900 2314 11970 2370
rect 11630 2228 11970 2314
rect 11630 2172 11702 2228
rect 11758 2172 11844 2228
rect 11900 2172 11970 2228
rect 11630 2086 11970 2172
rect 11630 2030 11702 2086
rect 11758 2030 11844 2086
rect 11900 2030 11970 2086
rect 11630 1944 11970 2030
rect 11630 1888 11702 1944
rect 11758 1888 11844 1944
rect 11900 1888 11970 1944
rect 11630 1802 11970 1888
rect 11630 1746 11702 1802
rect 11758 1746 11844 1802
rect 11900 1746 11970 1802
rect 11630 1660 11970 1746
rect 11630 1604 11702 1660
rect 11758 1604 11844 1660
rect 11900 1604 11970 1660
rect 11630 1518 11970 1604
rect 11630 1462 11702 1518
rect 11758 1462 11844 1518
rect 11900 1462 11970 1518
rect 11630 1376 11970 1462
rect 11630 1320 11702 1376
rect 11758 1320 11844 1376
rect 11900 1320 11970 1376
rect 11630 1234 11970 1320
rect 11630 1178 11702 1234
rect 11758 1178 11844 1234
rect 11900 1178 11970 1234
rect 11630 1092 11970 1178
rect 11630 1036 11702 1092
rect 11758 1036 11844 1092
rect 11900 1036 11970 1092
rect 11630 950 11970 1036
rect 11630 894 11702 950
rect 11758 894 11844 950
rect 11900 894 11970 950
rect 11630 808 11970 894
rect 11630 752 11702 808
rect 11758 752 11844 808
rect 11900 752 11970 808
rect 11630 666 11970 752
rect 11630 610 11702 666
rect 11758 610 11844 666
rect 11900 610 11970 666
rect 11630 524 11970 610
rect 11630 468 11702 524
rect 11758 468 11844 524
rect 11900 468 11970 524
rect 11630 400 11970 468
rect 12400 12358 13200 12400
rect 12400 12302 12526 12358
rect 12582 12302 12650 12358
rect 12706 12302 12774 12358
rect 12830 12302 12898 12358
rect 12954 12302 13022 12358
rect 13078 12302 13200 12358
rect 12400 12234 13200 12302
rect 12400 12178 12526 12234
rect 12582 12178 12650 12234
rect 12706 12178 12774 12234
rect 12830 12178 12898 12234
rect 12954 12178 13022 12234
rect 13078 12178 13200 12234
rect 12400 12110 13200 12178
rect 12400 12054 12526 12110
rect 12582 12054 12650 12110
rect 12706 12054 12774 12110
rect 12830 12054 12898 12110
rect 12954 12054 13022 12110
rect 13078 12054 13200 12110
rect 12400 11986 13200 12054
rect 12400 11930 12526 11986
rect 12582 11930 12650 11986
rect 12706 11930 12774 11986
rect 12830 11930 12898 11986
rect 12954 11930 13022 11986
rect 13078 11930 13200 11986
rect 12400 11862 13200 11930
rect 12400 11806 12526 11862
rect 12582 11806 12650 11862
rect 12706 11806 12774 11862
rect 12830 11806 12898 11862
rect 12954 11806 13022 11862
rect 13078 11806 13200 11862
rect 12400 11738 13200 11806
rect 12400 11682 12526 11738
rect 12582 11682 12650 11738
rect 12706 11682 12774 11738
rect 12830 11682 12898 11738
rect 12954 11682 13022 11738
rect 13078 11682 13200 11738
rect 12400 11614 13200 11682
rect 12400 11558 12526 11614
rect 12582 11558 12650 11614
rect 12706 11558 12774 11614
rect 12830 11558 12898 11614
rect 12954 11558 13022 11614
rect 13078 11558 13200 11614
rect 12400 11490 13200 11558
rect 12400 11434 12526 11490
rect 12582 11434 12650 11490
rect 12706 11434 12774 11490
rect 12830 11434 12898 11490
rect 12954 11434 13022 11490
rect 13078 11434 13200 11490
rect 12400 11366 13200 11434
rect 12400 11310 12526 11366
rect 12582 11310 12650 11366
rect 12706 11310 12774 11366
rect 12830 11310 12898 11366
rect 12954 11310 13022 11366
rect 13078 11310 13200 11366
rect 12400 11242 13200 11310
rect 12400 11186 12526 11242
rect 12582 11186 12650 11242
rect 12706 11186 12774 11242
rect 12830 11186 12898 11242
rect 12954 11186 13022 11242
rect 13078 11186 13200 11242
rect 12400 11118 13200 11186
rect 12400 11062 12526 11118
rect 12582 11062 12650 11118
rect 12706 11062 12774 11118
rect 12830 11062 12898 11118
rect 12954 11062 13022 11118
rect 13078 11062 13200 11118
rect 12400 10994 13200 11062
rect 12400 10938 12526 10994
rect 12582 10938 12650 10994
rect 12706 10938 12774 10994
rect 12830 10938 12898 10994
rect 12954 10938 13022 10994
rect 13078 10938 13200 10994
rect 12400 10870 13200 10938
rect 12400 10814 12526 10870
rect 12582 10814 12650 10870
rect 12706 10814 12774 10870
rect 12830 10814 12898 10870
rect 12954 10814 13022 10870
rect 13078 10814 13200 10870
rect 12400 10746 13200 10814
rect 12400 10690 12526 10746
rect 12582 10690 12650 10746
rect 12706 10690 12774 10746
rect 12830 10690 12898 10746
rect 12954 10690 13022 10746
rect 13078 10690 13200 10746
rect 12400 10622 13200 10690
rect 12400 10566 12526 10622
rect 12582 10566 12650 10622
rect 12706 10566 12774 10622
rect 12830 10566 12898 10622
rect 12954 10566 13022 10622
rect 13078 10566 13200 10622
rect 12400 10498 13200 10566
rect 12400 10442 12526 10498
rect 12582 10442 12650 10498
rect 12706 10442 12774 10498
rect 12830 10442 12898 10498
rect 12954 10442 13022 10498
rect 13078 10442 13200 10498
rect 12400 10374 13200 10442
rect 12400 10318 12526 10374
rect 12582 10318 12650 10374
rect 12706 10318 12774 10374
rect 12830 10318 12898 10374
rect 12954 10318 13022 10374
rect 13078 10318 13200 10374
rect 12400 10250 13200 10318
rect 12400 10194 12526 10250
rect 12582 10194 12650 10250
rect 12706 10194 12774 10250
rect 12830 10194 12898 10250
rect 12954 10194 13022 10250
rect 13078 10194 13200 10250
rect 12400 10126 13200 10194
rect 12400 10070 12526 10126
rect 12582 10070 12650 10126
rect 12706 10070 12774 10126
rect 12830 10070 12898 10126
rect 12954 10070 13022 10126
rect 13078 10070 13200 10126
rect 12400 10002 13200 10070
rect 12400 9946 12526 10002
rect 12582 9946 12650 10002
rect 12706 9946 12774 10002
rect 12830 9946 12898 10002
rect 12954 9946 13022 10002
rect 13078 9946 13200 10002
rect 12400 9878 13200 9946
rect 12400 9822 12526 9878
rect 12582 9822 12650 9878
rect 12706 9822 12774 9878
rect 12830 9822 12898 9878
rect 12954 9822 13022 9878
rect 13078 9822 13200 9878
rect 12400 9754 13200 9822
rect 12400 9698 12526 9754
rect 12582 9698 12650 9754
rect 12706 9698 12774 9754
rect 12830 9698 12898 9754
rect 12954 9698 13022 9754
rect 13078 9698 13200 9754
rect 12400 9630 13200 9698
rect 12400 9574 12526 9630
rect 12582 9574 12650 9630
rect 12706 9574 12774 9630
rect 12830 9574 12898 9630
rect 12954 9574 13022 9630
rect 13078 9574 13200 9630
rect 12400 9506 13200 9574
rect 12400 9450 12526 9506
rect 12582 9450 12650 9506
rect 12706 9450 12774 9506
rect 12830 9450 12898 9506
rect 12954 9450 13022 9506
rect 13078 9450 13200 9506
rect 12400 9382 13200 9450
rect 12400 9326 12526 9382
rect 12582 9326 12650 9382
rect 12706 9326 12774 9382
rect 12830 9326 12898 9382
rect 12954 9326 13022 9382
rect 13078 9326 13200 9382
rect 12400 9258 13200 9326
rect 12400 9202 12526 9258
rect 12582 9202 12650 9258
rect 12706 9202 12774 9258
rect 12830 9202 12898 9258
rect 12954 9202 13022 9258
rect 13078 9202 13200 9258
rect 12400 9134 13200 9202
rect 12400 9078 12526 9134
rect 12582 9078 12650 9134
rect 12706 9078 12774 9134
rect 12830 9078 12898 9134
rect 12954 9078 13022 9134
rect 13078 9078 13200 9134
rect 12400 9010 13200 9078
rect 12400 8954 12526 9010
rect 12582 8954 12650 9010
rect 12706 8954 12774 9010
rect 12830 8954 12898 9010
rect 12954 8954 13022 9010
rect 13078 8954 13200 9010
rect 12400 8886 13200 8954
rect 12400 8830 12526 8886
rect 12582 8830 12650 8886
rect 12706 8830 12774 8886
rect 12830 8830 12898 8886
rect 12954 8830 13022 8886
rect 13078 8830 13200 8886
rect 12400 8762 13200 8830
rect 12400 8706 12526 8762
rect 12582 8706 12650 8762
rect 12706 8706 12774 8762
rect 12830 8706 12898 8762
rect 12954 8706 13022 8762
rect 13078 8706 13200 8762
rect 12400 8638 13200 8706
rect 12400 8582 12526 8638
rect 12582 8582 12650 8638
rect 12706 8582 12774 8638
rect 12830 8582 12898 8638
rect 12954 8582 13022 8638
rect 13078 8582 13200 8638
rect 12400 8514 13200 8582
rect 12400 8458 12526 8514
rect 12582 8458 12650 8514
rect 12706 8458 12774 8514
rect 12830 8458 12898 8514
rect 12954 8458 13022 8514
rect 13078 8458 13200 8514
rect 12400 8390 13200 8458
rect 12400 8334 12526 8390
rect 12582 8334 12650 8390
rect 12706 8334 12774 8390
rect 12830 8334 12898 8390
rect 12954 8334 13022 8390
rect 13078 8334 13200 8390
rect 12400 8266 13200 8334
rect 12400 8210 12526 8266
rect 12582 8210 12650 8266
rect 12706 8210 12774 8266
rect 12830 8210 12898 8266
rect 12954 8210 13022 8266
rect 13078 8210 13200 8266
rect 12400 8142 13200 8210
rect 12400 8086 12526 8142
rect 12582 8086 12650 8142
rect 12706 8086 12774 8142
rect 12830 8086 12898 8142
rect 12954 8086 13022 8142
rect 13078 8086 13200 8142
rect 12400 8018 13200 8086
rect 12400 7962 12526 8018
rect 12582 7962 12650 8018
rect 12706 7962 12774 8018
rect 12830 7962 12898 8018
rect 12954 7962 13022 8018
rect 13078 7962 13200 8018
rect 12400 7894 13200 7962
rect 12400 7838 12526 7894
rect 12582 7838 12650 7894
rect 12706 7838 12774 7894
rect 12830 7838 12898 7894
rect 12954 7838 13022 7894
rect 13078 7838 13200 7894
rect 12400 7770 13200 7838
rect 12400 7714 12526 7770
rect 12582 7714 12650 7770
rect 12706 7714 12774 7770
rect 12830 7714 12898 7770
rect 12954 7714 13022 7770
rect 13078 7714 13200 7770
rect 12400 7646 13200 7714
rect 12400 7590 12526 7646
rect 12582 7590 12650 7646
rect 12706 7590 12774 7646
rect 12830 7590 12898 7646
rect 12954 7590 13022 7646
rect 13078 7590 13200 7646
rect 12400 7522 13200 7590
rect 12400 7466 12526 7522
rect 12582 7466 12650 7522
rect 12706 7466 12774 7522
rect 12830 7466 12898 7522
rect 12954 7466 13022 7522
rect 13078 7466 13200 7522
rect 12400 7398 13200 7466
rect 12400 7342 12526 7398
rect 12582 7342 12650 7398
rect 12706 7342 12774 7398
rect 12830 7342 12898 7398
rect 12954 7342 13022 7398
rect 13078 7342 13200 7398
rect 12400 7274 13200 7342
rect 12400 7218 12526 7274
rect 12582 7218 12650 7274
rect 12706 7218 12774 7274
rect 12830 7218 12898 7274
rect 12954 7218 13022 7274
rect 13078 7218 13200 7274
rect 12400 7150 13200 7218
rect 12400 7094 12526 7150
rect 12582 7094 12650 7150
rect 12706 7094 12774 7150
rect 12830 7094 12898 7150
rect 12954 7094 13022 7150
rect 13078 7094 13200 7150
rect 12400 7026 13200 7094
rect 12400 6970 12526 7026
rect 12582 6970 12650 7026
rect 12706 6970 12774 7026
rect 12830 6970 12898 7026
rect 12954 6970 13022 7026
rect 13078 6970 13200 7026
rect 12400 6902 13200 6970
rect 12400 6846 12526 6902
rect 12582 6846 12650 6902
rect 12706 6846 12774 6902
rect 12830 6846 12898 6902
rect 12954 6846 13022 6902
rect 13078 6846 13200 6902
rect 12400 6778 13200 6846
rect 12400 6722 12526 6778
rect 12582 6722 12650 6778
rect 12706 6722 12774 6778
rect 12830 6722 12898 6778
rect 12954 6722 13022 6778
rect 13078 6722 13200 6778
rect 12400 6654 13200 6722
rect 12400 6598 12526 6654
rect 12582 6598 12650 6654
rect 12706 6598 12774 6654
rect 12830 6598 12898 6654
rect 12954 6598 13022 6654
rect 13078 6598 13200 6654
rect 12400 6530 13200 6598
rect 12400 6474 12526 6530
rect 12582 6474 12650 6530
rect 12706 6474 12774 6530
rect 12830 6474 12898 6530
rect 12954 6474 13022 6530
rect 13078 6474 13200 6530
rect 12400 6406 13200 6474
rect 12400 6350 12526 6406
rect 12582 6350 12650 6406
rect 12706 6350 12774 6406
rect 12830 6350 12898 6406
rect 12954 6350 13022 6406
rect 13078 6350 13200 6406
rect 12400 6282 13200 6350
rect 12400 6226 12526 6282
rect 12582 6226 12650 6282
rect 12706 6226 12774 6282
rect 12830 6226 12898 6282
rect 12954 6226 13022 6282
rect 13078 6226 13200 6282
rect 12400 6158 13200 6226
rect 12400 6102 12526 6158
rect 12582 6102 12650 6158
rect 12706 6102 12774 6158
rect 12830 6102 12898 6158
rect 12954 6102 13022 6158
rect 13078 6102 13200 6158
rect 12400 6034 13200 6102
rect 12400 5978 12526 6034
rect 12582 5978 12650 6034
rect 12706 5978 12774 6034
rect 12830 5978 12898 6034
rect 12954 5978 13022 6034
rect 13078 5978 13200 6034
rect 12400 5910 13200 5978
rect 12400 5854 12526 5910
rect 12582 5854 12650 5910
rect 12706 5854 12774 5910
rect 12830 5854 12898 5910
rect 12954 5854 13022 5910
rect 13078 5854 13200 5910
rect 12400 5786 13200 5854
rect 12400 5730 12526 5786
rect 12582 5730 12650 5786
rect 12706 5730 12774 5786
rect 12830 5730 12898 5786
rect 12954 5730 13022 5786
rect 13078 5730 13200 5786
rect 12400 5662 13200 5730
rect 12400 5606 12526 5662
rect 12582 5606 12650 5662
rect 12706 5606 12774 5662
rect 12830 5606 12898 5662
rect 12954 5606 13022 5662
rect 13078 5606 13200 5662
rect 12400 5538 13200 5606
rect 12400 5482 12526 5538
rect 12582 5482 12650 5538
rect 12706 5482 12774 5538
rect 12830 5482 12898 5538
rect 12954 5482 13022 5538
rect 13078 5482 13200 5538
rect 12400 5414 13200 5482
rect 12400 5358 12526 5414
rect 12582 5358 12650 5414
rect 12706 5358 12774 5414
rect 12830 5358 12898 5414
rect 12954 5358 13022 5414
rect 13078 5358 13200 5414
rect 12400 5290 13200 5358
rect 12400 5234 12526 5290
rect 12582 5234 12650 5290
rect 12706 5234 12774 5290
rect 12830 5234 12898 5290
rect 12954 5234 13022 5290
rect 13078 5234 13200 5290
rect 12400 5166 13200 5234
rect 12400 5110 12526 5166
rect 12582 5110 12650 5166
rect 12706 5110 12774 5166
rect 12830 5110 12898 5166
rect 12954 5110 13022 5166
rect 13078 5110 13200 5166
rect 12400 5042 13200 5110
rect 12400 4986 12526 5042
rect 12582 4986 12650 5042
rect 12706 4986 12774 5042
rect 12830 4986 12898 5042
rect 12954 4986 13022 5042
rect 13078 4986 13200 5042
rect 12400 4918 13200 4986
rect 12400 4862 12526 4918
rect 12582 4862 12650 4918
rect 12706 4862 12774 4918
rect 12830 4862 12898 4918
rect 12954 4862 13022 4918
rect 13078 4862 13200 4918
rect 12400 4794 13200 4862
rect 12400 4738 12526 4794
rect 12582 4738 12650 4794
rect 12706 4738 12774 4794
rect 12830 4738 12898 4794
rect 12954 4738 13022 4794
rect 13078 4738 13200 4794
rect 12400 4670 13200 4738
rect 12400 4614 12526 4670
rect 12582 4614 12650 4670
rect 12706 4614 12774 4670
rect 12830 4614 12898 4670
rect 12954 4614 13022 4670
rect 13078 4614 13200 4670
rect 12400 4546 13200 4614
rect 12400 4490 12526 4546
rect 12582 4490 12650 4546
rect 12706 4490 12774 4546
rect 12830 4490 12898 4546
rect 12954 4490 13022 4546
rect 13078 4490 13200 4546
rect 12400 4422 13200 4490
rect 12400 4366 12526 4422
rect 12582 4366 12650 4422
rect 12706 4366 12774 4422
rect 12830 4366 12898 4422
rect 12954 4366 13022 4422
rect 13078 4366 13200 4422
rect 12400 4298 13200 4366
rect 12400 4242 12526 4298
rect 12582 4242 12650 4298
rect 12706 4242 12774 4298
rect 12830 4242 12898 4298
rect 12954 4242 13022 4298
rect 13078 4242 13200 4298
rect 12400 4174 13200 4242
rect 12400 4118 12526 4174
rect 12582 4118 12650 4174
rect 12706 4118 12774 4174
rect 12830 4118 12898 4174
rect 12954 4118 13022 4174
rect 13078 4118 13200 4174
rect 12400 4050 13200 4118
rect 12400 3994 12526 4050
rect 12582 3994 12650 4050
rect 12706 3994 12774 4050
rect 12830 3994 12898 4050
rect 12954 3994 13022 4050
rect 13078 3994 13200 4050
rect 12400 3926 13200 3994
rect 12400 3870 12526 3926
rect 12582 3870 12650 3926
rect 12706 3870 12774 3926
rect 12830 3870 12898 3926
rect 12954 3870 13022 3926
rect 13078 3870 13200 3926
rect 12400 3802 13200 3870
rect 12400 3746 12526 3802
rect 12582 3746 12650 3802
rect 12706 3746 12774 3802
rect 12830 3746 12898 3802
rect 12954 3746 13022 3802
rect 13078 3746 13200 3802
rect 12400 3678 13200 3746
rect 12400 3622 12526 3678
rect 12582 3622 12650 3678
rect 12706 3622 12774 3678
rect 12830 3622 12898 3678
rect 12954 3622 13022 3678
rect 13078 3622 13200 3678
rect 12400 3554 13200 3622
rect 12400 3498 12526 3554
rect 12582 3498 12650 3554
rect 12706 3498 12774 3554
rect 12830 3498 12898 3554
rect 12954 3498 13022 3554
rect 13078 3498 13200 3554
rect 12400 3430 13200 3498
rect 12400 3374 12526 3430
rect 12582 3374 12650 3430
rect 12706 3374 12774 3430
rect 12830 3374 12898 3430
rect 12954 3374 13022 3430
rect 13078 3374 13200 3430
rect 12400 3306 13200 3374
rect 12400 3250 12526 3306
rect 12582 3250 12650 3306
rect 12706 3250 12774 3306
rect 12830 3250 12898 3306
rect 12954 3250 13022 3306
rect 13078 3250 13200 3306
rect 12400 3182 13200 3250
rect 12400 3126 12526 3182
rect 12582 3126 12650 3182
rect 12706 3126 12774 3182
rect 12830 3126 12898 3182
rect 12954 3126 13022 3182
rect 13078 3126 13200 3182
rect 12400 3058 13200 3126
rect 12400 3002 12526 3058
rect 12582 3002 12650 3058
rect 12706 3002 12774 3058
rect 12830 3002 12898 3058
rect 12954 3002 13022 3058
rect 13078 3002 13200 3058
rect 12400 2934 13200 3002
rect 12400 2878 12526 2934
rect 12582 2878 12650 2934
rect 12706 2878 12774 2934
rect 12830 2878 12898 2934
rect 12954 2878 13022 2934
rect 13078 2878 13200 2934
rect 12400 2810 13200 2878
rect 12400 2754 12526 2810
rect 12582 2754 12650 2810
rect 12706 2754 12774 2810
rect 12830 2754 12898 2810
rect 12954 2754 13022 2810
rect 13078 2754 13200 2810
rect 12400 2686 13200 2754
rect 12400 2630 12526 2686
rect 12582 2630 12650 2686
rect 12706 2630 12774 2686
rect 12830 2630 12898 2686
rect 12954 2630 13022 2686
rect 13078 2630 13200 2686
rect 12400 2562 13200 2630
rect 12400 2506 12526 2562
rect 12582 2506 12650 2562
rect 12706 2506 12774 2562
rect 12830 2506 12898 2562
rect 12954 2506 13022 2562
rect 13078 2506 13200 2562
rect 12400 2438 13200 2506
rect 12400 2382 12526 2438
rect 12582 2382 12650 2438
rect 12706 2382 12774 2438
rect 12830 2382 12898 2438
rect 12954 2382 13022 2438
rect 13078 2382 13200 2438
rect 12400 2314 13200 2382
rect 12400 2258 12526 2314
rect 12582 2258 12650 2314
rect 12706 2258 12774 2314
rect 12830 2258 12898 2314
rect 12954 2258 13022 2314
rect 13078 2258 13200 2314
rect 12400 2190 13200 2258
rect 12400 2134 12526 2190
rect 12582 2134 12650 2190
rect 12706 2134 12774 2190
rect 12830 2134 12898 2190
rect 12954 2134 13022 2190
rect 13078 2134 13200 2190
rect 12400 2066 13200 2134
rect 12400 2010 12526 2066
rect 12582 2010 12650 2066
rect 12706 2010 12774 2066
rect 12830 2010 12898 2066
rect 12954 2010 13022 2066
rect 13078 2010 13200 2066
rect 12400 1942 13200 2010
rect 12400 1886 12526 1942
rect 12582 1886 12650 1942
rect 12706 1886 12774 1942
rect 12830 1886 12898 1942
rect 12954 1886 13022 1942
rect 13078 1886 13200 1942
rect 12400 1818 13200 1886
rect 12400 1762 12526 1818
rect 12582 1762 12650 1818
rect 12706 1762 12774 1818
rect 12830 1762 12898 1818
rect 12954 1762 13022 1818
rect 13078 1762 13200 1818
rect 12400 1694 13200 1762
rect 12400 1638 12526 1694
rect 12582 1638 12650 1694
rect 12706 1638 12774 1694
rect 12830 1638 12898 1694
rect 12954 1638 13022 1694
rect 13078 1638 13200 1694
rect 12400 1570 13200 1638
rect 12400 1514 12526 1570
rect 12582 1514 12650 1570
rect 12706 1514 12774 1570
rect 12830 1514 12898 1570
rect 12954 1514 13022 1570
rect 13078 1514 13200 1570
rect 12400 1446 13200 1514
rect 12400 1390 12526 1446
rect 12582 1390 12650 1446
rect 12706 1390 12774 1446
rect 12830 1390 12898 1446
rect 12954 1390 13022 1446
rect 13078 1390 13200 1446
rect 12400 1322 13200 1390
rect 12400 1266 12526 1322
rect 12582 1266 12650 1322
rect 12706 1266 12774 1322
rect 12830 1266 12898 1322
rect 12954 1266 13022 1322
rect 13078 1266 13200 1322
rect 12400 1198 13200 1266
rect 12400 1142 12526 1198
rect 12582 1142 12650 1198
rect 12706 1142 12774 1198
rect 12830 1142 12898 1198
rect 12954 1142 13022 1198
rect 13078 1142 13200 1198
rect 12400 1074 13200 1142
rect 12400 1018 12526 1074
rect 12582 1018 12650 1074
rect 12706 1018 12774 1074
rect 12830 1018 12898 1074
rect 12954 1018 13022 1074
rect 13078 1018 13200 1074
rect 12400 950 13200 1018
rect 12400 894 12526 950
rect 12582 894 12650 950
rect 12706 894 12774 950
rect 12830 894 12898 950
rect 12954 894 13022 950
rect 13078 894 13200 950
rect 12400 826 13200 894
rect 12400 770 12526 826
rect 12582 770 12650 826
rect 12706 770 12774 826
rect 12830 770 12898 826
rect 12954 770 13022 826
rect 13078 770 13200 826
rect 12400 702 13200 770
rect 12400 646 12526 702
rect 12582 646 12650 702
rect 12706 646 12774 702
rect 12830 646 12898 702
rect 12954 646 13022 702
rect 13078 646 13200 702
rect 12400 578 13200 646
rect 12400 522 12526 578
rect 12582 522 12650 578
rect 12706 522 12774 578
rect 12830 522 12898 578
rect 12954 522 13022 578
rect 13078 522 13200 578
rect 12400 454 13200 522
rect 12400 400 12526 454
rect 266 398 12526 400
rect 12582 398 12650 454
rect 12706 398 12774 454
rect 12830 398 12898 454
rect 12954 398 13022 454
rect 13078 398 13200 454
rect -400 330 13200 398
rect -400 274 -286 330
rect -230 274 -162 330
rect -106 274 -38 330
rect 18 274 86 330
rect 142 274 210 330
rect 266 302 12526 330
rect 266 274 415 302
rect -400 246 415 274
rect 471 246 557 302
rect 613 246 699 302
rect 755 246 841 302
rect 897 246 983 302
rect 1039 246 1125 302
rect 1181 246 1267 302
rect 1323 246 1409 302
rect 1465 246 1551 302
rect 1607 246 1693 302
rect 1749 246 1835 302
rect 1891 246 1977 302
rect 2033 246 2119 302
rect 2175 246 2261 302
rect 2317 246 2403 302
rect 2459 246 2545 302
rect 2601 246 2687 302
rect 2743 246 2829 302
rect 2885 246 2971 302
rect 3027 246 3113 302
rect 3169 246 3255 302
rect 3311 246 3397 302
rect 3453 246 3539 302
rect 3595 246 3681 302
rect 3737 246 3823 302
rect 3879 246 3965 302
rect 4021 246 4107 302
rect 4163 246 4249 302
rect 4305 246 4391 302
rect 4447 246 4533 302
rect 4589 246 4675 302
rect 4731 246 4817 302
rect 4873 246 4959 302
rect 5015 246 5101 302
rect 5157 246 5243 302
rect 5299 246 5385 302
rect 5441 246 5527 302
rect 5583 246 5669 302
rect 5725 246 5811 302
rect 5867 246 5953 302
rect 6009 246 6095 302
rect 6151 246 6237 302
rect 6293 246 6379 302
rect 6435 246 6521 302
rect 6577 246 6663 302
rect 6719 246 6805 302
rect 6861 246 6947 302
rect 7003 246 7089 302
rect 7145 246 7231 302
rect 7287 246 7373 302
rect 7429 246 7515 302
rect 7571 246 7657 302
rect 7713 246 7799 302
rect 7855 246 7941 302
rect 7997 246 8083 302
rect 8139 246 8225 302
rect 8281 246 8367 302
rect 8423 246 8509 302
rect 8565 246 8651 302
rect 8707 246 8793 302
rect 8849 246 8935 302
rect 8991 246 9077 302
rect 9133 246 9219 302
rect 9275 246 9361 302
rect 9417 246 9503 302
rect 9559 246 9645 302
rect 9701 246 9787 302
rect 9843 246 9929 302
rect 9985 246 10071 302
rect 10127 246 10213 302
rect 10269 246 10355 302
rect 10411 246 10497 302
rect 10553 246 10639 302
rect 10695 246 10781 302
rect 10837 246 10923 302
rect 10979 246 11065 302
rect 11121 246 11207 302
rect 11263 246 11349 302
rect 11405 246 11491 302
rect 11547 246 11633 302
rect 11689 246 11775 302
rect 11831 246 11917 302
rect 11973 246 12059 302
rect 12115 246 12201 302
rect 12257 246 12343 302
rect 12399 274 12526 302
rect 12582 274 12650 330
rect 12706 274 12774 330
rect 12830 274 12898 330
rect 12954 274 13022 330
rect 13078 274 13200 330
rect 12399 246 13200 274
rect -400 206 13200 246
rect -400 150 -286 206
rect -230 150 -162 206
rect -106 150 -38 206
rect 18 150 86 206
rect 142 150 210 206
rect 266 160 12526 206
rect 266 150 415 160
rect -400 104 415 150
rect 471 104 557 160
rect 613 104 699 160
rect 755 104 841 160
rect 897 104 983 160
rect 1039 104 1125 160
rect 1181 104 1267 160
rect 1323 104 1409 160
rect 1465 104 1551 160
rect 1607 104 1693 160
rect 1749 104 1835 160
rect 1891 104 1977 160
rect 2033 104 2119 160
rect 2175 104 2261 160
rect 2317 104 2403 160
rect 2459 104 2545 160
rect 2601 104 2687 160
rect 2743 104 2829 160
rect 2885 104 2971 160
rect 3027 104 3113 160
rect 3169 104 3255 160
rect 3311 104 3397 160
rect 3453 104 3539 160
rect 3595 104 3681 160
rect 3737 104 3823 160
rect 3879 104 3965 160
rect 4021 104 4107 160
rect 4163 104 4249 160
rect 4305 104 4391 160
rect 4447 104 4533 160
rect 4589 104 4675 160
rect 4731 104 4817 160
rect 4873 104 4959 160
rect 5015 104 5101 160
rect 5157 104 5243 160
rect 5299 104 5385 160
rect 5441 104 5527 160
rect 5583 104 5669 160
rect 5725 104 5811 160
rect 5867 104 5953 160
rect 6009 104 6095 160
rect 6151 104 6237 160
rect 6293 104 6379 160
rect 6435 104 6521 160
rect 6577 104 6663 160
rect 6719 104 6805 160
rect 6861 104 6947 160
rect 7003 104 7089 160
rect 7145 104 7231 160
rect 7287 104 7373 160
rect 7429 104 7515 160
rect 7571 104 7657 160
rect 7713 104 7799 160
rect 7855 104 7941 160
rect 7997 104 8083 160
rect 8139 104 8225 160
rect 8281 104 8367 160
rect 8423 104 8509 160
rect 8565 104 8651 160
rect 8707 104 8793 160
rect 8849 104 8935 160
rect 8991 104 9077 160
rect 9133 104 9219 160
rect 9275 104 9361 160
rect 9417 104 9503 160
rect 9559 104 9645 160
rect 9701 104 9787 160
rect 9843 104 9929 160
rect 9985 104 10071 160
rect 10127 104 10213 160
rect 10269 104 10355 160
rect 10411 104 10497 160
rect 10553 104 10639 160
rect 10695 104 10781 160
rect 10837 104 10923 160
rect 10979 104 11065 160
rect 11121 104 11207 160
rect 11263 104 11349 160
rect 11405 104 11491 160
rect 11547 104 11633 160
rect 11689 104 11775 160
rect 11831 104 11917 160
rect 11973 104 12059 160
rect 12115 104 12201 160
rect 12257 104 12343 160
rect 12399 150 12526 160
rect 12582 150 12650 206
rect 12706 150 12774 206
rect 12830 150 12898 206
rect 12954 150 13022 206
rect 13078 150 13200 206
rect 12399 104 13200 150
rect -400 0 13200 104
<< via2 >>
rect -254 12893 -198 12949
rect -130 12893 -74 12949
rect -6 12893 50 12949
rect 118 12893 174 12949
rect 242 12893 298 12949
rect 366 12893 422 12949
rect 490 12893 546 12949
rect 614 12893 670 12949
rect 738 12893 794 12949
rect 862 12893 918 12949
rect 986 12893 1042 12949
rect 1110 12893 1166 12949
rect 1234 12893 1290 12949
rect 1358 12893 1414 12949
rect 1482 12893 1538 12949
rect 1606 12893 1662 12949
rect 1730 12893 1786 12949
rect 1854 12893 1910 12949
rect 1978 12893 2034 12949
rect 2102 12893 2158 12949
rect 2226 12893 2282 12949
rect 2350 12893 2406 12949
rect 2474 12893 2530 12949
rect 2598 12893 2654 12949
rect 2722 12893 2778 12949
rect 2846 12893 2902 12949
rect 2970 12893 3026 12949
rect 3094 12893 3150 12949
rect 3218 12893 3274 12949
rect 3342 12893 3398 12949
rect 3466 12893 3522 12949
rect 3590 12893 3646 12949
rect 3714 12893 3770 12949
rect 3838 12893 3894 12949
rect 3962 12893 4018 12949
rect 4086 12893 4142 12949
rect 4210 12893 4266 12949
rect 4334 12893 4390 12949
rect 4458 12893 4514 12949
rect 4582 12893 4638 12949
rect 4706 12893 4762 12949
rect 4830 12893 4886 12949
rect 4954 12893 5010 12949
rect 5078 12893 5134 12949
rect 5202 12893 5258 12949
rect 5326 12893 5382 12949
rect 5450 12893 5506 12949
rect 5574 12893 5630 12949
rect 5698 12893 5754 12949
rect 5822 12893 5878 12949
rect 5946 12893 6002 12949
rect 6070 12893 6126 12949
rect 6194 12893 6250 12949
rect 6318 12893 6374 12949
rect 6442 12893 6498 12949
rect 6566 12893 6622 12949
rect 6690 12893 6746 12949
rect 6814 12893 6870 12949
rect 6938 12893 6994 12949
rect 7062 12893 7118 12949
rect 7186 12893 7242 12949
rect 7310 12893 7366 12949
rect 7434 12893 7490 12949
rect 7558 12893 7614 12949
rect 7682 12893 7738 12949
rect 7806 12893 7862 12949
rect 7930 12893 7986 12949
rect 8054 12893 8110 12949
rect 8178 12893 8234 12949
rect 8302 12893 8358 12949
rect 8426 12893 8482 12949
rect 8550 12893 8606 12949
rect 8674 12893 8730 12949
rect 8798 12893 8854 12949
rect 8922 12893 8978 12949
rect 9046 12893 9102 12949
rect 9170 12893 9226 12949
rect 9294 12893 9350 12949
rect 9418 12893 9474 12949
rect 9542 12893 9598 12949
rect 9666 12893 9722 12949
rect 9790 12893 9846 12949
rect 9914 12893 9970 12949
rect 10038 12893 10094 12949
rect 10162 12893 10218 12949
rect 10286 12893 10342 12949
rect 10410 12893 10466 12949
rect 10534 12893 10590 12949
rect 10658 12893 10714 12949
rect 10782 12893 10838 12949
rect 10906 12893 10962 12949
rect 11030 12893 11086 12949
rect 11154 12893 11210 12949
rect 11278 12893 11334 12949
rect 11402 12893 11458 12949
rect 11526 12893 11582 12949
rect 11650 12893 11706 12949
rect 11774 12893 11830 12949
rect 11898 12893 11954 12949
rect 12022 12893 12078 12949
rect 12146 12893 12202 12949
rect 12270 12893 12326 12949
rect 12394 12893 12450 12949
rect 12518 12893 12574 12949
rect 12642 12893 12698 12949
rect 12766 12893 12822 12949
rect 12890 12893 12946 12949
rect 13014 12893 13070 12949
rect -254 12769 -198 12825
rect -130 12769 -74 12825
rect -6 12769 50 12825
rect 118 12769 174 12825
rect 242 12769 298 12825
rect 366 12769 422 12825
rect 490 12769 546 12825
rect 614 12769 670 12825
rect 738 12769 794 12825
rect 862 12769 918 12825
rect 986 12769 1042 12825
rect 1110 12769 1166 12825
rect 1234 12769 1290 12825
rect 1358 12769 1414 12825
rect 1482 12769 1538 12825
rect 1606 12769 1662 12825
rect 1730 12769 1786 12825
rect 1854 12769 1910 12825
rect 1978 12769 2034 12825
rect 2102 12769 2158 12825
rect 2226 12769 2282 12825
rect 2350 12769 2406 12825
rect 2474 12769 2530 12825
rect 2598 12769 2654 12825
rect 2722 12769 2778 12825
rect 2846 12769 2902 12825
rect 2970 12769 3026 12825
rect 3094 12769 3150 12825
rect 3218 12769 3274 12825
rect 3342 12769 3398 12825
rect 3466 12769 3522 12825
rect 3590 12769 3646 12825
rect 3714 12769 3770 12825
rect 3838 12769 3894 12825
rect 3962 12769 4018 12825
rect 4086 12769 4142 12825
rect 4210 12769 4266 12825
rect 4334 12769 4390 12825
rect 4458 12769 4514 12825
rect 4582 12769 4638 12825
rect 4706 12769 4762 12825
rect 4830 12769 4886 12825
rect 4954 12769 5010 12825
rect 5078 12769 5134 12825
rect 5202 12769 5258 12825
rect 5326 12769 5382 12825
rect 5450 12769 5506 12825
rect 5574 12769 5630 12825
rect 5698 12769 5754 12825
rect 5822 12769 5878 12825
rect 5946 12769 6002 12825
rect 6070 12769 6126 12825
rect 6194 12769 6250 12825
rect 6318 12769 6374 12825
rect 6442 12769 6498 12825
rect 6566 12769 6622 12825
rect 6690 12769 6746 12825
rect 6814 12769 6870 12825
rect 6938 12769 6994 12825
rect 7062 12769 7118 12825
rect 7186 12769 7242 12825
rect 7310 12769 7366 12825
rect 7434 12769 7490 12825
rect 7558 12769 7614 12825
rect 7682 12769 7738 12825
rect 7806 12769 7862 12825
rect 7930 12769 7986 12825
rect 8054 12769 8110 12825
rect 8178 12769 8234 12825
rect 8302 12769 8358 12825
rect 8426 12769 8482 12825
rect 8550 12769 8606 12825
rect 8674 12769 8730 12825
rect 8798 12769 8854 12825
rect 8922 12769 8978 12825
rect 9046 12769 9102 12825
rect 9170 12769 9226 12825
rect 9294 12769 9350 12825
rect 9418 12769 9474 12825
rect 9542 12769 9598 12825
rect 9666 12769 9722 12825
rect 9790 12769 9846 12825
rect 9914 12769 9970 12825
rect 10038 12769 10094 12825
rect 10162 12769 10218 12825
rect 10286 12769 10342 12825
rect 10410 12769 10466 12825
rect 10534 12769 10590 12825
rect 10658 12769 10714 12825
rect 10782 12769 10838 12825
rect 10906 12769 10962 12825
rect 11030 12769 11086 12825
rect 11154 12769 11210 12825
rect 11278 12769 11334 12825
rect 11402 12769 11458 12825
rect 11526 12769 11582 12825
rect 11650 12769 11706 12825
rect 11774 12769 11830 12825
rect 11898 12769 11954 12825
rect 12022 12769 12078 12825
rect 12146 12769 12202 12825
rect 12270 12769 12326 12825
rect 12394 12769 12450 12825
rect 12518 12769 12574 12825
rect 12642 12769 12698 12825
rect 12766 12769 12822 12825
rect 12890 12769 12946 12825
rect 13014 12769 13070 12825
rect -254 12645 -198 12701
rect -130 12645 -74 12701
rect -6 12645 50 12701
rect 118 12645 174 12701
rect 242 12645 298 12701
rect 366 12645 422 12701
rect 490 12645 546 12701
rect 614 12645 670 12701
rect 738 12645 794 12701
rect 862 12645 918 12701
rect 986 12645 1042 12701
rect 1110 12645 1166 12701
rect 1234 12645 1290 12701
rect 1358 12645 1414 12701
rect 1482 12645 1538 12701
rect 1606 12645 1662 12701
rect 1730 12645 1786 12701
rect 1854 12645 1910 12701
rect 1978 12645 2034 12701
rect 2102 12645 2158 12701
rect 2226 12645 2282 12701
rect 2350 12645 2406 12701
rect 2474 12645 2530 12701
rect 2598 12645 2654 12701
rect 2722 12645 2778 12701
rect 2846 12645 2902 12701
rect 2970 12645 3026 12701
rect 3094 12645 3150 12701
rect 3218 12645 3274 12701
rect 3342 12645 3398 12701
rect 3466 12645 3522 12701
rect 3590 12645 3646 12701
rect 3714 12645 3770 12701
rect 3838 12645 3894 12701
rect 3962 12645 4018 12701
rect 4086 12645 4142 12701
rect 4210 12645 4266 12701
rect 4334 12645 4390 12701
rect 4458 12645 4514 12701
rect 4582 12645 4638 12701
rect 4706 12645 4762 12701
rect 4830 12645 4886 12701
rect 4954 12645 5010 12701
rect 5078 12645 5134 12701
rect 5202 12645 5258 12701
rect 5326 12645 5382 12701
rect 5450 12645 5506 12701
rect 5574 12645 5630 12701
rect 5698 12645 5754 12701
rect 5822 12645 5878 12701
rect 5946 12645 6002 12701
rect 6070 12645 6126 12701
rect 6194 12645 6250 12701
rect 6318 12645 6374 12701
rect 6442 12645 6498 12701
rect 6566 12645 6622 12701
rect 6690 12645 6746 12701
rect 6814 12645 6870 12701
rect 6938 12645 6994 12701
rect 7062 12645 7118 12701
rect 7186 12645 7242 12701
rect 7310 12645 7366 12701
rect 7434 12645 7490 12701
rect 7558 12645 7614 12701
rect 7682 12645 7738 12701
rect 7806 12645 7862 12701
rect 7930 12645 7986 12701
rect 8054 12645 8110 12701
rect 8178 12645 8234 12701
rect 8302 12645 8358 12701
rect 8426 12645 8482 12701
rect 8550 12645 8606 12701
rect 8674 12645 8730 12701
rect 8798 12645 8854 12701
rect 8922 12645 8978 12701
rect 9046 12645 9102 12701
rect 9170 12645 9226 12701
rect 9294 12645 9350 12701
rect 9418 12645 9474 12701
rect 9542 12645 9598 12701
rect 9666 12645 9722 12701
rect 9790 12645 9846 12701
rect 9914 12645 9970 12701
rect 10038 12645 10094 12701
rect 10162 12645 10218 12701
rect 10286 12645 10342 12701
rect 10410 12645 10466 12701
rect 10534 12645 10590 12701
rect 10658 12645 10714 12701
rect 10782 12645 10838 12701
rect 10906 12645 10962 12701
rect 11030 12645 11086 12701
rect 11154 12645 11210 12701
rect 11278 12645 11334 12701
rect 11402 12645 11458 12701
rect 11526 12645 11582 12701
rect 11650 12645 11706 12701
rect 11774 12645 11830 12701
rect 11898 12645 11954 12701
rect 12022 12645 12078 12701
rect 12146 12645 12202 12701
rect 12270 12645 12326 12701
rect 12394 12645 12450 12701
rect 12518 12645 12574 12701
rect 12642 12645 12698 12701
rect 12766 12645 12822 12701
rect 12890 12645 12946 12701
rect 13014 12645 13070 12701
rect -254 12521 -198 12577
rect -130 12521 -74 12577
rect -6 12521 50 12577
rect 118 12521 174 12577
rect 242 12521 298 12577
rect 366 12521 422 12577
rect 490 12521 546 12577
rect 614 12521 670 12577
rect 738 12521 794 12577
rect 862 12521 918 12577
rect 986 12521 1042 12577
rect 1110 12521 1166 12577
rect 1234 12521 1290 12577
rect 1358 12521 1414 12577
rect 1482 12521 1538 12577
rect 1606 12521 1662 12577
rect 1730 12521 1786 12577
rect 1854 12521 1910 12577
rect 1978 12521 2034 12577
rect 2102 12521 2158 12577
rect 2226 12521 2282 12577
rect 2350 12521 2406 12577
rect 2474 12521 2530 12577
rect 2598 12521 2654 12577
rect 2722 12521 2778 12577
rect 2846 12521 2902 12577
rect 2970 12521 3026 12577
rect 3094 12521 3150 12577
rect 3218 12521 3274 12577
rect 3342 12521 3398 12577
rect 3466 12521 3522 12577
rect 3590 12521 3646 12577
rect 3714 12521 3770 12577
rect 3838 12521 3894 12577
rect 3962 12521 4018 12577
rect 4086 12521 4142 12577
rect 4210 12521 4266 12577
rect 4334 12521 4390 12577
rect 4458 12521 4514 12577
rect 4582 12521 4638 12577
rect 4706 12521 4762 12577
rect 4830 12521 4886 12577
rect 4954 12521 5010 12577
rect 5078 12521 5134 12577
rect 5202 12521 5258 12577
rect 5326 12521 5382 12577
rect 5450 12521 5506 12577
rect 5574 12521 5630 12577
rect 5698 12521 5754 12577
rect 5822 12521 5878 12577
rect 5946 12521 6002 12577
rect 6070 12521 6126 12577
rect 6194 12521 6250 12577
rect 6318 12521 6374 12577
rect 6442 12521 6498 12577
rect 6566 12521 6622 12577
rect 6690 12521 6746 12577
rect 6814 12521 6870 12577
rect 6938 12521 6994 12577
rect 7062 12521 7118 12577
rect 7186 12521 7242 12577
rect 7310 12521 7366 12577
rect 7434 12521 7490 12577
rect 7558 12521 7614 12577
rect 7682 12521 7738 12577
rect 7806 12521 7862 12577
rect 7930 12521 7986 12577
rect 8054 12521 8110 12577
rect 8178 12521 8234 12577
rect 8302 12521 8358 12577
rect 8426 12521 8482 12577
rect 8550 12521 8606 12577
rect 8674 12521 8730 12577
rect 8798 12521 8854 12577
rect 8922 12521 8978 12577
rect 9046 12521 9102 12577
rect 9170 12521 9226 12577
rect 9294 12521 9350 12577
rect 9418 12521 9474 12577
rect 9542 12521 9598 12577
rect 9666 12521 9722 12577
rect 9790 12521 9846 12577
rect 9914 12521 9970 12577
rect 10038 12521 10094 12577
rect 10162 12521 10218 12577
rect 10286 12521 10342 12577
rect 10410 12521 10466 12577
rect 10534 12521 10590 12577
rect 10658 12521 10714 12577
rect 10782 12521 10838 12577
rect 10906 12521 10962 12577
rect 11030 12521 11086 12577
rect 11154 12521 11210 12577
rect 11278 12521 11334 12577
rect 11402 12521 11458 12577
rect 11526 12521 11582 12577
rect 11650 12521 11706 12577
rect 11774 12521 11830 12577
rect 11898 12521 11954 12577
rect 12022 12521 12078 12577
rect 12146 12521 12202 12577
rect 12270 12521 12326 12577
rect 12394 12521 12450 12577
rect 12518 12521 12574 12577
rect 12642 12521 12698 12577
rect 12766 12521 12822 12577
rect 12890 12521 12946 12577
rect 13014 12521 13070 12577
rect -286 12302 -230 12358
rect -162 12302 -106 12358
rect -38 12302 18 12358
rect 86 12302 142 12358
rect 210 12302 266 12358
rect -286 12178 -230 12234
rect -162 12178 -106 12234
rect -38 12178 18 12234
rect 86 12178 142 12234
rect 210 12178 266 12234
rect -286 12054 -230 12110
rect -162 12054 -106 12110
rect -38 12054 18 12110
rect 86 12054 142 12110
rect 210 12054 266 12110
rect -286 11930 -230 11986
rect -162 11930 -106 11986
rect -38 11930 18 11986
rect 86 11930 142 11986
rect 210 11930 266 11986
rect -286 11806 -230 11862
rect -162 11806 -106 11862
rect -38 11806 18 11862
rect 86 11806 142 11862
rect 210 11806 266 11862
rect -286 11682 -230 11738
rect -162 11682 -106 11738
rect -38 11682 18 11738
rect 86 11682 142 11738
rect 210 11682 266 11738
rect -286 11558 -230 11614
rect -162 11558 -106 11614
rect -38 11558 18 11614
rect 86 11558 142 11614
rect 210 11558 266 11614
rect -286 11434 -230 11490
rect -162 11434 -106 11490
rect -38 11434 18 11490
rect 86 11434 142 11490
rect 210 11434 266 11490
rect -286 11310 -230 11366
rect -162 11310 -106 11366
rect -38 11310 18 11366
rect 86 11310 142 11366
rect 210 11310 266 11366
rect -286 11186 -230 11242
rect -162 11186 -106 11242
rect -38 11186 18 11242
rect 86 11186 142 11242
rect 210 11186 266 11242
rect -286 11062 -230 11118
rect -162 11062 -106 11118
rect -38 11062 18 11118
rect 86 11062 142 11118
rect 210 11062 266 11118
rect -286 10938 -230 10994
rect -162 10938 -106 10994
rect -38 10938 18 10994
rect 86 10938 142 10994
rect 210 10938 266 10994
rect -286 10814 -230 10870
rect -162 10814 -106 10870
rect -38 10814 18 10870
rect 86 10814 142 10870
rect 210 10814 266 10870
rect -286 10690 -230 10746
rect -162 10690 -106 10746
rect -38 10690 18 10746
rect 86 10690 142 10746
rect 210 10690 266 10746
rect -286 10566 -230 10622
rect -162 10566 -106 10622
rect -38 10566 18 10622
rect 86 10566 142 10622
rect 210 10566 266 10622
rect -286 10442 -230 10498
rect -162 10442 -106 10498
rect -38 10442 18 10498
rect 86 10442 142 10498
rect 210 10442 266 10498
rect -286 10318 -230 10374
rect -162 10318 -106 10374
rect -38 10318 18 10374
rect 86 10318 142 10374
rect 210 10318 266 10374
rect -286 10194 -230 10250
rect -162 10194 -106 10250
rect -38 10194 18 10250
rect 86 10194 142 10250
rect 210 10194 266 10250
rect -286 10070 -230 10126
rect -162 10070 -106 10126
rect -38 10070 18 10126
rect 86 10070 142 10126
rect 210 10070 266 10126
rect -286 9946 -230 10002
rect -162 9946 -106 10002
rect -38 9946 18 10002
rect 86 9946 142 10002
rect 210 9946 266 10002
rect -286 9822 -230 9878
rect -162 9822 -106 9878
rect -38 9822 18 9878
rect 86 9822 142 9878
rect 210 9822 266 9878
rect -286 9698 -230 9754
rect -162 9698 -106 9754
rect -38 9698 18 9754
rect 86 9698 142 9754
rect 210 9698 266 9754
rect -286 9574 -230 9630
rect -162 9574 -106 9630
rect -38 9574 18 9630
rect 86 9574 142 9630
rect 210 9574 266 9630
rect -286 9450 -230 9506
rect -162 9450 -106 9506
rect -38 9450 18 9506
rect 86 9450 142 9506
rect 210 9450 266 9506
rect -286 9326 -230 9382
rect -162 9326 -106 9382
rect -38 9326 18 9382
rect 86 9326 142 9382
rect 210 9326 266 9382
rect -286 9202 -230 9258
rect -162 9202 -106 9258
rect -38 9202 18 9258
rect 86 9202 142 9258
rect 210 9202 266 9258
rect -286 9078 -230 9134
rect -162 9078 -106 9134
rect -38 9078 18 9134
rect 86 9078 142 9134
rect 210 9078 266 9134
rect -286 8954 -230 9010
rect -162 8954 -106 9010
rect -38 8954 18 9010
rect 86 8954 142 9010
rect 210 8954 266 9010
rect -286 8830 -230 8886
rect -162 8830 -106 8886
rect -38 8830 18 8886
rect 86 8830 142 8886
rect 210 8830 266 8886
rect -286 8706 -230 8762
rect -162 8706 -106 8762
rect -38 8706 18 8762
rect 86 8706 142 8762
rect 210 8706 266 8762
rect -286 8582 -230 8638
rect -162 8582 -106 8638
rect -38 8582 18 8638
rect 86 8582 142 8638
rect 210 8582 266 8638
rect -286 8458 -230 8514
rect -162 8458 -106 8514
rect -38 8458 18 8514
rect 86 8458 142 8514
rect 210 8458 266 8514
rect -286 8334 -230 8390
rect -162 8334 -106 8390
rect -38 8334 18 8390
rect 86 8334 142 8390
rect 210 8334 266 8390
rect -286 8210 -230 8266
rect -162 8210 -106 8266
rect -38 8210 18 8266
rect 86 8210 142 8266
rect 210 8210 266 8266
rect -286 8086 -230 8142
rect -162 8086 -106 8142
rect -38 8086 18 8142
rect 86 8086 142 8142
rect 210 8086 266 8142
rect -286 7962 -230 8018
rect -162 7962 -106 8018
rect -38 7962 18 8018
rect 86 7962 142 8018
rect 210 7962 266 8018
rect -286 7838 -230 7894
rect -162 7838 -106 7894
rect -38 7838 18 7894
rect 86 7838 142 7894
rect 210 7838 266 7894
rect -286 7714 -230 7770
rect -162 7714 -106 7770
rect -38 7714 18 7770
rect 86 7714 142 7770
rect 210 7714 266 7770
rect -286 7590 -230 7646
rect -162 7590 -106 7646
rect -38 7590 18 7646
rect 86 7590 142 7646
rect 210 7590 266 7646
rect -286 7466 -230 7522
rect -162 7466 -106 7522
rect -38 7466 18 7522
rect 86 7466 142 7522
rect 210 7466 266 7522
rect -286 7342 -230 7398
rect -162 7342 -106 7398
rect -38 7342 18 7398
rect 86 7342 142 7398
rect 210 7342 266 7398
rect -286 7218 -230 7274
rect -162 7218 -106 7274
rect -38 7218 18 7274
rect 86 7218 142 7274
rect 210 7218 266 7274
rect -286 7094 -230 7150
rect -162 7094 -106 7150
rect -38 7094 18 7150
rect 86 7094 142 7150
rect 210 7094 266 7150
rect -286 6970 -230 7026
rect -162 6970 -106 7026
rect -38 6970 18 7026
rect 86 6970 142 7026
rect 210 6970 266 7026
rect -286 6846 -230 6902
rect -162 6846 -106 6902
rect -38 6846 18 6902
rect 86 6846 142 6902
rect 210 6846 266 6902
rect -286 6722 -230 6778
rect -162 6722 -106 6778
rect -38 6722 18 6778
rect 86 6722 142 6778
rect 210 6722 266 6778
rect -286 6598 -230 6654
rect -162 6598 -106 6654
rect -38 6598 18 6654
rect 86 6598 142 6654
rect 210 6598 266 6654
rect -286 6474 -230 6530
rect -162 6474 -106 6530
rect -38 6474 18 6530
rect 86 6474 142 6530
rect 210 6474 266 6530
rect -286 6350 -230 6406
rect -162 6350 -106 6406
rect -38 6350 18 6406
rect 86 6350 142 6406
rect 210 6350 266 6406
rect -286 6226 -230 6282
rect -162 6226 -106 6282
rect -38 6226 18 6282
rect 86 6226 142 6282
rect 210 6226 266 6282
rect -286 6102 -230 6158
rect -162 6102 -106 6158
rect -38 6102 18 6158
rect 86 6102 142 6158
rect 210 6102 266 6158
rect -286 5978 -230 6034
rect -162 5978 -106 6034
rect -38 5978 18 6034
rect 86 5978 142 6034
rect 210 5978 266 6034
rect -286 5854 -230 5910
rect -162 5854 -106 5910
rect -38 5854 18 5910
rect 86 5854 142 5910
rect 210 5854 266 5910
rect -286 5730 -230 5786
rect -162 5730 -106 5786
rect -38 5730 18 5786
rect 86 5730 142 5786
rect 210 5730 266 5786
rect -286 5606 -230 5662
rect -162 5606 -106 5662
rect -38 5606 18 5662
rect 86 5606 142 5662
rect 210 5606 266 5662
rect -286 5482 -230 5538
rect -162 5482 -106 5538
rect -38 5482 18 5538
rect 86 5482 142 5538
rect 210 5482 266 5538
rect -286 5358 -230 5414
rect -162 5358 -106 5414
rect -38 5358 18 5414
rect 86 5358 142 5414
rect 210 5358 266 5414
rect -286 5234 -230 5290
rect -162 5234 -106 5290
rect -38 5234 18 5290
rect 86 5234 142 5290
rect 210 5234 266 5290
rect -286 5110 -230 5166
rect -162 5110 -106 5166
rect -38 5110 18 5166
rect 86 5110 142 5166
rect 210 5110 266 5166
rect -286 4986 -230 5042
rect -162 4986 -106 5042
rect -38 4986 18 5042
rect 86 4986 142 5042
rect 210 4986 266 5042
rect -286 4862 -230 4918
rect -162 4862 -106 4918
rect -38 4862 18 4918
rect 86 4862 142 4918
rect 210 4862 266 4918
rect -286 4738 -230 4794
rect -162 4738 -106 4794
rect -38 4738 18 4794
rect 86 4738 142 4794
rect 210 4738 266 4794
rect -286 4614 -230 4670
rect -162 4614 -106 4670
rect -38 4614 18 4670
rect 86 4614 142 4670
rect 210 4614 266 4670
rect -286 4490 -230 4546
rect -162 4490 -106 4546
rect -38 4490 18 4546
rect 86 4490 142 4546
rect 210 4490 266 4546
rect -286 4366 -230 4422
rect -162 4366 -106 4422
rect -38 4366 18 4422
rect 86 4366 142 4422
rect 210 4366 266 4422
rect -286 4242 -230 4298
rect -162 4242 -106 4298
rect -38 4242 18 4298
rect 86 4242 142 4298
rect 210 4242 266 4298
rect -286 4118 -230 4174
rect -162 4118 -106 4174
rect -38 4118 18 4174
rect 86 4118 142 4174
rect 210 4118 266 4174
rect -286 3994 -230 4050
rect -162 3994 -106 4050
rect -38 3994 18 4050
rect 86 3994 142 4050
rect 210 3994 266 4050
rect -286 3870 -230 3926
rect -162 3870 -106 3926
rect -38 3870 18 3926
rect 86 3870 142 3926
rect 210 3870 266 3926
rect -286 3746 -230 3802
rect -162 3746 -106 3802
rect -38 3746 18 3802
rect 86 3746 142 3802
rect 210 3746 266 3802
rect -286 3622 -230 3678
rect -162 3622 -106 3678
rect -38 3622 18 3678
rect 86 3622 142 3678
rect 210 3622 266 3678
rect -286 3498 -230 3554
rect -162 3498 -106 3554
rect -38 3498 18 3554
rect 86 3498 142 3554
rect 210 3498 266 3554
rect -286 3374 -230 3430
rect -162 3374 -106 3430
rect -38 3374 18 3430
rect 86 3374 142 3430
rect 210 3374 266 3430
rect -286 3250 -230 3306
rect -162 3250 -106 3306
rect -38 3250 18 3306
rect 86 3250 142 3306
rect 210 3250 266 3306
rect -286 3126 -230 3182
rect -162 3126 -106 3182
rect -38 3126 18 3182
rect 86 3126 142 3182
rect 210 3126 266 3182
rect -286 3002 -230 3058
rect -162 3002 -106 3058
rect -38 3002 18 3058
rect 86 3002 142 3058
rect 210 3002 266 3058
rect -286 2878 -230 2934
rect -162 2878 -106 2934
rect -38 2878 18 2934
rect 86 2878 142 2934
rect 210 2878 266 2934
rect -286 2754 -230 2810
rect -162 2754 -106 2810
rect -38 2754 18 2810
rect 86 2754 142 2810
rect 210 2754 266 2810
rect -286 2630 -230 2686
rect -162 2630 -106 2686
rect -38 2630 18 2686
rect 86 2630 142 2686
rect 210 2630 266 2686
rect -286 2506 -230 2562
rect -162 2506 -106 2562
rect -38 2506 18 2562
rect 86 2506 142 2562
rect 210 2506 266 2562
rect -286 2382 -230 2438
rect -162 2382 -106 2438
rect -38 2382 18 2438
rect 86 2382 142 2438
rect 210 2382 266 2438
rect -286 2258 -230 2314
rect -162 2258 -106 2314
rect -38 2258 18 2314
rect 86 2258 142 2314
rect 210 2258 266 2314
rect -286 2134 -230 2190
rect -162 2134 -106 2190
rect -38 2134 18 2190
rect 86 2134 142 2190
rect 210 2134 266 2190
rect -286 2010 -230 2066
rect -162 2010 -106 2066
rect -38 2010 18 2066
rect 86 2010 142 2066
rect 210 2010 266 2066
rect -286 1886 -230 1942
rect -162 1886 -106 1942
rect -38 1886 18 1942
rect 86 1886 142 1942
rect 210 1886 266 1942
rect -286 1762 -230 1818
rect -162 1762 -106 1818
rect -38 1762 18 1818
rect 86 1762 142 1818
rect 210 1762 266 1818
rect -286 1638 -230 1694
rect -162 1638 -106 1694
rect -38 1638 18 1694
rect 86 1638 142 1694
rect 210 1638 266 1694
rect -286 1514 -230 1570
rect -162 1514 -106 1570
rect -38 1514 18 1570
rect 86 1514 142 1570
rect 210 1514 266 1570
rect -286 1390 -230 1446
rect -162 1390 -106 1446
rect -38 1390 18 1446
rect 86 1390 142 1446
rect 210 1390 266 1446
rect -286 1266 -230 1322
rect -162 1266 -106 1322
rect -38 1266 18 1322
rect 86 1266 142 1322
rect 210 1266 266 1322
rect -286 1142 -230 1198
rect -162 1142 -106 1198
rect -38 1142 18 1198
rect 86 1142 142 1198
rect 210 1142 266 1198
rect -286 1018 -230 1074
rect -162 1018 -106 1074
rect -38 1018 18 1074
rect 86 1018 142 1074
rect 210 1018 266 1074
rect -286 894 -230 950
rect -162 894 -106 950
rect -38 894 18 950
rect 86 894 142 950
rect 210 894 266 950
rect -286 770 -230 826
rect -162 770 -106 826
rect -38 770 18 826
rect 86 770 142 826
rect 210 770 266 826
rect -286 646 -230 702
rect -162 646 -106 702
rect -38 646 18 702
rect 86 646 142 702
rect 210 646 266 702
rect -286 522 -230 578
rect -162 522 -106 578
rect -38 522 18 578
rect 86 522 142 578
rect 210 522 266 578
rect -286 398 -230 454
rect -162 398 -106 454
rect -38 398 18 454
rect 86 398 142 454
rect 210 398 266 454
rect 903 12254 959 12310
rect 1045 12254 1101 12310
rect 903 12112 959 12168
rect 1045 12112 1101 12168
rect 903 11970 959 12026
rect 1045 11970 1101 12026
rect 903 11828 959 11884
rect 1045 11828 1101 11884
rect 903 11686 959 11742
rect 1045 11686 1101 11742
rect 903 11544 959 11600
rect 1045 11544 1101 11600
rect 903 11402 959 11458
rect 1045 11402 1101 11458
rect 903 11260 959 11316
rect 1045 11260 1101 11316
rect 903 11118 959 11174
rect 1045 11118 1101 11174
rect 903 10976 959 11032
rect 1045 10976 1101 11032
rect 903 10834 959 10890
rect 1045 10834 1101 10890
rect 903 10692 959 10748
rect 1045 10692 1101 10748
rect 903 10550 959 10606
rect 1045 10550 1101 10606
rect 903 10408 959 10464
rect 1045 10408 1101 10464
rect 903 10266 959 10322
rect 1045 10266 1101 10322
rect 903 10124 959 10180
rect 1045 10124 1101 10180
rect 903 9982 959 10038
rect 1045 9982 1101 10038
rect 903 9840 959 9896
rect 1045 9840 1101 9896
rect 903 9698 959 9754
rect 1045 9698 1101 9754
rect 903 9556 959 9612
rect 1045 9556 1101 9612
rect 903 9414 959 9470
rect 1045 9414 1101 9470
rect 903 9272 959 9328
rect 1045 9272 1101 9328
rect 903 9130 959 9186
rect 1045 9130 1101 9186
rect 903 8988 959 9044
rect 1045 8988 1101 9044
rect 903 8846 959 8902
rect 1045 8846 1101 8902
rect 903 8704 959 8760
rect 1045 8704 1101 8760
rect 903 8562 959 8618
rect 1045 8562 1101 8618
rect 903 8420 959 8476
rect 1045 8420 1101 8476
rect 903 8278 959 8334
rect 1045 8278 1101 8334
rect 903 8136 959 8192
rect 1045 8136 1101 8192
rect 903 7994 959 8050
rect 1045 7994 1101 8050
rect 903 7852 959 7908
rect 1045 7852 1101 7908
rect 903 7710 959 7766
rect 1045 7710 1101 7766
rect 903 7568 959 7624
rect 1045 7568 1101 7624
rect 903 7426 959 7482
rect 1045 7426 1101 7482
rect 903 7284 959 7340
rect 1045 7284 1101 7340
rect 903 7142 959 7198
rect 1045 7142 1101 7198
rect 903 7000 959 7056
rect 1045 7000 1101 7056
rect 903 6858 959 6914
rect 1045 6858 1101 6914
rect 903 6716 959 6772
rect 1045 6716 1101 6772
rect 903 6574 959 6630
rect 1045 6574 1101 6630
rect 903 6432 959 6488
rect 1045 6432 1101 6488
rect 903 6290 959 6346
rect 1045 6290 1101 6346
rect 903 6148 959 6204
rect 1045 6148 1101 6204
rect 903 6006 959 6062
rect 1045 6006 1101 6062
rect 903 5864 959 5920
rect 1045 5864 1101 5920
rect 903 5722 959 5778
rect 1045 5722 1101 5778
rect 903 5580 959 5636
rect 1045 5580 1101 5636
rect 903 5438 959 5494
rect 1045 5438 1101 5494
rect 903 5296 959 5352
rect 1045 5296 1101 5352
rect 903 5154 959 5210
rect 1045 5154 1101 5210
rect 903 5012 959 5068
rect 1045 5012 1101 5068
rect 903 4870 959 4926
rect 1045 4870 1101 4926
rect 903 4728 959 4784
rect 1045 4728 1101 4784
rect 903 4586 959 4642
rect 1045 4586 1101 4642
rect 903 4444 959 4500
rect 1045 4444 1101 4500
rect 903 4302 959 4358
rect 1045 4302 1101 4358
rect 903 4160 959 4216
rect 1045 4160 1101 4216
rect 903 4018 959 4074
rect 1045 4018 1101 4074
rect 903 3876 959 3932
rect 1045 3876 1101 3932
rect 903 3734 959 3790
rect 1045 3734 1101 3790
rect 903 3592 959 3648
rect 1045 3592 1101 3648
rect 903 3450 959 3506
rect 1045 3450 1101 3506
rect 903 3308 959 3364
rect 1045 3308 1101 3364
rect 903 3166 959 3222
rect 1045 3166 1101 3222
rect 903 3024 959 3080
rect 1045 3024 1101 3080
rect 903 2882 959 2938
rect 1045 2882 1101 2938
rect 903 2740 959 2796
rect 1045 2740 1101 2796
rect 903 2598 959 2654
rect 1045 2598 1101 2654
rect 903 2456 959 2512
rect 1045 2456 1101 2512
rect 903 2314 959 2370
rect 1045 2314 1101 2370
rect 903 2172 959 2228
rect 1045 2172 1101 2228
rect 903 2030 959 2086
rect 1045 2030 1101 2086
rect 903 1888 959 1944
rect 1045 1888 1101 1944
rect 903 1746 959 1802
rect 1045 1746 1101 1802
rect 903 1604 959 1660
rect 1045 1604 1101 1660
rect 903 1462 959 1518
rect 1045 1462 1101 1518
rect 903 1320 959 1376
rect 1045 1320 1101 1376
rect 903 1178 959 1234
rect 1045 1178 1101 1234
rect 903 1036 959 1092
rect 1045 1036 1101 1092
rect 903 894 959 950
rect 1045 894 1101 950
rect 903 752 959 808
rect 1045 752 1101 808
rect 903 610 959 666
rect 1045 610 1101 666
rect 903 468 959 524
rect 1045 468 1101 524
rect 1444 12254 1500 12310
rect 1586 12254 1642 12310
rect 1444 12112 1500 12168
rect 1586 12112 1642 12168
rect 1444 11970 1500 12026
rect 1586 11970 1642 12026
rect 1444 11828 1500 11884
rect 1586 11828 1642 11884
rect 1444 11686 1500 11742
rect 1586 11686 1642 11742
rect 1444 11544 1500 11600
rect 1586 11544 1642 11600
rect 1444 11402 1500 11458
rect 1586 11402 1642 11458
rect 1444 11260 1500 11316
rect 1586 11260 1642 11316
rect 1444 11118 1500 11174
rect 1586 11118 1642 11174
rect 1444 10976 1500 11032
rect 1586 10976 1642 11032
rect 1444 10834 1500 10890
rect 1586 10834 1642 10890
rect 1444 10692 1500 10748
rect 1586 10692 1642 10748
rect 1444 10550 1500 10606
rect 1586 10550 1642 10606
rect 1444 10408 1500 10464
rect 1586 10408 1642 10464
rect 1444 10266 1500 10322
rect 1586 10266 1642 10322
rect 1444 10124 1500 10180
rect 1586 10124 1642 10180
rect 1444 9982 1500 10038
rect 1586 9982 1642 10038
rect 1444 9840 1500 9896
rect 1586 9840 1642 9896
rect 1444 9698 1500 9754
rect 1586 9698 1642 9754
rect 1444 9556 1500 9612
rect 1586 9556 1642 9612
rect 1444 9414 1500 9470
rect 1586 9414 1642 9470
rect 1444 9272 1500 9328
rect 1586 9272 1642 9328
rect 1444 9130 1500 9186
rect 1586 9130 1642 9186
rect 1444 8988 1500 9044
rect 1586 8988 1642 9044
rect 1444 8846 1500 8902
rect 1586 8846 1642 8902
rect 1444 8704 1500 8760
rect 1586 8704 1642 8760
rect 1444 8562 1500 8618
rect 1586 8562 1642 8618
rect 1444 8420 1500 8476
rect 1586 8420 1642 8476
rect 1444 8278 1500 8334
rect 1586 8278 1642 8334
rect 1444 8136 1500 8192
rect 1586 8136 1642 8192
rect 1444 7994 1500 8050
rect 1586 7994 1642 8050
rect 1444 7852 1500 7908
rect 1586 7852 1642 7908
rect 1444 7710 1500 7766
rect 1586 7710 1642 7766
rect 1444 7568 1500 7624
rect 1586 7568 1642 7624
rect 1444 7426 1500 7482
rect 1586 7426 1642 7482
rect 1444 7284 1500 7340
rect 1586 7284 1642 7340
rect 1444 7142 1500 7198
rect 1586 7142 1642 7198
rect 1444 7000 1500 7056
rect 1586 7000 1642 7056
rect 1444 6858 1500 6914
rect 1586 6858 1642 6914
rect 1444 6716 1500 6772
rect 1586 6716 1642 6772
rect 1444 6574 1500 6630
rect 1586 6574 1642 6630
rect 1444 6432 1500 6488
rect 1586 6432 1642 6488
rect 1444 6290 1500 6346
rect 1586 6290 1642 6346
rect 1444 6148 1500 6204
rect 1586 6148 1642 6204
rect 1444 6006 1500 6062
rect 1586 6006 1642 6062
rect 1444 5864 1500 5920
rect 1586 5864 1642 5920
rect 1444 5722 1500 5778
rect 1586 5722 1642 5778
rect 1444 5580 1500 5636
rect 1586 5580 1642 5636
rect 1444 5438 1500 5494
rect 1586 5438 1642 5494
rect 1444 5296 1500 5352
rect 1586 5296 1642 5352
rect 1444 5154 1500 5210
rect 1586 5154 1642 5210
rect 1444 5012 1500 5068
rect 1586 5012 1642 5068
rect 1444 4870 1500 4926
rect 1586 4870 1642 4926
rect 1444 4728 1500 4784
rect 1586 4728 1642 4784
rect 1444 4586 1500 4642
rect 1586 4586 1642 4642
rect 1444 4444 1500 4500
rect 1586 4444 1642 4500
rect 1444 4302 1500 4358
rect 1586 4302 1642 4358
rect 1444 4160 1500 4216
rect 1586 4160 1642 4216
rect 1444 4018 1500 4074
rect 1586 4018 1642 4074
rect 1444 3876 1500 3932
rect 1586 3876 1642 3932
rect 1444 3734 1500 3790
rect 1586 3734 1642 3790
rect 1444 3592 1500 3648
rect 1586 3592 1642 3648
rect 1444 3450 1500 3506
rect 1586 3450 1642 3506
rect 1444 3308 1500 3364
rect 1586 3308 1642 3364
rect 1444 3166 1500 3222
rect 1586 3166 1642 3222
rect 1444 3024 1500 3080
rect 1586 3024 1642 3080
rect 1444 2882 1500 2938
rect 1586 2882 1642 2938
rect 1444 2740 1500 2796
rect 1586 2740 1642 2796
rect 1444 2598 1500 2654
rect 1586 2598 1642 2654
rect 1444 2456 1500 2512
rect 1586 2456 1642 2512
rect 1444 2314 1500 2370
rect 1586 2314 1642 2370
rect 1444 2172 1500 2228
rect 1586 2172 1642 2228
rect 1444 2030 1500 2086
rect 1586 2030 1642 2086
rect 1444 1888 1500 1944
rect 1586 1888 1642 1944
rect 1444 1746 1500 1802
rect 1586 1746 1642 1802
rect 1444 1604 1500 1660
rect 1586 1604 1642 1660
rect 1444 1462 1500 1518
rect 1586 1462 1642 1518
rect 1444 1320 1500 1376
rect 1586 1320 1642 1376
rect 1444 1178 1500 1234
rect 1586 1178 1642 1234
rect 1444 1036 1500 1092
rect 1586 1036 1642 1092
rect 1444 894 1500 950
rect 1586 894 1642 950
rect 1444 752 1500 808
rect 1586 752 1642 808
rect 1444 610 1500 666
rect 1586 610 1642 666
rect 1444 468 1500 524
rect 1586 468 1642 524
rect 1984 12254 2040 12310
rect 2126 12254 2182 12310
rect 1984 12112 2040 12168
rect 2126 12112 2182 12168
rect 1984 11970 2040 12026
rect 2126 11970 2182 12026
rect 1984 11828 2040 11884
rect 2126 11828 2182 11884
rect 1984 11686 2040 11742
rect 2126 11686 2182 11742
rect 1984 11544 2040 11600
rect 2126 11544 2182 11600
rect 1984 11402 2040 11458
rect 2126 11402 2182 11458
rect 1984 11260 2040 11316
rect 2126 11260 2182 11316
rect 1984 11118 2040 11174
rect 2126 11118 2182 11174
rect 1984 10976 2040 11032
rect 2126 10976 2182 11032
rect 1984 10834 2040 10890
rect 2126 10834 2182 10890
rect 1984 10692 2040 10748
rect 2126 10692 2182 10748
rect 1984 10550 2040 10606
rect 2126 10550 2182 10606
rect 1984 10408 2040 10464
rect 2126 10408 2182 10464
rect 1984 10266 2040 10322
rect 2126 10266 2182 10322
rect 1984 10124 2040 10180
rect 2126 10124 2182 10180
rect 1984 9982 2040 10038
rect 2126 9982 2182 10038
rect 1984 9840 2040 9896
rect 2126 9840 2182 9896
rect 1984 9698 2040 9754
rect 2126 9698 2182 9754
rect 1984 9556 2040 9612
rect 2126 9556 2182 9612
rect 1984 9414 2040 9470
rect 2126 9414 2182 9470
rect 1984 9272 2040 9328
rect 2126 9272 2182 9328
rect 1984 9130 2040 9186
rect 2126 9130 2182 9186
rect 1984 8988 2040 9044
rect 2126 8988 2182 9044
rect 1984 8846 2040 8902
rect 2126 8846 2182 8902
rect 1984 8704 2040 8760
rect 2126 8704 2182 8760
rect 1984 8562 2040 8618
rect 2126 8562 2182 8618
rect 1984 8420 2040 8476
rect 2126 8420 2182 8476
rect 1984 8278 2040 8334
rect 2126 8278 2182 8334
rect 1984 8136 2040 8192
rect 2126 8136 2182 8192
rect 1984 7994 2040 8050
rect 2126 7994 2182 8050
rect 1984 7852 2040 7908
rect 2126 7852 2182 7908
rect 1984 7710 2040 7766
rect 2126 7710 2182 7766
rect 1984 7568 2040 7624
rect 2126 7568 2182 7624
rect 1984 7426 2040 7482
rect 2126 7426 2182 7482
rect 1984 7284 2040 7340
rect 2126 7284 2182 7340
rect 1984 7142 2040 7198
rect 2126 7142 2182 7198
rect 1984 7000 2040 7056
rect 2126 7000 2182 7056
rect 1984 6858 2040 6914
rect 2126 6858 2182 6914
rect 1984 6716 2040 6772
rect 2126 6716 2182 6772
rect 1984 6574 2040 6630
rect 2126 6574 2182 6630
rect 1984 6432 2040 6488
rect 2126 6432 2182 6488
rect 1984 6290 2040 6346
rect 2126 6290 2182 6346
rect 1984 6148 2040 6204
rect 2126 6148 2182 6204
rect 1984 6006 2040 6062
rect 2126 6006 2182 6062
rect 1984 5864 2040 5920
rect 2126 5864 2182 5920
rect 1984 5722 2040 5778
rect 2126 5722 2182 5778
rect 1984 5580 2040 5636
rect 2126 5580 2182 5636
rect 1984 5438 2040 5494
rect 2126 5438 2182 5494
rect 1984 5296 2040 5352
rect 2126 5296 2182 5352
rect 1984 5154 2040 5210
rect 2126 5154 2182 5210
rect 1984 5012 2040 5068
rect 2126 5012 2182 5068
rect 1984 4870 2040 4926
rect 2126 4870 2182 4926
rect 1984 4728 2040 4784
rect 2126 4728 2182 4784
rect 1984 4586 2040 4642
rect 2126 4586 2182 4642
rect 1984 4444 2040 4500
rect 2126 4444 2182 4500
rect 1984 4302 2040 4358
rect 2126 4302 2182 4358
rect 1984 4160 2040 4216
rect 2126 4160 2182 4216
rect 1984 4018 2040 4074
rect 2126 4018 2182 4074
rect 1984 3876 2040 3932
rect 2126 3876 2182 3932
rect 1984 3734 2040 3790
rect 2126 3734 2182 3790
rect 1984 3592 2040 3648
rect 2126 3592 2182 3648
rect 1984 3450 2040 3506
rect 2126 3450 2182 3506
rect 1984 3308 2040 3364
rect 2126 3308 2182 3364
rect 1984 3166 2040 3222
rect 2126 3166 2182 3222
rect 1984 3024 2040 3080
rect 2126 3024 2182 3080
rect 1984 2882 2040 2938
rect 2126 2882 2182 2938
rect 1984 2740 2040 2796
rect 2126 2740 2182 2796
rect 1984 2598 2040 2654
rect 2126 2598 2182 2654
rect 1984 2456 2040 2512
rect 2126 2456 2182 2512
rect 1984 2314 2040 2370
rect 2126 2314 2182 2370
rect 1984 2172 2040 2228
rect 2126 2172 2182 2228
rect 1984 2030 2040 2086
rect 2126 2030 2182 2086
rect 1984 1888 2040 1944
rect 2126 1888 2182 1944
rect 1984 1746 2040 1802
rect 2126 1746 2182 1802
rect 1984 1604 2040 1660
rect 2126 1604 2182 1660
rect 1984 1462 2040 1518
rect 2126 1462 2182 1518
rect 1984 1320 2040 1376
rect 2126 1320 2182 1376
rect 1984 1178 2040 1234
rect 2126 1178 2182 1234
rect 1984 1036 2040 1092
rect 2126 1036 2182 1092
rect 1984 894 2040 950
rect 2126 894 2182 950
rect 1984 752 2040 808
rect 2126 752 2182 808
rect 1984 610 2040 666
rect 2126 610 2182 666
rect 1984 468 2040 524
rect 2126 468 2182 524
rect 2521 12254 2577 12310
rect 2663 12254 2719 12310
rect 2521 12112 2577 12168
rect 2663 12112 2719 12168
rect 2521 11970 2577 12026
rect 2663 11970 2719 12026
rect 2521 11828 2577 11884
rect 2663 11828 2719 11884
rect 2521 11686 2577 11742
rect 2663 11686 2719 11742
rect 2521 11544 2577 11600
rect 2663 11544 2719 11600
rect 2521 11402 2577 11458
rect 2663 11402 2719 11458
rect 2521 11260 2577 11316
rect 2663 11260 2719 11316
rect 2521 11118 2577 11174
rect 2663 11118 2719 11174
rect 2521 10976 2577 11032
rect 2663 10976 2719 11032
rect 2521 10834 2577 10890
rect 2663 10834 2719 10890
rect 2521 10692 2577 10748
rect 2663 10692 2719 10748
rect 2521 10550 2577 10606
rect 2663 10550 2719 10606
rect 2521 10408 2577 10464
rect 2663 10408 2719 10464
rect 2521 10266 2577 10322
rect 2663 10266 2719 10322
rect 2521 10124 2577 10180
rect 2663 10124 2719 10180
rect 2521 9982 2577 10038
rect 2663 9982 2719 10038
rect 2521 9840 2577 9896
rect 2663 9840 2719 9896
rect 2521 9698 2577 9754
rect 2663 9698 2719 9754
rect 2521 9556 2577 9612
rect 2663 9556 2719 9612
rect 2521 9414 2577 9470
rect 2663 9414 2719 9470
rect 2521 9272 2577 9328
rect 2663 9272 2719 9328
rect 2521 9130 2577 9186
rect 2663 9130 2719 9186
rect 2521 8988 2577 9044
rect 2663 8988 2719 9044
rect 2521 8846 2577 8902
rect 2663 8846 2719 8902
rect 2521 8704 2577 8760
rect 2663 8704 2719 8760
rect 2521 8562 2577 8618
rect 2663 8562 2719 8618
rect 2521 8420 2577 8476
rect 2663 8420 2719 8476
rect 2521 8278 2577 8334
rect 2663 8278 2719 8334
rect 2521 8136 2577 8192
rect 2663 8136 2719 8192
rect 2521 7994 2577 8050
rect 2663 7994 2719 8050
rect 2521 7852 2577 7908
rect 2663 7852 2719 7908
rect 2521 7710 2577 7766
rect 2663 7710 2719 7766
rect 2521 7568 2577 7624
rect 2663 7568 2719 7624
rect 2521 7426 2577 7482
rect 2663 7426 2719 7482
rect 2521 7284 2577 7340
rect 2663 7284 2719 7340
rect 2521 7142 2577 7198
rect 2663 7142 2719 7198
rect 2521 7000 2577 7056
rect 2663 7000 2719 7056
rect 2521 6858 2577 6914
rect 2663 6858 2719 6914
rect 2521 6716 2577 6772
rect 2663 6716 2719 6772
rect 2521 6574 2577 6630
rect 2663 6574 2719 6630
rect 2521 6432 2577 6488
rect 2663 6432 2719 6488
rect 2521 6290 2577 6346
rect 2663 6290 2719 6346
rect 2521 6148 2577 6204
rect 2663 6148 2719 6204
rect 2521 6006 2577 6062
rect 2663 6006 2719 6062
rect 2521 5864 2577 5920
rect 2663 5864 2719 5920
rect 2521 5722 2577 5778
rect 2663 5722 2719 5778
rect 2521 5580 2577 5636
rect 2663 5580 2719 5636
rect 2521 5438 2577 5494
rect 2663 5438 2719 5494
rect 2521 5296 2577 5352
rect 2663 5296 2719 5352
rect 2521 5154 2577 5210
rect 2663 5154 2719 5210
rect 2521 5012 2577 5068
rect 2663 5012 2719 5068
rect 2521 4870 2577 4926
rect 2663 4870 2719 4926
rect 2521 4728 2577 4784
rect 2663 4728 2719 4784
rect 2521 4586 2577 4642
rect 2663 4586 2719 4642
rect 2521 4444 2577 4500
rect 2663 4444 2719 4500
rect 2521 4302 2577 4358
rect 2663 4302 2719 4358
rect 2521 4160 2577 4216
rect 2663 4160 2719 4216
rect 2521 4018 2577 4074
rect 2663 4018 2719 4074
rect 2521 3876 2577 3932
rect 2663 3876 2719 3932
rect 2521 3734 2577 3790
rect 2663 3734 2719 3790
rect 2521 3592 2577 3648
rect 2663 3592 2719 3648
rect 2521 3450 2577 3506
rect 2663 3450 2719 3506
rect 2521 3308 2577 3364
rect 2663 3308 2719 3364
rect 2521 3166 2577 3222
rect 2663 3166 2719 3222
rect 2521 3024 2577 3080
rect 2663 3024 2719 3080
rect 2521 2882 2577 2938
rect 2663 2882 2719 2938
rect 2521 2740 2577 2796
rect 2663 2740 2719 2796
rect 2521 2598 2577 2654
rect 2663 2598 2719 2654
rect 2521 2456 2577 2512
rect 2663 2456 2719 2512
rect 2521 2314 2577 2370
rect 2663 2314 2719 2370
rect 2521 2172 2577 2228
rect 2663 2172 2719 2228
rect 2521 2030 2577 2086
rect 2663 2030 2719 2086
rect 2521 1888 2577 1944
rect 2663 1888 2719 1944
rect 2521 1746 2577 1802
rect 2663 1746 2719 1802
rect 2521 1604 2577 1660
rect 2663 1604 2719 1660
rect 2521 1462 2577 1518
rect 2663 1462 2719 1518
rect 2521 1320 2577 1376
rect 2663 1320 2719 1376
rect 2521 1178 2577 1234
rect 2663 1178 2719 1234
rect 2521 1036 2577 1092
rect 2663 1036 2719 1092
rect 2521 894 2577 950
rect 2663 894 2719 950
rect 2521 752 2577 808
rect 2663 752 2719 808
rect 2521 610 2577 666
rect 2663 610 2719 666
rect 2521 468 2577 524
rect 2663 468 2719 524
rect 3058 12254 3114 12310
rect 3200 12254 3256 12310
rect 3058 12112 3114 12168
rect 3200 12112 3256 12168
rect 3058 11970 3114 12026
rect 3200 11970 3256 12026
rect 3058 11828 3114 11884
rect 3200 11828 3256 11884
rect 3058 11686 3114 11742
rect 3200 11686 3256 11742
rect 3058 11544 3114 11600
rect 3200 11544 3256 11600
rect 3058 11402 3114 11458
rect 3200 11402 3256 11458
rect 3058 11260 3114 11316
rect 3200 11260 3256 11316
rect 3058 11118 3114 11174
rect 3200 11118 3256 11174
rect 3058 10976 3114 11032
rect 3200 10976 3256 11032
rect 3058 10834 3114 10890
rect 3200 10834 3256 10890
rect 3058 10692 3114 10748
rect 3200 10692 3256 10748
rect 3058 10550 3114 10606
rect 3200 10550 3256 10606
rect 3058 10408 3114 10464
rect 3200 10408 3256 10464
rect 3058 10266 3114 10322
rect 3200 10266 3256 10322
rect 3058 10124 3114 10180
rect 3200 10124 3256 10180
rect 3058 9982 3114 10038
rect 3200 9982 3256 10038
rect 3058 9840 3114 9896
rect 3200 9840 3256 9896
rect 3058 9698 3114 9754
rect 3200 9698 3256 9754
rect 3058 9556 3114 9612
rect 3200 9556 3256 9612
rect 3058 9414 3114 9470
rect 3200 9414 3256 9470
rect 3058 9272 3114 9328
rect 3200 9272 3256 9328
rect 3058 9130 3114 9186
rect 3200 9130 3256 9186
rect 3058 8988 3114 9044
rect 3200 8988 3256 9044
rect 3058 8846 3114 8902
rect 3200 8846 3256 8902
rect 3058 8704 3114 8760
rect 3200 8704 3256 8760
rect 3058 8562 3114 8618
rect 3200 8562 3256 8618
rect 3058 8420 3114 8476
rect 3200 8420 3256 8476
rect 3058 8278 3114 8334
rect 3200 8278 3256 8334
rect 3058 8136 3114 8192
rect 3200 8136 3256 8192
rect 3058 7994 3114 8050
rect 3200 7994 3256 8050
rect 3058 7852 3114 7908
rect 3200 7852 3256 7908
rect 3058 7710 3114 7766
rect 3200 7710 3256 7766
rect 3058 7568 3114 7624
rect 3200 7568 3256 7624
rect 3058 7426 3114 7482
rect 3200 7426 3256 7482
rect 3058 7284 3114 7340
rect 3200 7284 3256 7340
rect 3058 7142 3114 7198
rect 3200 7142 3256 7198
rect 3058 7000 3114 7056
rect 3200 7000 3256 7056
rect 3058 6858 3114 6914
rect 3200 6858 3256 6914
rect 3058 6716 3114 6772
rect 3200 6716 3256 6772
rect 3058 6574 3114 6630
rect 3200 6574 3256 6630
rect 3058 6432 3114 6488
rect 3200 6432 3256 6488
rect 3058 6290 3114 6346
rect 3200 6290 3256 6346
rect 3058 6148 3114 6204
rect 3200 6148 3256 6204
rect 3058 6006 3114 6062
rect 3200 6006 3256 6062
rect 3058 5864 3114 5920
rect 3200 5864 3256 5920
rect 3058 5722 3114 5778
rect 3200 5722 3256 5778
rect 3058 5580 3114 5636
rect 3200 5580 3256 5636
rect 3058 5438 3114 5494
rect 3200 5438 3256 5494
rect 3058 5296 3114 5352
rect 3200 5296 3256 5352
rect 3058 5154 3114 5210
rect 3200 5154 3256 5210
rect 3058 5012 3114 5068
rect 3200 5012 3256 5068
rect 3058 4870 3114 4926
rect 3200 4870 3256 4926
rect 3058 4728 3114 4784
rect 3200 4728 3256 4784
rect 3058 4586 3114 4642
rect 3200 4586 3256 4642
rect 3058 4444 3114 4500
rect 3200 4444 3256 4500
rect 3058 4302 3114 4358
rect 3200 4302 3256 4358
rect 3058 4160 3114 4216
rect 3200 4160 3256 4216
rect 3058 4018 3114 4074
rect 3200 4018 3256 4074
rect 3058 3876 3114 3932
rect 3200 3876 3256 3932
rect 3058 3734 3114 3790
rect 3200 3734 3256 3790
rect 3058 3592 3114 3648
rect 3200 3592 3256 3648
rect 3058 3450 3114 3506
rect 3200 3450 3256 3506
rect 3058 3308 3114 3364
rect 3200 3308 3256 3364
rect 3058 3166 3114 3222
rect 3200 3166 3256 3222
rect 3058 3024 3114 3080
rect 3200 3024 3256 3080
rect 3058 2882 3114 2938
rect 3200 2882 3256 2938
rect 3058 2740 3114 2796
rect 3200 2740 3256 2796
rect 3058 2598 3114 2654
rect 3200 2598 3256 2654
rect 3058 2456 3114 2512
rect 3200 2456 3256 2512
rect 3058 2314 3114 2370
rect 3200 2314 3256 2370
rect 3058 2172 3114 2228
rect 3200 2172 3256 2228
rect 3058 2030 3114 2086
rect 3200 2030 3256 2086
rect 3058 1888 3114 1944
rect 3200 1888 3256 1944
rect 3058 1746 3114 1802
rect 3200 1746 3256 1802
rect 3058 1604 3114 1660
rect 3200 1604 3256 1660
rect 3058 1462 3114 1518
rect 3200 1462 3256 1518
rect 3058 1320 3114 1376
rect 3200 1320 3256 1376
rect 3058 1178 3114 1234
rect 3200 1178 3256 1234
rect 3058 1036 3114 1092
rect 3200 1036 3256 1092
rect 3058 894 3114 950
rect 3200 894 3256 950
rect 3058 752 3114 808
rect 3200 752 3256 808
rect 3058 610 3114 666
rect 3200 610 3256 666
rect 3058 468 3114 524
rect 3200 468 3256 524
rect 3602 12254 3658 12310
rect 3744 12254 3800 12310
rect 3602 12112 3658 12168
rect 3744 12112 3800 12168
rect 3602 11970 3658 12026
rect 3744 11970 3800 12026
rect 3602 11828 3658 11884
rect 3744 11828 3800 11884
rect 3602 11686 3658 11742
rect 3744 11686 3800 11742
rect 3602 11544 3658 11600
rect 3744 11544 3800 11600
rect 3602 11402 3658 11458
rect 3744 11402 3800 11458
rect 3602 11260 3658 11316
rect 3744 11260 3800 11316
rect 3602 11118 3658 11174
rect 3744 11118 3800 11174
rect 3602 10976 3658 11032
rect 3744 10976 3800 11032
rect 3602 10834 3658 10890
rect 3744 10834 3800 10890
rect 3602 10692 3658 10748
rect 3744 10692 3800 10748
rect 3602 10550 3658 10606
rect 3744 10550 3800 10606
rect 3602 10408 3658 10464
rect 3744 10408 3800 10464
rect 3602 10266 3658 10322
rect 3744 10266 3800 10322
rect 3602 10124 3658 10180
rect 3744 10124 3800 10180
rect 3602 9982 3658 10038
rect 3744 9982 3800 10038
rect 3602 9840 3658 9896
rect 3744 9840 3800 9896
rect 3602 9698 3658 9754
rect 3744 9698 3800 9754
rect 3602 9556 3658 9612
rect 3744 9556 3800 9612
rect 3602 9414 3658 9470
rect 3744 9414 3800 9470
rect 3602 9272 3658 9328
rect 3744 9272 3800 9328
rect 3602 9130 3658 9186
rect 3744 9130 3800 9186
rect 3602 8988 3658 9044
rect 3744 8988 3800 9044
rect 3602 8846 3658 8902
rect 3744 8846 3800 8902
rect 3602 8704 3658 8760
rect 3744 8704 3800 8760
rect 3602 8562 3658 8618
rect 3744 8562 3800 8618
rect 3602 8420 3658 8476
rect 3744 8420 3800 8476
rect 3602 8278 3658 8334
rect 3744 8278 3800 8334
rect 3602 8136 3658 8192
rect 3744 8136 3800 8192
rect 3602 7994 3658 8050
rect 3744 7994 3800 8050
rect 3602 7852 3658 7908
rect 3744 7852 3800 7908
rect 3602 7710 3658 7766
rect 3744 7710 3800 7766
rect 3602 7568 3658 7624
rect 3744 7568 3800 7624
rect 3602 7426 3658 7482
rect 3744 7426 3800 7482
rect 3602 7284 3658 7340
rect 3744 7284 3800 7340
rect 3602 7142 3658 7198
rect 3744 7142 3800 7198
rect 3602 7000 3658 7056
rect 3744 7000 3800 7056
rect 3602 6858 3658 6914
rect 3744 6858 3800 6914
rect 3602 6716 3658 6772
rect 3744 6716 3800 6772
rect 3602 6574 3658 6630
rect 3744 6574 3800 6630
rect 3602 6432 3658 6488
rect 3744 6432 3800 6488
rect 3602 6290 3658 6346
rect 3744 6290 3800 6346
rect 3602 6148 3658 6204
rect 3744 6148 3800 6204
rect 3602 6006 3658 6062
rect 3744 6006 3800 6062
rect 3602 5864 3658 5920
rect 3744 5864 3800 5920
rect 3602 5722 3658 5778
rect 3744 5722 3800 5778
rect 3602 5580 3658 5636
rect 3744 5580 3800 5636
rect 3602 5438 3658 5494
rect 3744 5438 3800 5494
rect 3602 5296 3658 5352
rect 3744 5296 3800 5352
rect 3602 5154 3658 5210
rect 3744 5154 3800 5210
rect 3602 5012 3658 5068
rect 3744 5012 3800 5068
rect 3602 4870 3658 4926
rect 3744 4870 3800 4926
rect 3602 4728 3658 4784
rect 3744 4728 3800 4784
rect 3602 4586 3658 4642
rect 3744 4586 3800 4642
rect 3602 4444 3658 4500
rect 3744 4444 3800 4500
rect 3602 4302 3658 4358
rect 3744 4302 3800 4358
rect 3602 4160 3658 4216
rect 3744 4160 3800 4216
rect 3602 4018 3658 4074
rect 3744 4018 3800 4074
rect 3602 3876 3658 3932
rect 3744 3876 3800 3932
rect 3602 3734 3658 3790
rect 3744 3734 3800 3790
rect 3602 3592 3658 3648
rect 3744 3592 3800 3648
rect 3602 3450 3658 3506
rect 3744 3450 3800 3506
rect 3602 3308 3658 3364
rect 3744 3308 3800 3364
rect 3602 3166 3658 3222
rect 3744 3166 3800 3222
rect 3602 3024 3658 3080
rect 3744 3024 3800 3080
rect 3602 2882 3658 2938
rect 3744 2882 3800 2938
rect 3602 2740 3658 2796
rect 3744 2740 3800 2796
rect 3602 2598 3658 2654
rect 3744 2598 3800 2654
rect 3602 2456 3658 2512
rect 3744 2456 3800 2512
rect 3602 2314 3658 2370
rect 3744 2314 3800 2370
rect 3602 2172 3658 2228
rect 3744 2172 3800 2228
rect 3602 2030 3658 2086
rect 3744 2030 3800 2086
rect 3602 1888 3658 1944
rect 3744 1888 3800 1944
rect 3602 1746 3658 1802
rect 3744 1746 3800 1802
rect 3602 1604 3658 1660
rect 3744 1604 3800 1660
rect 3602 1462 3658 1518
rect 3744 1462 3800 1518
rect 3602 1320 3658 1376
rect 3744 1320 3800 1376
rect 3602 1178 3658 1234
rect 3744 1178 3800 1234
rect 3602 1036 3658 1092
rect 3744 1036 3800 1092
rect 3602 894 3658 950
rect 3744 894 3800 950
rect 3602 752 3658 808
rect 3744 752 3800 808
rect 3602 610 3658 666
rect 3744 610 3800 666
rect 3602 468 3658 524
rect 3744 468 3800 524
rect 4138 12254 4194 12310
rect 4280 12254 4336 12310
rect 4138 12112 4194 12168
rect 4280 12112 4336 12168
rect 4138 11970 4194 12026
rect 4280 11970 4336 12026
rect 4138 11828 4194 11884
rect 4280 11828 4336 11884
rect 4138 11686 4194 11742
rect 4280 11686 4336 11742
rect 4138 11544 4194 11600
rect 4280 11544 4336 11600
rect 4138 11402 4194 11458
rect 4280 11402 4336 11458
rect 4138 11260 4194 11316
rect 4280 11260 4336 11316
rect 4138 11118 4194 11174
rect 4280 11118 4336 11174
rect 4138 10976 4194 11032
rect 4280 10976 4336 11032
rect 4138 10834 4194 10890
rect 4280 10834 4336 10890
rect 4138 10692 4194 10748
rect 4280 10692 4336 10748
rect 4138 10550 4194 10606
rect 4280 10550 4336 10606
rect 4138 10408 4194 10464
rect 4280 10408 4336 10464
rect 4138 10266 4194 10322
rect 4280 10266 4336 10322
rect 4138 10124 4194 10180
rect 4280 10124 4336 10180
rect 4138 9982 4194 10038
rect 4280 9982 4336 10038
rect 4138 9840 4194 9896
rect 4280 9840 4336 9896
rect 4138 9698 4194 9754
rect 4280 9698 4336 9754
rect 4138 9556 4194 9612
rect 4280 9556 4336 9612
rect 4138 9414 4194 9470
rect 4280 9414 4336 9470
rect 4138 9272 4194 9328
rect 4280 9272 4336 9328
rect 4138 9130 4194 9186
rect 4280 9130 4336 9186
rect 4138 8988 4194 9044
rect 4280 8988 4336 9044
rect 4138 8846 4194 8902
rect 4280 8846 4336 8902
rect 4138 8704 4194 8760
rect 4280 8704 4336 8760
rect 4138 8562 4194 8618
rect 4280 8562 4336 8618
rect 4138 8420 4194 8476
rect 4280 8420 4336 8476
rect 4138 8278 4194 8334
rect 4280 8278 4336 8334
rect 4138 8136 4194 8192
rect 4280 8136 4336 8192
rect 4138 7994 4194 8050
rect 4280 7994 4336 8050
rect 4138 7852 4194 7908
rect 4280 7852 4336 7908
rect 4138 7710 4194 7766
rect 4280 7710 4336 7766
rect 4138 7568 4194 7624
rect 4280 7568 4336 7624
rect 4138 7426 4194 7482
rect 4280 7426 4336 7482
rect 4138 7284 4194 7340
rect 4280 7284 4336 7340
rect 4138 7142 4194 7198
rect 4280 7142 4336 7198
rect 4138 7000 4194 7056
rect 4280 7000 4336 7056
rect 4138 6858 4194 6914
rect 4280 6858 4336 6914
rect 4138 6716 4194 6772
rect 4280 6716 4336 6772
rect 4138 6574 4194 6630
rect 4280 6574 4336 6630
rect 4138 6432 4194 6488
rect 4280 6432 4336 6488
rect 4138 6290 4194 6346
rect 4280 6290 4336 6346
rect 4138 6148 4194 6204
rect 4280 6148 4336 6204
rect 4138 6006 4194 6062
rect 4280 6006 4336 6062
rect 4138 5864 4194 5920
rect 4280 5864 4336 5920
rect 4138 5722 4194 5778
rect 4280 5722 4336 5778
rect 4138 5580 4194 5636
rect 4280 5580 4336 5636
rect 4138 5438 4194 5494
rect 4280 5438 4336 5494
rect 4138 5296 4194 5352
rect 4280 5296 4336 5352
rect 4138 5154 4194 5210
rect 4280 5154 4336 5210
rect 4138 5012 4194 5068
rect 4280 5012 4336 5068
rect 4138 4870 4194 4926
rect 4280 4870 4336 4926
rect 4138 4728 4194 4784
rect 4280 4728 4336 4784
rect 4138 4586 4194 4642
rect 4280 4586 4336 4642
rect 4138 4444 4194 4500
rect 4280 4444 4336 4500
rect 4138 4302 4194 4358
rect 4280 4302 4336 4358
rect 4138 4160 4194 4216
rect 4280 4160 4336 4216
rect 4138 4018 4194 4074
rect 4280 4018 4336 4074
rect 4138 3876 4194 3932
rect 4280 3876 4336 3932
rect 4138 3734 4194 3790
rect 4280 3734 4336 3790
rect 4138 3592 4194 3648
rect 4280 3592 4336 3648
rect 4138 3450 4194 3506
rect 4280 3450 4336 3506
rect 4138 3308 4194 3364
rect 4280 3308 4336 3364
rect 4138 3166 4194 3222
rect 4280 3166 4336 3222
rect 4138 3024 4194 3080
rect 4280 3024 4336 3080
rect 4138 2882 4194 2938
rect 4280 2882 4336 2938
rect 4138 2740 4194 2796
rect 4280 2740 4336 2796
rect 4138 2598 4194 2654
rect 4280 2598 4336 2654
rect 4138 2456 4194 2512
rect 4280 2456 4336 2512
rect 4138 2314 4194 2370
rect 4280 2314 4336 2370
rect 4138 2172 4194 2228
rect 4280 2172 4336 2228
rect 4138 2030 4194 2086
rect 4280 2030 4336 2086
rect 4138 1888 4194 1944
rect 4280 1888 4336 1944
rect 4138 1746 4194 1802
rect 4280 1746 4336 1802
rect 4138 1604 4194 1660
rect 4280 1604 4336 1660
rect 4138 1462 4194 1518
rect 4280 1462 4336 1518
rect 4138 1320 4194 1376
rect 4280 1320 4336 1376
rect 4138 1178 4194 1234
rect 4280 1178 4336 1234
rect 4138 1036 4194 1092
rect 4280 1036 4336 1092
rect 4138 894 4194 950
rect 4280 894 4336 950
rect 4138 752 4194 808
rect 4280 752 4336 808
rect 4138 610 4194 666
rect 4280 610 4336 666
rect 4138 468 4194 524
rect 4280 468 4336 524
rect 4678 12254 4734 12310
rect 4820 12254 4876 12310
rect 4678 12112 4734 12168
rect 4820 12112 4876 12168
rect 4678 11970 4734 12026
rect 4820 11970 4876 12026
rect 4678 11828 4734 11884
rect 4820 11828 4876 11884
rect 4678 11686 4734 11742
rect 4820 11686 4876 11742
rect 4678 11544 4734 11600
rect 4820 11544 4876 11600
rect 4678 11402 4734 11458
rect 4820 11402 4876 11458
rect 4678 11260 4734 11316
rect 4820 11260 4876 11316
rect 4678 11118 4734 11174
rect 4820 11118 4876 11174
rect 4678 10976 4734 11032
rect 4820 10976 4876 11032
rect 4678 10834 4734 10890
rect 4820 10834 4876 10890
rect 4678 10692 4734 10748
rect 4820 10692 4876 10748
rect 4678 10550 4734 10606
rect 4820 10550 4876 10606
rect 4678 10408 4734 10464
rect 4820 10408 4876 10464
rect 4678 10266 4734 10322
rect 4820 10266 4876 10322
rect 4678 10124 4734 10180
rect 4820 10124 4876 10180
rect 4678 9982 4734 10038
rect 4820 9982 4876 10038
rect 4678 9840 4734 9896
rect 4820 9840 4876 9896
rect 4678 9698 4734 9754
rect 4820 9698 4876 9754
rect 4678 9556 4734 9612
rect 4820 9556 4876 9612
rect 4678 9414 4734 9470
rect 4820 9414 4876 9470
rect 4678 9272 4734 9328
rect 4820 9272 4876 9328
rect 4678 9130 4734 9186
rect 4820 9130 4876 9186
rect 4678 8988 4734 9044
rect 4820 8988 4876 9044
rect 4678 8846 4734 8902
rect 4820 8846 4876 8902
rect 4678 8704 4734 8760
rect 4820 8704 4876 8760
rect 4678 8562 4734 8618
rect 4820 8562 4876 8618
rect 4678 8420 4734 8476
rect 4820 8420 4876 8476
rect 4678 8278 4734 8334
rect 4820 8278 4876 8334
rect 4678 8136 4734 8192
rect 4820 8136 4876 8192
rect 4678 7994 4734 8050
rect 4820 7994 4876 8050
rect 4678 7852 4734 7908
rect 4820 7852 4876 7908
rect 4678 7710 4734 7766
rect 4820 7710 4876 7766
rect 4678 7568 4734 7624
rect 4820 7568 4876 7624
rect 4678 7426 4734 7482
rect 4820 7426 4876 7482
rect 4678 7284 4734 7340
rect 4820 7284 4876 7340
rect 4678 7142 4734 7198
rect 4820 7142 4876 7198
rect 4678 7000 4734 7056
rect 4820 7000 4876 7056
rect 4678 6858 4734 6914
rect 4820 6858 4876 6914
rect 4678 6716 4734 6772
rect 4820 6716 4876 6772
rect 4678 6574 4734 6630
rect 4820 6574 4876 6630
rect 4678 6432 4734 6488
rect 4820 6432 4876 6488
rect 4678 6290 4734 6346
rect 4820 6290 4876 6346
rect 4678 6148 4734 6204
rect 4820 6148 4876 6204
rect 4678 6006 4734 6062
rect 4820 6006 4876 6062
rect 4678 5864 4734 5920
rect 4820 5864 4876 5920
rect 4678 5722 4734 5778
rect 4820 5722 4876 5778
rect 4678 5580 4734 5636
rect 4820 5580 4876 5636
rect 4678 5438 4734 5494
rect 4820 5438 4876 5494
rect 4678 5296 4734 5352
rect 4820 5296 4876 5352
rect 4678 5154 4734 5210
rect 4820 5154 4876 5210
rect 4678 5012 4734 5068
rect 4820 5012 4876 5068
rect 4678 4870 4734 4926
rect 4820 4870 4876 4926
rect 4678 4728 4734 4784
rect 4820 4728 4876 4784
rect 4678 4586 4734 4642
rect 4820 4586 4876 4642
rect 4678 4444 4734 4500
rect 4820 4444 4876 4500
rect 4678 4302 4734 4358
rect 4820 4302 4876 4358
rect 4678 4160 4734 4216
rect 4820 4160 4876 4216
rect 4678 4018 4734 4074
rect 4820 4018 4876 4074
rect 4678 3876 4734 3932
rect 4820 3876 4876 3932
rect 4678 3734 4734 3790
rect 4820 3734 4876 3790
rect 4678 3592 4734 3648
rect 4820 3592 4876 3648
rect 4678 3450 4734 3506
rect 4820 3450 4876 3506
rect 4678 3308 4734 3364
rect 4820 3308 4876 3364
rect 4678 3166 4734 3222
rect 4820 3166 4876 3222
rect 4678 3024 4734 3080
rect 4820 3024 4876 3080
rect 4678 2882 4734 2938
rect 4820 2882 4876 2938
rect 4678 2740 4734 2796
rect 4820 2740 4876 2796
rect 4678 2598 4734 2654
rect 4820 2598 4876 2654
rect 4678 2456 4734 2512
rect 4820 2456 4876 2512
rect 4678 2314 4734 2370
rect 4820 2314 4876 2370
rect 4678 2172 4734 2228
rect 4820 2172 4876 2228
rect 4678 2030 4734 2086
rect 4820 2030 4876 2086
rect 4678 1888 4734 1944
rect 4820 1888 4876 1944
rect 4678 1746 4734 1802
rect 4820 1746 4876 1802
rect 4678 1604 4734 1660
rect 4820 1604 4876 1660
rect 4678 1462 4734 1518
rect 4820 1462 4876 1518
rect 4678 1320 4734 1376
rect 4820 1320 4876 1376
rect 4678 1178 4734 1234
rect 4820 1178 4876 1234
rect 4678 1036 4734 1092
rect 4820 1036 4876 1092
rect 4678 894 4734 950
rect 4820 894 4876 950
rect 4678 752 4734 808
rect 4820 752 4876 808
rect 4678 610 4734 666
rect 4820 610 4876 666
rect 4678 468 4734 524
rect 4820 468 4876 524
rect 5215 12254 5271 12310
rect 5357 12254 5413 12310
rect 5215 12112 5271 12168
rect 5357 12112 5413 12168
rect 5215 11970 5271 12026
rect 5357 11970 5413 12026
rect 5215 11828 5271 11884
rect 5357 11828 5413 11884
rect 5215 11686 5271 11742
rect 5357 11686 5413 11742
rect 5215 11544 5271 11600
rect 5357 11544 5413 11600
rect 5215 11402 5271 11458
rect 5357 11402 5413 11458
rect 5215 11260 5271 11316
rect 5357 11260 5413 11316
rect 5215 11118 5271 11174
rect 5357 11118 5413 11174
rect 5215 10976 5271 11032
rect 5357 10976 5413 11032
rect 5215 10834 5271 10890
rect 5357 10834 5413 10890
rect 5215 10692 5271 10748
rect 5357 10692 5413 10748
rect 5215 10550 5271 10606
rect 5357 10550 5413 10606
rect 5215 10408 5271 10464
rect 5357 10408 5413 10464
rect 5215 10266 5271 10322
rect 5357 10266 5413 10322
rect 5215 10124 5271 10180
rect 5357 10124 5413 10180
rect 5215 9982 5271 10038
rect 5357 9982 5413 10038
rect 5215 9840 5271 9896
rect 5357 9840 5413 9896
rect 5215 9698 5271 9754
rect 5357 9698 5413 9754
rect 5215 9556 5271 9612
rect 5357 9556 5413 9612
rect 5215 9414 5271 9470
rect 5357 9414 5413 9470
rect 5215 9272 5271 9328
rect 5357 9272 5413 9328
rect 5215 9130 5271 9186
rect 5357 9130 5413 9186
rect 5215 8988 5271 9044
rect 5357 8988 5413 9044
rect 5215 8846 5271 8902
rect 5357 8846 5413 8902
rect 5215 8704 5271 8760
rect 5357 8704 5413 8760
rect 5215 8562 5271 8618
rect 5357 8562 5413 8618
rect 5215 8420 5271 8476
rect 5357 8420 5413 8476
rect 5215 8278 5271 8334
rect 5357 8278 5413 8334
rect 5215 8136 5271 8192
rect 5357 8136 5413 8192
rect 5215 7994 5271 8050
rect 5357 7994 5413 8050
rect 5215 7852 5271 7908
rect 5357 7852 5413 7908
rect 5215 7710 5271 7766
rect 5357 7710 5413 7766
rect 5215 7568 5271 7624
rect 5357 7568 5413 7624
rect 5215 7426 5271 7482
rect 5357 7426 5413 7482
rect 5215 7284 5271 7340
rect 5357 7284 5413 7340
rect 5215 7142 5271 7198
rect 5357 7142 5413 7198
rect 5215 7000 5271 7056
rect 5357 7000 5413 7056
rect 5215 6858 5271 6914
rect 5357 6858 5413 6914
rect 5215 6716 5271 6772
rect 5357 6716 5413 6772
rect 5215 6574 5271 6630
rect 5357 6574 5413 6630
rect 5215 6432 5271 6488
rect 5357 6432 5413 6488
rect 5215 6290 5271 6346
rect 5357 6290 5413 6346
rect 5215 6148 5271 6204
rect 5357 6148 5413 6204
rect 5215 6006 5271 6062
rect 5357 6006 5413 6062
rect 5215 5864 5271 5920
rect 5357 5864 5413 5920
rect 5215 5722 5271 5778
rect 5357 5722 5413 5778
rect 5215 5580 5271 5636
rect 5357 5580 5413 5636
rect 5215 5438 5271 5494
rect 5357 5438 5413 5494
rect 5215 5296 5271 5352
rect 5357 5296 5413 5352
rect 5215 5154 5271 5210
rect 5357 5154 5413 5210
rect 5215 5012 5271 5068
rect 5357 5012 5413 5068
rect 5215 4870 5271 4926
rect 5357 4870 5413 4926
rect 5215 4728 5271 4784
rect 5357 4728 5413 4784
rect 5215 4586 5271 4642
rect 5357 4586 5413 4642
rect 5215 4444 5271 4500
rect 5357 4444 5413 4500
rect 5215 4302 5271 4358
rect 5357 4302 5413 4358
rect 5215 4160 5271 4216
rect 5357 4160 5413 4216
rect 5215 4018 5271 4074
rect 5357 4018 5413 4074
rect 5215 3876 5271 3932
rect 5357 3876 5413 3932
rect 5215 3734 5271 3790
rect 5357 3734 5413 3790
rect 5215 3592 5271 3648
rect 5357 3592 5413 3648
rect 5215 3450 5271 3506
rect 5357 3450 5413 3506
rect 5215 3308 5271 3364
rect 5357 3308 5413 3364
rect 5215 3166 5271 3222
rect 5357 3166 5413 3222
rect 5215 3024 5271 3080
rect 5357 3024 5413 3080
rect 5215 2882 5271 2938
rect 5357 2882 5413 2938
rect 5215 2740 5271 2796
rect 5357 2740 5413 2796
rect 5215 2598 5271 2654
rect 5357 2598 5413 2654
rect 5215 2456 5271 2512
rect 5357 2456 5413 2512
rect 5215 2314 5271 2370
rect 5357 2314 5413 2370
rect 5215 2172 5271 2228
rect 5357 2172 5413 2228
rect 5215 2030 5271 2086
rect 5357 2030 5413 2086
rect 5215 1888 5271 1944
rect 5357 1888 5413 1944
rect 5215 1746 5271 1802
rect 5357 1746 5413 1802
rect 5215 1604 5271 1660
rect 5357 1604 5413 1660
rect 5215 1462 5271 1518
rect 5357 1462 5413 1518
rect 5215 1320 5271 1376
rect 5357 1320 5413 1376
rect 5215 1178 5271 1234
rect 5357 1178 5413 1234
rect 5215 1036 5271 1092
rect 5357 1036 5413 1092
rect 5215 894 5271 950
rect 5357 894 5413 950
rect 5215 752 5271 808
rect 5357 752 5413 808
rect 5215 610 5271 666
rect 5357 610 5413 666
rect 5215 468 5271 524
rect 5357 468 5413 524
rect 5760 12254 5816 12310
rect 5902 12254 5958 12310
rect 5760 12112 5816 12168
rect 5902 12112 5958 12168
rect 5760 11970 5816 12026
rect 5902 11970 5958 12026
rect 5760 11828 5816 11884
rect 5902 11828 5958 11884
rect 5760 11686 5816 11742
rect 5902 11686 5958 11742
rect 5760 11544 5816 11600
rect 5902 11544 5958 11600
rect 5760 11402 5816 11458
rect 5902 11402 5958 11458
rect 5760 11260 5816 11316
rect 5902 11260 5958 11316
rect 5760 11118 5816 11174
rect 5902 11118 5958 11174
rect 5760 10976 5816 11032
rect 5902 10976 5958 11032
rect 5760 10834 5816 10890
rect 5902 10834 5958 10890
rect 5760 10692 5816 10748
rect 5902 10692 5958 10748
rect 5760 10550 5816 10606
rect 5902 10550 5958 10606
rect 5760 10408 5816 10464
rect 5902 10408 5958 10464
rect 5760 10266 5816 10322
rect 5902 10266 5958 10322
rect 5760 10124 5816 10180
rect 5902 10124 5958 10180
rect 5760 9982 5816 10038
rect 5902 9982 5958 10038
rect 5760 9840 5816 9896
rect 5902 9840 5958 9896
rect 5760 9698 5816 9754
rect 5902 9698 5958 9754
rect 5760 9556 5816 9612
rect 5902 9556 5958 9612
rect 5760 9414 5816 9470
rect 5902 9414 5958 9470
rect 5760 9272 5816 9328
rect 5902 9272 5958 9328
rect 5760 9130 5816 9186
rect 5902 9130 5958 9186
rect 5760 8988 5816 9044
rect 5902 8988 5958 9044
rect 5760 8846 5816 8902
rect 5902 8846 5958 8902
rect 5760 8704 5816 8760
rect 5902 8704 5958 8760
rect 5760 8562 5816 8618
rect 5902 8562 5958 8618
rect 5760 8420 5816 8476
rect 5902 8420 5958 8476
rect 5760 8278 5816 8334
rect 5902 8278 5958 8334
rect 5760 8136 5816 8192
rect 5902 8136 5958 8192
rect 5760 7994 5816 8050
rect 5902 7994 5958 8050
rect 5760 7852 5816 7908
rect 5902 7852 5958 7908
rect 5760 7710 5816 7766
rect 5902 7710 5958 7766
rect 5760 7568 5816 7624
rect 5902 7568 5958 7624
rect 5760 7426 5816 7482
rect 5902 7426 5958 7482
rect 5760 7284 5816 7340
rect 5902 7284 5958 7340
rect 5760 7142 5816 7198
rect 5902 7142 5958 7198
rect 5760 7000 5816 7056
rect 5902 7000 5958 7056
rect 5760 6858 5816 6914
rect 5902 6858 5958 6914
rect 5760 6716 5816 6772
rect 5902 6716 5958 6772
rect 5760 6574 5816 6630
rect 5902 6574 5958 6630
rect 5760 6432 5816 6488
rect 5902 6432 5958 6488
rect 5760 6290 5816 6346
rect 5902 6290 5958 6346
rect 5760 6148 5816 6204
rect 5902 6148 5958 6204
rect 5760 6006 5816 6062
rect 5902 6006 5958 6062
rect 5760 5864 5816 5920
rect 5902 5864 5958 5920
rect 5760 5722 5816 5778
rect 5902 5722 5958 5778
rect 5760 5580 5816 5636
rect 5902 5580 5958 5636
rect 5760 5438 5816 5494
rect 5902 5438 5958 5494
rect 5760 5296 5816 5352
rect 5902 5296 5958 5352
rect 5760 5154 5816 5210
rect 5902 5154 5958 5210
rect 5760 5012 5816 5068
rect 5902 5012 5958 5068
rect 5760 4870 5816 4926
rect 5902 4870 5958 4926
rect 5760 4728 5816 4784
rect 5902 4728 5958 4784
rect 5760 4586 5816 4642
rect 5902 4586 5958 4642
rect 5760 4444 5816 4500
rect 5902 4444 5958 4500
rect 5760 4302 5816 4358
rect 5902 4302 5958 4358
rect 5760 4160 5816 4216
rect 5902 4160 5958 4216
rect 5760 4018 5816 4074
rect 5902 4018 5958 4074
rect 5760 3876 5816 3932
rect 5902 3876 5958 3932
rect 5760 3734 5816 3790
rect 5902 3734 5958 3790
rect 5760 3592 5816 3648
rect 5902 3592 5958 3648
rect 5760 3450 5816 3506
rect 5902 3450 5958 3506
rect 5760 3308 5816 3364
rect 5902 3308 5958 3364
rect 5760 3166 5816 3222
rect 5902 3166 5958 3222
rect 5760 3024 5816 3080
rect 5902 3024 5958 3080
rect 5760 2882 5816 2938
rect 5902 2882 5958 2938
rect 5760 2740 5816 2796
rect 5902 2740 5958 2796
rect 5760 2598 5816 2654
rect 5902 2598 5958 2654
rect 5760 2456 5816 2512
rect 5902 2456 5958 2512
rect 5760 2314 5816 2370
rect 5902 2314 5958 2370
rect 5760 2172 5816 2228
rect 5902 2172 5958 2228
rect 5760 2030 5816 2086
rect 5902 2030 5958 2086
rect 5760 1888 5816 1944
rect 5902 1888 5958 1944
rect 5760 1746 5816 1802
rect 5902 1746 5958 1802
rect 5760 1604 5816 1660
rect 5902 1604 5958 1660
rect 5760 1462 5816 1518
rect 5902 1462 5958 1518
rect 5760 1320 5816 1376
rect 5902 1320 5958 1376
rect 5760 1178 5816 1234
rect 5902 1178 5958 1234
rect 5760 1036 5816 1092
rect 5902 1036 5958 1092
rect 5760 894 5816 950
rect 5902 894 5958 950
rect 5760 752 5816 808
rect 5902 752 5958 808
rect 5760 610 5816 666
rect 5902 610 5958 666
rect 5760 468 5816 524
rect 5902 468 5958 524
rect 6300 12254 6356 12310
rect 6442 12254 6498 12310
rect 6300 12112 6356 12168
rect 6442 12112 6498 12168
rect 6300 11970 6356 12026
rect 6442 11970 6498 12026
rect 6300 11828 6356 11884
rect 6442 11828 6498 11884
rect 6300 11686 6356 11742
rect 6442 11686 6498 11742
rect 6300 11544 6356 11600
rect 6442 11544 6498 11600
rect 6300 11402 6356 11458
rect 6442 11402 6498 11458
rect 6300 11260 6356 11316
rect 6442 11260 6498 11316
rect 6300 11118 6356 11174
rect 6442 11118 6498 11174
rect 6300 10976 6356 11032
rect 6442 10976 6498 11032
rect 6300 10834 6356 10890
rect 6442 10834 6498 10890
rect 6300 10692 6356 10748
rect 6442 10692 6498 10748
rect 6300 10550 6356 10606
rect 6442 10550 6498 10606
rect 6300 10408 6356 10464
rect 6442 10408 6498 10464
rect 6300 10266 6356 10322
rect 6442 10266 6498 10322
rect 6300 10124 6356 10180
rect 6442 10124 6498 10180
rect 6300 9982 6356 10038
rect 6442 9982 6498 10038
rect 6300 9840 6356 9896
rect 6442 9840 6498 9896
rect 6300 9698 6356 9754
rect 6442 9698 6498 9754
rect 6300 9556 6356 9612
rect 6442 9556 6498 9612
rect 6300 9414 6356 9470
rect 6442 9414 6498 9470
rect 6300 9272 6356 9328
rect 6442 9272 6498 9328
rect 6300 9130 6356 9186
rect 6442 9130 6498 9186
rect 6300 8988 6356 9044
rect 6442 8988 6498 9044
rect 6300 8846 6356 8902
rect 6442 8846 6498 8902
rect 6300 8704 6356 8760
rect 6442 8704 6498 8760
rect 6300 8562 6356 8618
rect 6442 8562 6498 8618
rect 6300 8420 6356 8476
rect 6442 8420 6498 8476
rect 6300 8278 6356 8334
rect 6442 8278 6498 8334
rect 6300 8136 6356 8192
rect 6442 8136 6498 8192
rect 6300 7994 6356 8050
rect 6442 7994 6498 8050
rect 6300 7852 6356 7908
rect 6442 7852 6498 7908
rect 6300 7710 6356 7766
rect 6442 7710 6498 7766
rect 6300 7568 6356 7624
rect 6442 7568 6498 7624
rect 6300 7426 6356 7482
rect 6442 7426 6498 7482
rect 6300 7284 6356 7340
rect 6442 7284 6498 7340
rect 6300 7142 6356 7198
rect 6442 7142 6498 7198
rect 6300 7000 6356 7056
rect 6442 7000 6498 7056
rect 6300 6858 6356 6914
rect 6442 6858 6498 6914
rect 6300 6716 6356 6772
rect 6442 6716 6498 6772
rect 6300 6574 6356 6630
rect 6442 6574 6498 6630
rect 6300 6432 6356 6488
rect 6442 6432 6498 6488
rect 6300 6290 6356 6346
rect 6442 6290 6498 6346
rect 6300 6148 6356 6204
rect 6442 6148 6498 6204
rect 6300 6006 6356 6062
rect 6442 6006 6498 6062
rect 6300 5864 6356 5920
rect 6442 5864 6498 5920
rect 6300 5722 6356 5778
rect 6442 5722 6498 5778
rect 6300 5580 6356 5636
rect 6442 5580 6498 5636
rect 6300 5438 6356 5494
rect 6442 5438 6498 5494
rect 6300 5296 6356 5352
rect 6442 5296 6498 5352
rect 6300 5154 6356 5210
rect 6442 5154 6498 5210
rect 6300 5012 6356 5068
rect 6442 5012 6498 5068
rect 6300 4870 6356 4926
rect 6442 4870 6498 4926
rect 6300 4728 6356 4784
rect 6442 4728 6498 4784
rect 6300 4586 6356 4642
rect 6442 4586 6498 4642
rect 6300 4444 6356 4500
rect 6442 4444 6498 4500
rect 6300 4302 6356 4358
rect 6442 4302 6498 4358
rect 6300 4160 6356 4216
rect 6442 4160 6498 4216
rect 6300 4018 6356 4074
rect 6442 4018 6498 4074
rect 6300 3876 6356 3932
rect 6442 3876 6498 3932
rect 6300 3734 6356 3790
rect 6442 3734 6498 3790
rect 6300 3592 6356 3648
rect 6442 3592 6498 3648
rect 6300 3450 6356 3506
rect 6442 3450 6498 3506
rect 6300 3308 6356 3364
rect 6442 3308 6498 3364
rect 6300 3166 6356 3222
rect 6442 3166 6498 3222
rect 6300 3024 6356 3080
rect 6442 3024 6498 3080
rect 6300 2882 6356 2938
rect 6442 2882 6498 2938
rect 6300 2740 6356 2796
rect 6442 2740 6498 2796
rect 6300 2598 6356 2654
rect 6442 2598 6498 2654
rect 6300 2456 6356 2512
rect 6442 2456 6498 2512
rect 6300 2314 6356 2370
rect 6442 2314 6498 2370
rect 6300 2172 6356 2228
rect 6442 2172 6498 2228
rect 6300 2030 6356 2086
rect 6442 2030 6498 2086
rect 6300 1888 6356 1944
rect 6442 1888 6498 1944
rect 6300 1746 6356 1802
rect 6442 1746 6498 1802
rect 6300 1604 6356 1660
rect 6442 1604 6498 1660
rect 6300 1462 6356 1518
rect 6442 1462 6498 1518
rect 6300 1320 6356 1376
rect 6442 1320 6498 1376
rect 6300 1178 6356 1234
rect 6442 1178 6498 1234
rect 6300 1036 6356 1092
rect 6442 1036 6498 1092
rect 6300 894 6356 950
rect 6442 894 6498 950
rect 6300 752 6356 808
rect 6442 752 6498 808
rect 6300 610 6356 666
rect 6442 610 6498 666
rect 6300 468 6356 524
rect 6442 468 6498 524
rect 6845 12254 6901 12310
rect 6987 12254 7043 12310
rect 6845 12112 6901 12168
rect 6987 12112 7043 12168
rect 6845 11970 6901 12026
rect 6987 11970 7043 12026
rect 6845 11828 6901 11884
rect 6987 11828 7043 11884
rect 6845 11686 6901 11742
rect 6987 11686 7043 11742
rect 6845 11544 6901 11600
rect 6987 11544 7043 11600
rect 6845 11402 6901 11458
rect 6987 11402 7043 11458
rect 6845 11260 6901 11316
rect 6987 11260 7043 11316
rect 6845 11118 6901 11174
rect 6987 11118 7043 11174
rect 6845 10976 6901 11032
rect 6987 10976 7043 11032
rect 6845 10834 6901 10890
rect 6987 10834 7043 10890
rect 6845 10692 6901 10748
rect 6987 10692 7043 10748
rect 6845 10550 6901 10606
rect 6987 10550 7043 10606
rect 6845 10408 6901 10464
rect 6987 10408 7043 10464
rect 6845 10266 6901 10322
rect 6987 10266 7043 10322
rect 6845 10124 6901 10180
rect 6987 10124 7043 10180
rect 6845 9982 6901 10038
rect 6987 9982 7043 10038
rect 6845 9840 6901 9896
rect 6987 9840 7043 9896
rect 6845 9698 6901 9754
rect 6987 9698 7043 9754
rect 6845 9556 6901 9612
rect 6987 9556 7043 9612
rect 6845 9414 6901 9470
rect 6987 9414 7043 9470
rect 6845 9272 6901 9328
rect 6987 9272 7043 9328
rect 6845 9130 6901 9186
rect 6987 9130 7043 9186
rect 6845 8988 6901 9044
rect 6987 8988 7043 9044
rect 6845 8846 6901 8902
rect 6987 8846 7043 8902
rect 6845 8704 6901 8760
rect 6987 8704 7043 8760
rect 6845 8562 6901 8618
rect 6987 8562 7043 8618
rect 6845 8420 6901 8476
rect 6987 8420 7043 8476
rect 6845 8278 6901 8334
rect 6987 8278 7043 8334
rect 6845 8136 6901 8192
rect 6987 8136 7043 8192
rect 6845 7994 6901 8050
rect 6987 7994 7043 8050
rect 6845 7852 6901 7908
rect 6987 7852 7043 7908
rect 6845 7710 6901 7766
rect 6987 7710 7043 7766
rect 6845 7568 6901 7624
rect 6987 7568 7043 7624
rect 6845 7426 6901 7482
rect 6987 7426 7043 7482
rect 6845 7284 6901 7340
rect 6987 7284 7043 7340
rect 6845 7142 6901 7198
rect 6987 7142 7043 7198
rect 6845 7000 6901 7056
rect 6987 7000 7043 7056
rect 6845 6858 6901 6914
rect 6987 6858 7043 6914
rect 6845 6716 6901 6772
rect 6987 6716 7043 6772
rect 6845 6574 6901 6630
rect 6987 6574 7043 6630
rect 6845 6432 6901 6488
rect 6987 6432 7043 6488
rect 6845 6290 6901 6346
rect 6987 6290 7043 6346
rect 6845 6148 6901 6204
rect 6987 6148 7043 6204
rect 6845 6006 6901 6062
rect 6987 6006 7043 6062
rect 6845 5864 6901 5920
rect 6987 5864 7043 5920
rect 6845 5722 6901 5778
rect 6987 5722 7043 5778
rect 6845 5580 6901 5636
rect 6987 5580 7043 5636
rect 6845 5438 6901 5494
rect 6987 5438 7043 5494
rect 6845 5296 6901 5352
rect 6987 5296 7043 5352
rect 6845 5154 6901 5210
rect 6987 5154 7043 5210
rect 6845 5012 6901 5068
rect 6987 5012 7043 5068
rect 6845 4870 6901 4926
rect 6987 4870 7043 4926
rect 6845 4728 6901 4784
rect 6987 4728 7043 4784
rect 6845 4586 6901 4642
rect 6987 4586 7043 4642
rect 6845 4444 6901 4500
rect 6987 4444 7043 4500
rect 6845 4302 6901 4358
rect 6987 4302 7043 4358
rect 6845 4160 6901 4216
rect 6987 4160 7043 4216
rect 6845 4018 6901 4074
rect 6987 4018 7043 4074
rect 6845 3876 6901 3932
rect 6987 3876 7043 3932
rect 6845 3734 6901 3790
rect 6987 3734 7043 3790
rect 6845 3592 6901 3648
rect 6987 3592 7043 3648
rect 6845 3450 6901 3506
rect 6987 3450 7043 3506
rect 6845 3308 6901 3364
rect 6987 3308 7043 3364
rect 6845 3166 6901 3222
rect 6987 3166 7043 3222
rect 6845 3024 6901 3080
rect 6987 3024 7043 3080
rect 6845 2882 6901 2938
rect 6987 2882 7043 2938
rect 6845 2740 6901 2796
rect 6987 2740 7043 2796
rect 6845 2598 6901 2654
rect 6987 2598 7043 2654
rect 6845 2456 6901 2512
rect 6987 2456 7043 2512
rect 6845 2314 6901 2370
rect 6987 2314 7043 2370
rect 6845 2172 6901 2228
rect 6987 2172 7043 2228
rect 6845 2030 6901 2086
rect 6987 2030 7043 2086
rect 6845 1888 6901 1944
rect 6987 1888 7043 1944
rect 6845 1746 6901 1802
rect 6987 1746 7043 1802
rect 6845 1604 6901 1660
rect 6987 1604 7043 1660
rect 6845 1462 6901 1518
rect 6987 1462 7043 1518
rect 6845 1320 6901 1376
rect 6987 1320 7043 1376
rect 6845 1178 6901 1234
rect 6987 1178 7043 1234
rect 6845 1036 6901 1092
rect 6987 1036 7043 1092
rect 6845 894 6901 950
rect 6987 894 7043 950
rect 6845 752 6901 808
rect 6987 752 7043 808
rect 6845 610 6901 666
rect 6987 610 7043 666
rect 6845 468 6901 524
rect 6987 468 7043 524
rect 7382 12254 7438 12310
rect 7524 12254 7580 12310
rect 7382 12112 7438 12168
rect 7524 12112 7580 12168
rect 7382 11970 7438 12026
rect 7524 11970 7580 12026
rect 7382 11828 7438 11884
rect 7524 11828 7580 11884
rect 7382 11686 7438 11742
rect 7524 11686 7580 11742
rect 7382 11544 7438 11600
rect 7524 11544 7580 11600
rect 7382 11402 7438 11458
rect 7524 11402 7580 11458
rect 7382 11260 7438 11316
rect 7524 11260 7580 11316
rect 7382 11118 7438 11174
rect 7524 11118 7580 11174
rect 7382 10976 7438 11032
rect 7524 10976 7580 11032
rect 7382 10834 7438 10890
rect 7524 10834 7580 10890
rect 7382 10692 7438 10748
rect 7524 10692 7580 10748
rect 7382 10550 7438 10606
rect 7524 10550 7580 10606
rect 7382 10408 7438 10464
rect 7524 10408 7580 10464
rect 7382 10266 7438 10322
rect 7524 10266 7580 10322
rect 7382 10124 7438 10180
rect 7524 10124 7580 10180
rect 7382 9982 7438 10038
rect 7524 9982 7580 10038
rect 7382 9840 7438 9896
rect 7524 9840 7580 9896
rect 7382 9698 7438 9754
rect 7524 9698 7580 9754
rect 7382 9556 7438 9612
rect 7524 9556 7580 9612
rect 7382 9414 7438 9470
rect 7524 9414 7580 9470
rect 7382 9272 7438 9328
rect 7524 9272 7580 9328
rect 7382 9130 7438 9186
rect 7524 9130 7580 9186
rect 7382 8988 7438 9044
rect 7524 8988 7580 9044
rect 7382 8846 7438 8902
rect 7524 8846 7580 8902
rect 7382 8704 7438 8760
rect 7524 8704 7580 8760
rect 7382 8562 7438 8618
rect 7524 8562 7580 8618
rect 7382 8420 7438 8476
rect 7524 8420 7580 8476
rect 7382 8278 7438 8334
rect 7524 8278 7580 8334
rect 7382 8136 7438 8192
rect 7524 8136 7580 8192
rect 7382 7994 7438 8050
rect 7524 7994 7580 8050
rect 7382 7852 7438 7908
rect 7524 7852 7580 7908
rect 7382 7710 7438 7766
rect 7524 7710 7580 7766
rect 7382 7568 7438 7624
rect 7524 7568 7580 7624
rect 7382 7426 7438 7482
rect 7524 7426 7580 7482
rect 7382 7284 7438 7340
rect 7524 7284 7580 7340
rect 7382 7142 7438 7198
rect 7524 7142 7580 7198
rect 7382 7000 7438 7056
rect 7524 7000 7580 7056
rect 7382 6858 7438 6914
rect 7524 6858 7580 6914
rect 7382 6716 7438 6772
rect 7524 6716 7580 6772
rect 7382 6574 7438 6630
rect 7524 6574 7580 6630
rect 7382 6432 7438 6488
rect 7524 6432 7580 6488
rect 7382 6290 7438 6346
rect 7524 6290 7580 6346
rect 7382 6148 7438 6204
rect 7524 6148 7580 6204
rect 7382 6006 7438 6062
rect 7524 6006 7580 6062
rect 7382 5864 7438 5920
rect 7524 5864 7580 5920
rect 7382 5722 7438 5778
rect 7524 5722 7580 5778
rect 7382 5580 7438 5636
rect 7524 5580 7580 5636
rect 7382 5438 7438 5494
rect 7524 5438 7580 5494
rect 7382 5296 7438 5352
rect 7524 5296 7580 5352
rect 7382 5154 7438 5210
rect 7524 5154 7580 5210
rect 7382 5012 7438 5068
rect 7524 5012 7580 5068
rect 7382 4870 7438 4926
rect 7524 4870 7580 4926
rect 7382 4728 7438 4784
rect 7524 4728 7580 4784
rect 7382 4586 7438 4642
rect 7524 4586 7580 4642
rect 7382 4444 7438 4500
rect 7524 4444 7580 4500
rect 7382 4302 7438 4358
rect 7524 4302 7580 4358
rect 7382 4160 7438 4216
rect 7524 4160 7580 4216
rect 7382 4018 7438 4074
rect 7524 4018 7580 4074
rect 7382 3876 7438 3932
rect 7524 3876 7580 3932
rect 7382 3734 7438 3790
rect 7524 3734 7580 3790
rect 7382 3592 7438 3648
rect 7524 3592 7580 3648
rect 7382 3450 7438 3506
rect 7524 3450 7580 3506
rect 7382 3308 7438 3364
rect 7524 3308 7580 3364
rect 7382 3166 7438 3222
rect 7524 3166 7580 3222
rect 7382 3024 7438 3080
rect 7524 3024 7580 3080
rect 7382 2882 7438 2938
rect 7524 2882 7580 2938
rect 7382 2740 7438 2796
rect 7524 2740 7580 2796
rect 7382 2598 7438 2654
rect 7524 2598 7580 2654
rect 7382 2456 7438 2512
rect 7524 2456 7580 2512
rect 7382 2314 7438 2370
rect 7524 2314 7580 2370
rect 7382 2172 7438 2228
rect 7524 2172 7580 2228
rect 7382 2030 7438 2086
rect 7524 2030 7580 2086
rect 7382 1888 7438 1944
rect 7524 1888 7580 1944
rect 7382 1746 7438 1802
rect 7524 1746 7580 1802
rect 7382 1604 7438 1660
rect 7524 1604 7580 1660
rect 7382 1462 7438 1518
rect 7524 1462 7580 1518
rect 7382 1320 7438 1376
rect 7524 1320 7580 1376
rect 7382 1178 7438 1234
rect 7524 1178 7580 1234
rect 7382 1036 7438 1092
rect 7524 1036 7580 1092
rect 7382 894 7438 950
rect 7524 894 7580 950
rect 7382 752 7438 808
rect 7524 752 7580 808
rect 7382 610 7438 666
rect 7524 610 7580 666
rect 7382 468 7438 524
rect 7524 468 7580 524
rect 7919 12254 7975 12310
rect 8061 12254 8117 12310
rect 7919 12112 7975 12168
rect 8061 12112 8117 12168
rect 7919 11970 7975 12026
rect 8061 11970 8117 12026
rect 7919 11828 7975 11884
rect 8061 11828 8117 11884
rect 7919 11686 7975 11742
rect 8061 11686 8117 11742
rect 7919 11544 7975 11600
rect 8061 11544 8117 11600
rect 7919 11402 7975 11458
rect 8061 11402 8117 11458
rect 7919 11260 7975 11316
rect 8061 11260 8117 11316
rect 7919 11118 7975 11174
rect 8061 11118 8117 11174
rect 7919 10976 7975 11032
rect 8061 10976 8117 11032
rect 7919 10834 7975 10890
rect 8061 10834 8117 10890
rect 7919 10692 7975 10748
rect 8061 10692 8117 10748
rect 7919 10550 7975 10606
rect 8061 10550 8117 10606
rect 7919 10408 7975 10464
rect 8061 10408 8117 10464
rect 7919 10266 7975 10322
rect 8061 10266 8117 10322
rect 7919 10124 7975 10180
rect 8061 10124 8117 10180
rect 7919 9982 7975 10038
rect 8061 9982 8117 10038
rect 7919 9840 7975 9896
rect 8061 9840 8117 9896
rect 7919 9698 7975 9754
rect 8061 9698 8117 9754
rect 7919 9556 7975 9612
rect 8061 9556 8117 9612
rect 7919 9414 7975 9470
rect 8061 9414 8117 9470
rect 7919 9272 7975 9328
rect 8061 9272 8117 9328
rect 7919 9130 7975 9186
rect 8061 9130 8117 9186
rect 7919 8988 7975 9044
rect 8061 8988 8117 9044
rect 7919 8846 7975 8902
rect 8061 8846 8117 8902
rect 7919 8704 7975 8760
rect 8061 8704 8117 8760
rect 7919 8562 7975 8618
rect 8061 8562 8117 8618
rect 7919 8420 7975 8476
rect 8061 8420 8117 8476
rect 7919 8278 7975 8334
rect 8061 8278 8117 8334
rect 7919 8136 7975 8192
rect 8061 8136 8117 8192
rect 7919 7994 7975 8050
rect 8061 7994 8117 8050
rect 7919 7852 7975 7908
rect 8061 7852 8117 7908
rect 7919 7710 7975 7766
rect 8061 7710 8117 7766
rect 7919 7568 7975 7624
rect 8061 7568 8117 7624
rect 7919 7426 7975 7482
rect 8061 7426 8117 7482
rect 7919 7284 7975 7340
rect 8061 7284 8117 7340
rect 7919 7142 7975 7198
rect 8061 7142 8117 7198
rect 7919 7000 7975 7056
rect 8061 7000 8117 7056
rect 7919 6858 7975 6914
rect 8061 6858 8117 6914
rect 7919 6716 7975 6772
rect 8061 6716 8117 6772
rect 7919 6574 7975 6630
rect 8061 6574 8117 6630
rect 7919 6432 7975 6488
rect 8061 6432 8117 6488
rect 7919 6290 7975 6346
rect 8061 6290 8117 6346
rect 7919 6148 7975 6204
rect 8061 6148 8117 6204
rect 7919 6006 7975 6062
rect 8061 6006 8117 6062
rect 7919 5864 7975 5920
rect 8061 5864 8117 5920
rect 7919 5722 7975 5778
rect 8061 5722 8117 5778
rect 7919 5580 7975 5636
rect 8061 5580 8117 5636
rect 7919 5438 7975 5494
rect 8061 5438 8117 5494
rect 7919 5296 7975 5352
rect 8061 5296 8117 5352
rect 7919 5154 7975 5210
rect 8061 5154 8117 5210
rect 7919 5012 7975 5068
rect 8061 5012 8117 5068
rect 7919 4870 7975 4926
rect 8061 4870 8117 4926
rect 7919 4728 7975 4784
rect 8061 4728 8117 4784
rect 7919 4586 7975 4642
rect 8061 4586 8117 4642
rect 7919 4444 7975 4500
rect 8061 4444 8117 4500
rect 7919 4302 7975 4358
rect 8061 4302 8117 4358
rect 7919 4160 7975 4216
rect 8061 4160 8117 4216
rect 7919 4018 7975 4074
rect 8061 4018 8117 4074
rect 7919 3876 7975 3932
rect 8061 3876 8117 3932
rect 7919 3734 7975 3790
rect 8061 3734 8117 3790
rect 7919 3592 7975 3648
rect 8061 3592 8117 3648
rect 7919 3450 7975 3506
rect 8061 3450 8117 3506
rect 7919 3308 7975 3364
rect 8061 3308 8117 3364
rect 7919 3166 7975 3222
rect 8061 3166 8117 3222
rect 7919 3024 7975 3080
rect 8061 3024 8117 3080
rect 7919 2882 7975 2938
rect 8061 2882 8117 2938
rect 7919 2740 7975 2796
rect 8061 2740 8117 2796
rect 7919 2598 7975 2654
rect 8061 2598 8117 2654
rect 7919 2456 7975 2512
rect 8061 2456 8117 2512
rect 7919 2314 7975 2370
rect 8061 2314 8117 2370
rect 7919 2172 7975 2228
rect 8061 2172 8117 2228
rect 7919 2030 7975 2086
rect 8061 2030 8117 2086
rect 7919 1888 7975 1944
rect 8061 1888 8117 1944
rect 7919 1746 7975 1802
rect 8061 1746 8117 1802
rect 7919 1604 7975 1660
rect 8061 1604 8117 1660
rect 7919 1462 7975 1518
rect 8061 1462 8117 1518
rect 7919 1320 7975 1376
rect 8061 1320 8117 1376
rect 7919 1178 7975 1234
rect 8061 1178 8117 1234
rect 7919 1036 7975 1092
rect 8061 1036 8117 1092
rect 7919 894 7975 950
rect 8061 894 8117 950
rect 7919 752 7975 808
rect 8061 752 8117 808
rect 7919 610 7975 666
rect 8061 610 8117 666
rect 7919 468 7975 524
rect 8061 468 8117 524
rect 8462 12254 8518 12310
rect 8604 12254 8660 12310
rect 8462 12112 8518 12168
rect 8604 12112 8660 12168
rect 8462 11970 8518 12026
rect 8604 11970 8660 12026
rect 8462 11828 8518 11884
rect 8604 11828 8660 11884
rect 8462 11686 8518 11742
rect 8604 11686 8660 11742
rect 8462 11544 8518 11600
rect 8604 11544 8660 11600
rect 8462 11402 8518 11458
rect 8604 11402 8660 11458
rect 8462 11260 8518 11316
rect 8604 11260 8660 11316
rect 8462 11118 8518 11174
rect 8604 11118 8660 11174
rect 8462 10976 8518 11032
rect 8604 10976 8660 11032
rect 8462 10834 8518 10890
rect 8604 10834 8660 10890
rect 8462 10692 8518 10748
rect 8604 10692 8660 10748
rect 8462 10550 8518 10606
rect 8604 10550 8660 10606
rect 8462 10408 8518 10464
rect 8604 10408 8660 10464
rect 8462 10266 8518 10322
rect 8604 10266 8660 10322
rect 8462 10124 8518 10180
rect 8604 10124 8660 10180
rect 8462 9982 8518 10038
rect 8604 9982 8660 10038
rect 8462 9840 8518 9896
rect 8604 9840 8660 9896
rect 8462 9698 8518 9754
rect 8604 9698 8660 9754
rect 8462 9556 8518 9612
rect 8604 9556 8660 9612
rect 8462 9414 8518 9470
rect 8604 9414 8660 9470
rect 8462 9272 8518 9328
rect 8604 9272 8660 9328
rect 8462 9130 8518 9186
rect 8604 9130 8660 9186
rect 8462 8988 8518 9044
rect 8604 8988 8660 9044
rect 8462 8846 8518 8902
rect 8604 8846 8660 8902
rect 8462 8704 8518 8760
rect 8604 8704 8660 8760
rect 8462 8562 8518 8618
rect 8604 8562 8660 8618
rect 8462 8420 8518 8476
rect 8604 8420 8660 8476
rect 8462 8278 8518 8334
rect 8604 8278 8660 8334
rect 8462 8136 8518 8192
rect 8604 8136 8660 8192
rect 8462 7994 8518 8050
rect 8604 7994 8660 8050
rect 8462 7852 8518 7908
rect 8604 7852 8660 7908
rect 8462 7710 8518 7766
rect 8604 7710 8660 7766
rect 8462 7568 8518 7624
rect 8604 7568 8660 7624
rect 8462 7426 8518 7482
rect 8604 7426 8660 7482
rect 8462 7284 8518 7340
rect 8604 7284 8660 7340
rect 8462 7142 8518 7198
rect 8604 7142 8660 7198
rect 8462 7000 8518 7056
rect 8604 7000 8660 7056
rect 8462 6858 8518 6914
rect 8604 6858 8660 6914
rect 8462 6716 8518 6772
rect 8604 6716 8660 6772
rect 8462 6574 8518 6630
rect 8604 6574 8660 6630
rect 8462 6432 8518 6488
rect 8604 6432 8660 6488
rect 8462 6290 8518 6346
rect 8604 6290 8660 6346
rect 8462 6148 8518 6204
rect 8604 6148 8660 6204
rect 8462 6006 8518 6062
rect 8604 6006 8660 6062
rect 8462 5864 8518 5920
rect 8604 5864 8660 5920
rect 8462 5722 8518 5778
rect 8604 5722 8660 5778
rect 8462 5580 8518 5636
rect 8604 5580 8660 5636
rect 8462 5438 8518 5494
rect 8604 5438 8660 5494
rect 8462 5296 8518 5352
rect 8604 5296 8660 5352
rect 8462 5154 8518 5210
rect 8604 5154 8660 5210
rect 8462 5012 8518 5068
rect 8604 5012 8660 5068
rect 8462 4870 8518 4926
rect 8604 4870 8660 4926
rect 8462 4728 8518 4784
rect 8604 4728 8660 4784
rect 8462 4586 8518 4642
rect 8604 4586 8660 4642
rect 8462 4444 8518 4500
rect 8604 4444 8660 4500
rect 8462 4302 8518 4358
rect 8604 4302 8660 4358
rect 8462 4160 8518 4216
rect 8604 4160 8660 4216
rect 8462 4018 8518 4074
rect 8604 4018 8660 4074
rect 8462 3876 8518 3932
rect 8604 3876 8660 3932
rect 8462 3734 8518 3790
rect 8604 3734 8660 3790
rect 8462 3592 8518 3648
rect 8604 3592 8660 3648
rect 8462 3450 8518 3506
rect 8604 3450 8660 3506
rect 8462 3308 8518 3364
rect 8604 3308 8660 3364
rect 8462 3166 8518 3222
rect 8604 3166 8660 3222
rect 8462 3024 8518 3080
rect 8604 3024 8660 3080
rect 8462 2882 8518 2938
rect 8604 2882 8660 2938
rect 8462 2740 8518 2796
rect 8604 2740 8660 2796
rect 8462 2598 8518 2654
rect 8604 2598 8660 2654
rect 8462 2456 8518 2512
rect 8604 2456 8660 2512
rect 8462 2314 8518 2370
rect 8604 2314 8660 2370
rect 8462 2172 8518 2228
rect 8604 2172 8660 2228
rect 8462 2030 8518 2086
rect 8604 2030 8660 2086
rect 8462 1888 8518 1944
rect 8604 1888 8660 1944
rect 8462 1746 8518 1802
rect 8604 1746 8660 1802
rect 8462 1604 8518 1660
rect 8604 1604 8660 1660
rect 8462 1462 8518 1518
rect 8604 1462 8660 1518
rect 8462 1320 8518 1376
rect 8604 1320 8660 1376
rect 8462 1178 8518 1234
rect 8604 1178 8660 1234
rect 8462 1036 8518 1092
rect 8604 1036 8660 1092
rect 8462 894 8518 950
rect 8604 894 8660 950
rect 8462 752 8518 808
rect 8604 752 8660 808
rect 8462 610 8518 666
rect 8604 610 8660 666
rect 8462 468 8518 524
rect 8604 468 8660 524
rect 9004 12254 9060 12310
rect 9146 12254 9202 12310
rect 9004 12112 9060 12168
rect 9146 12112 9202 12168
rect 9004 11970 9060 12026
rect 9146 11970 9202 12026
rect 9004 11828 9060 11884
rect 9146 11828 9202 11884
rect 9004 11686 9060 11742
rect 9146 11686 9202 11742
rect 9004 11544 9060 11600
rect 9146 11544 9202 11600
rect 9004 11402 9060 11458
rect 9146 11402 9202 11458
rect 9004 11260 9060 11316
rect 9146 11260 9202 11316
rect 9004 11118 9060 11174
rect 9146 11118 9202 11174
rect 9004 10976 9060 11032
rect 9146 10976 9202 11032
rect 9004 10834 9060 10890
rect 9146 10834 9202 10890
rect 9004 10692 9060 10748
rect 9146 10692 9202 10748
rect 9004 10550 9060 10606
rect 9146 10550 9202 10606
rect 9004 10408 9060 10464
rect 9146 10408 9202 10464
rect 9004 10266 9060 10322
rect 9146 10266 9202 10322
rect 9004 10124 9060 10180
rect 9146 10124 9202 10180
rect 9004 9982 9060 10038
rect 9146 9982 9202 10038
rect 9004 9840 9060 9896
rect 9146 9840 9202 9896
rect 9004 9698 9060 9754
rect 9146 9698 9202 9754
rect 9004 9556 9060 9612
rect 9146 9556 9202 9612
rect 9004 9414 9060 9470
rect 9146 9414 9202 9470
rect 9004 9272 9060 9328
rect 9146 9272 9202 9328
rect 9004 9130 9060 9186
rect 9146 9130 9202 9186
rect 9004 8988 9060 9044
rect 9146 8988 9202 9044
rect 9004 8846 9060 8902
rect 9146 8846 9202 8902
rect 9004 8704 9060 8760
rect 9146 8704 9202 8760
rect 9004 8562 9060 8618
rect 9146 8562 9202 8618
rect 9004 8420 9060 8476
rect 9146 8420 9202 8476
rect 9004 8278 9060 8334
rect 9146 8278 9202 8334
rect 9004 8136 9060 8192
rect 9146 8136 9202 8192
rect 9004 7994 9060 8050
rect 9146 7994 9202 8050
rect 9004 7852 9060 7908
rect 9146 7852 9202 7908
rect 9004 7710 9060 7766
rect 9146 7710 9202 7766
rect 9004 7568 9060 7624
rect 9146 7568 9202 7624
rect 9004 7426 9060 7482
rect 9146 7426 9202 7482
rect 9004 7284 9060 7340
rect 9146 7284 9202 7340
rect 9004 7142 9060 7198
rect 9146 7142 9202 7198
rect 9004 7000 9060 7056
rect 9146 7000 9202 7056
rect 9004 6858 9060 6914
rect 9146 6858 9202 6914
rect 9004 6716 9060 6772
rect 9146 6716 9202 6772
rect 9004 6574 9060 6630
rect 9146 6574 9202 6630
rect 9004 6432 9060 6488
rect 9146 6432 9202 6488
rect 9004 6290 9060 6346
rect 9146 6290 9202 6346
rect 9004 6148 9060 6204
rect 9146 6148 9202 6204
rect 9004 6006 9060 6062
rect 9146 6006 9202 6062
rect 9004 5864 9060 5920
rect 9146 5864 9202 5920
rect 9004 5722 9060 5778
rect 9146 5722 9202 5778
rect 9004 5580 9060 5636
rect 9146 5580 9202 5636
rect 9004 5438 9060 5494
rect 9146 5438 9202 5494
rect 9004 5296 9060 5352
rect 9146 5296 9202 5352
rect 9004 5154 9060 5210
rect 9146 5154 9202 5210
rect 9004 5012 9060 5068
rect 9146 5012 9202 5068
rect 9004 4870 9060 4926
rect 9146 4870 9202 4926
rect 9004 4728 9060 4784
rect 9146 4728 9202 4784
rect 9004 4586 9060 4642
rect 9146 4586 9202 4642
rect 9004 4444 9060 4500
rect 9146 4444 9202 4500
rect 9004 4302 9060 4358
rect 9146 4302 9202 4358
rect 9004 4160 9060 4216
rect 9146 4160 9202 4216
rect 9004 4018 9060 4074
rect 9146 4018 9202 4074
rect 9004 3876 9060 3932
rect 9146 3876 9202 3932
rect 9004 3734 9060 3790
rect 9146 3734 9202 3790
rect 9004 3592 9060 3648
rect 9146 3592 9202 3648
rect 9004 3450 9060 3506
rect 9146 3450 9202 3506
rect 9004 3308 9060 3364
rect 9146 3308 9202 3364
rect 9004 3166 9060 3222
rect 9146 3166 9202 3222
rect 9004 3024 9060 3080
rect 9146 3024 9202 3080
rect 9004 2882 9060 2938
rect 9146 2882 9202 2938
rect 9004 2740 9060 2796
rect 9146 2740 9202 2796
rect 9004 2598 9060 2654
rect 9146 2598 9202 2654
rect 9004 2456 9060 2512
rect 9146 2456 9202 2512
rect 9004 2314 9060 2370
rect 9146 2314 9202 2370
rect 9004 2172 9060 2228
rect 9146 2172 9202 2228
rect 9004 2030 9060 2086
rect 9146 2030 9202 2086
rect 9004 1888 9060 1944
rect 9146 1888 9202 1944
rect 9004 1746 9060 1802
rect 9146 1746 9202 1802
rect 9004 1604 9060 1660
rect 9146 1604 9202 1660
rect 9004 1462 9060 1518
rect 9146 1462 9202 1518
rect 9004 1320 9060 1376
rect 9146 1320 9202 1376
rect 9004 1178 9060 1234
rect 9146 1178 9202 1234
rect 9004 1036 9060 1092
rect 9146 1036 9202 1092
rect 9004 894 9060 950
rect 9146 894 9202 950
rect 9004 752 9060 808
rect 9146 752 9202 808
rect 9004 610 9060 666
rect 9146 610 9202 666
rect 9004 468 9060 524
rect 9146 468 9202 524
rect 9547 12254 9603 12310
rect 9689 12254 9745 12310
rect 9547 12112 9603 12168
rect 9689 12112 9745 12168
rect 9547 11970 9603 12026
rect 9689 11970 9745 12026
rect 9547 11828 9603 11884
rect 9689 11828 9745 11884
rect 9547 11686 9603 11742
rect 9689 11686 9745 11742
rect 9547 11544 9603 11600
rect 9689 11544 9745 11600
rect 9547 11402 9603 11458
rect 9689 11402 9745 11458
rect 9547 11260 9603 11316
rect 9689 11260 9745 11316
rect 9547 11118 9603 11174
rect 9689 11118 9745 11174
rect 9547 10976 9603 11032
rect 9689 10976 9745 11032
rect 9547 10834 9603 10890
rect 9689 10834 9745 10890
rect 9547 10692 9603 10748
rect 9689 10692 9745 10748
rect 9547 10550 9603 10606
rect 9689 10550 9745 10606
rect 9547 10408 9603 10464
rect 9689 10408 9745 10464
rect 9547 10266 9603 10322
rect 9689 10266 9745 10322
rect 9547 10124 9603 10180
rect 9689 10124 9745 10180
rect 9547 9982 9603 10038
rect 9689 9982 9745 10038
rect 9547 9840 9603 9896
rect 9689 9840 9745 9896
rect 9547 9698 9603 9754
rect 9689 9698 9745 9754
rect 9547 9556 9603 9612
rect 9689 9556 9745 9612
rect 9547 9414 9603 9470
rect 9689 9414 9745 9470
rect 9547 9272 9603 9328
rect 9689 9272 9745 9328
rect 9547 9130 9603 9186
rect 9689 9130 9745 9186
rect 9547 8988 9603 9044
rect 9689 8988 9745 9044
rect 9547 8846 9603 8902
rect 9689 8846 9745 8902
rect 9547 8704 9603 8760
rect 9689 8704 9745 8760
rect 9547 8562 9603 8618
rect 9689 8562 9745 8618
rect 9547 8420 9603 8476
rect 9689 8420 9745 8476
rect 9547 8278 9603 8334
rect 9689 8278 9745 8334
rect 9547 8136 9603 8192
rect 9689 8136 9745 8192
rect 9547 7994 9603 8050
rect 9689 7994 9745 8050
rect 9547 7852 9603 7908
rect 9689 7852 9745 7908
rect 9547 7710 9603 7766
rect 9689 7710 9745 7766
rect 9547 7568 9603 7624
rect 9689 7568 9745 7624
rect 9547 7426 9603 7482
rect 9689 7426 9745 7482
rect 9547 7284 9603 7340
rect 9689 7284 9745 7340
rect 9547 7142 9603 7198
rect 9689 7142 9745 7198
rect 9547 7000 9603 7056
rect 9689 7000 9745 7056
rect 9547 6858 9603 6914
rect 9689 6858 9745 6914
rect 9547 6716 9603 6772
rect 9689 6716 9745 6772
rect 9547 6574 9603 6630
rect 9689 6574 9745 6630
rect 9547 6432 9603 6488
rect 9689 6432 9745 6488
rect 9547 6290 9603 6346
rect 9689 6290 9745 6346
rect 9547 6148 9603 6204
rect 9689 6148 9745 6204
rect 9547 6006 9603 6062
rect 9689 6006 9745 6062
rect 9547 5864 9603 5920
rect 9689 5864 9745 5920
rect 9547 5722 9603 5778
rect 9689 5722 9745 5778
rect 9547 5580 9603 5636
rect 9689 5580 9745 5636
rect 9547 5438 9603 5494
rect 9689 5438 9745 5494
rect 9547 5296 9603 5352
rect 9689 5296 9745 5352
rect 9547 5154 9603 5210
rect 9689 5154 9745 5210
rect 9547 5012 9603 5068
rect 9689 5012 9745 5068
rect 9547 4870 9603 4926
rect 9689 4870 9745 4926
rect 9547 4728 9603 4784
rect 9689 4728 9745 4784
rect 9547 4586 9603 4642
rect 9689 4586 9745 4642
rect 9547 4444 9603 4500
rect 9689 4444 9745 4500
rect 9547 4302 9603 4358
rect 9689 4302 9745 4358
rect 9547 4160 9603 4216
rect 9689 4160 9745 4216
rect 9547 4018 9603 4074
rect 9689 4018 9745 4074
rect 9547 3876 9603 3932
rect 9689 3876 9745 3932
rect 9547 3734 9603 3790
rect 9689 3734 9745 3790
rect 9547 3592 9603 3648
rect 9689 3592 9745 3648
rect 9547 3450 9603 3506
rect 9689 3450 9745 3506
rect 9547 3308 9603 3364
rect 9689 3308 9745 3364
rect 9547 3166 9603 3222
rect 9689 3166 9745 3222
rect 9547 3024 9603 3080
rect 9689 3024 9745 3080
rect 9547 2882 9603 2938
rect 9689 2882 9745 2938
rect 9547 2740 9603 2796
rect 9689 2740 9745 2796
rect 9547 2598 9603 2654
rect 9689 2598 9745 2654
rect 9547 2456 9603 2512
rect 9689 2456 9745 2512
rect 9547 2314 9603 2370
rect 9689 2314 9745 2370
rect 9547 2172 9603 2228
rect 9689 2172 9745 2228
rect 9547 2030 9603 2086
rect 9689 2030 9745 2086
rect 9547 1888 9603 1944
rect 9689 1888 9745 1944
rect 9547 1746 9603 1802
rect 9689 1746 9745 1802
rect 9547 1604 9603 1660
rect 9689 1604 9745 1660
rect 9547 1462 9603 1518
rect 9689 1462 9745 1518
rect 9547 1320 9603 1376
rect 9689 1320 9745 1376
rect 9547 1178 9603 1234
rect 9689 1178 9745 1234
rect 9547 1036 9603 1092
rect 9689 1036 9745 1092
rect 9547 894 9603 950
rect 9689 894 9745 950
rect 9547 752 9603 808
rect 9689 752 9745 808
rect 9547 610 9603 666
rect 9689 610 9745 666
rect 9547 468 9603 524
rect 9689 468 9745 524
rect 10081 12254 10137 12310
rect 10223 12254 10279 12310
rect 10081 12112 10137 12168
rect 10223 12112 10279 12168
rect 10081 11970 10137 12026
rect 10223 11970 10279 12026
rect 10081 11828 10137 11884
rect 10223 11828 10279 11884
rect 10081 11686 10137 11742
rect 10223 11686 10279 11742
rect 10081 11544 10137 11600
rect 10223 11544 10279 11600
rect 10081 11402 10137 11458
rect 10223 11402 10279 11458
rect 10081 11260 10137 11316
rect 10223 11260 10279 11316
rect 10081 11118 10137 11174
rect 10223 11118 10279 11174
rect 10081 10976 10137 11032
rect 10223 10976 10279 11032
rect 10081 10834 10137 10890
rect 10223 10834 10279 10890
rect 10081 10692 10137 10748
rect 10223 10692 10279 10748
rect 10081 10550 10137 10606
rect 10223 10550 10279 10606
rect 10081 10408 10137 10464
rect 10223 10408 10279 10464
rect 10081 10266 10137 10322
rect 10223 10266 10279 10322
rect 10081 10124 10137 10180
rect 10223 10124 10279 10180
rect 10081 9982 10137 10038
rect 10223 9982 10279 10038
rect 10081 9840 10137 9896
rect 10223 9840 10279 9896
rect 10081 9698 10137 9754
rect 10223 9698 10279 9754
rect 10081 9556 10137 9612
rect 10223 9556 10279 9612
rect 10081 9414 10137 9470
rect 10223 9414 10279 9470
rect 10081 9272 10137 9328
rect 10223 9272 10279 9328
rect 10081 9130 10137 9186
rect 10223 9130 10279 9186
rect 10081 8988 10137 9044
rect 10223 8988 10279 9044
rect 10081 8846 10137 8902
rect 10223 8846 10279 8902
rect 10081 8704 10137 8760
rect 10223 8704 10279 8760
rect 10081 8562 10137 8618
rect 10223 8562 10279 8618
rect 10081 8420 10137 8476
rect 10223 8420 10279 8476
rect 10081 8278 10137 8334
rect 10223 8278 10279 8334
rect 10081 8136 10137 8192
rect 10223 8136 10279 8192
rect 10081 7994 10137 8050
rect 10223 7994 10279 8050
rect 10081 7852 10137 7908
rect 10223 7852 10279 7908
rect 10081 7710 10137 7766
rect 10223 7710 10279 7766
rect 10081 7568 10137 7624
rect 10223 7568 10279 7624
rect 10081 7426 10137 7482
rect 10223 7426 10279 7482
rect 10081 7284 10137 7340
rect 10223 7284 10279 7340
rect 10081 7142 10137 7198
rect 10223 7142 10279 7198
rect 10081 7000 10137 7056
rect 10223 7000 10279 7056
rect 10081 6858 10137 6914
rect 10223 6858 10279 6914
rect 10081 6716 10137 6772
rect 10223 6716 10279 6772
rect 10081 6574 10137 6630
rect 10223 6574 10279 6630
rect 10081 6432 10137 6488
rect 10223 6432 10279 6488
rect 10081 6290 10137 6346
rect 10223 6290 10279 6346
rect 10081 6148 10137 6204
rect 10223 6148 10279 6204
rect 10081 6006 10137 6062
rect 10223 6006 10279 6062
rect 10081 5864 10137 5920
rect 10223 5864 10279 5920
rect 10081 5722 10137 5778
rect 10223 5722 10279 5778
rect 10081 5580 10137 5636
rect 10223 5580 10279 5636
rect 10081 5438 10137 5494
rect 10223 5438 10279 5494
rect 10081 5296 10137 5352
rect 10223 5296 10279 5352
rect 10081 5154 10137 5210
rect 10223 5154 10279 5210
rect 10081 5012 10137 5068
rect 10223 5012 10279 5068
rect 10081 4870 10137 4926
rect 10223 4870 10279 4926
rect 10081 4728 10137 4784
rect 10223 4728 10279 4784
rect 10081 4586 10137 4642
rect 10223 4586 10279 4642
rect 10081 4444 10137 4500
rect 10223 4444 10279 4500
rect 10081 4302 10137 4358
rect 10223 4302 10279 4358
rect 10081 4160 10137 4216
rect 10223 4160 10279 4216
rect 10081 4018 10137 4074
rect 10223 4018 10279 4074
rect 10081 3876 10137 3932
rect 10223 3876 10279 3932
rect 10081 3734 10137 3790
rect 10223 3734 10279 3790
rect 10081 3592 10137 3648
rect 10223 3592 10279 3648
rect 10081 3450 10137 3506
rect 10223 3450 10279 3506
rect 10081 3308 10137 3364
rect 10223 3308 10279 3364
rect 10081 3166 10137 3222
rect 10223 3166 10279 3222
rect 10081 3024 10137 3080
rect 10223 3024 10279 3080
rect 10081 2882 10137 2938
rect 10223 2882 10279 2938
rect 10081 2740 10137 2796
rect 10223 2740 10279 2796
rect 10081 2598 10137 2654
rect 10223 2598 10279 2654
rect 10081 2456 10137 2512
rect 10223 2456 10279 2512
rect 10081 2314 10137 2370
rect 10223 2314 10279 2370
rect 10081 2172 10137 2228
rect 10223 2172 10279 2228
rect 10081 2030 10137 2086
rect 10223 2030 10279 2086
rect 10081 1888 10137 1944
rect 10223 1888 10279 1944
rect 10081 1746 10137 1802
rect 10223 1746 10279 1802
rect 10081 1604 10137 1660
rect 10223 1604 10279 1660
rect 10081 1462 10137 1518
rect 10223 1462 10279 1518
rect 10081 1320 10137 1376
rect 10223 1320 10279 1376
rect 10081 1178 10137 1234
rect 10223 1178 10279 1234
rect 10081 1036 10137 1092
rect 10223 1036 10279 1092
rect 10081 894 10137 950
rect 10223 894 10279 950
rect 10081 752 10137 808
rect 10223 752 10279 808
rect 10081 610 10137 666
rect 10223 610 10279 666
rect 10081 468 10137 524
rect 10223 468 10279 524
rect 10622 12254 10678 12310
rect 10764 12254 10820 12310
rect 10622 12112 10678 12168
rect 10764 12112 10820 12168
rect 10622 11970 10678 12026
rect 10764 11970 10820 12026
rect 10622 11828 10678 11884
rect 10764 11828 10820 11884
rect 10622 11686 10678 11742
rect 10764 11686 10820 11742
rect 10622 11544 10678 11600
rect 10764 11544 10820 11600
rect 10622 11402 10678 11458
rect 10764 11402 10820 11458
rect 10622 11260 10678 11316
rect 10764 11260 10820 11316
rect 10622 11118 10678 11174
rect 10764 11118 10820 11174
rect 10622 10976 10678 11032
rect 10764 10976 10820 11032
rect 10622 10834 10678 10890
rect 10764 10834 10820 10890
rect 10622 10692 10678 10748
rect 10764 10692 10820 10748
rect 10622 10550 10678 10606
rect 10764 10550 10820 10606
rect 10622 10408 10678 10464
rect 10764 10408 10820 10464
rect 10622 10266 10678 10322
rect 10764 10266 10820 10322
rect 10622 10124 10678 10180
rect 10764 10124 10820 10180
rect 10622 9982 10678 10038
rect 10764 9982 10820 10038
rect 10622 9840 10678 9896
rect 10764 9840 10820 9896
rect 10622 9698 10678 9754
rect 10764 9698 10820 9754
rect 10622 9556 10678 9612
rect 10764 9556 10820 9612
rect 10622 9414 10678 9470
rect 10764 9414 10820 9470
rect 10622 9272 10678 9328
rect 10764 9272 10820 9328
rect 10622 9130 10678 9186
rect 10764 9130 10820 9186
rect 10622 8988 10678 9044
rect 10764 8988 10820 9044
rect 10622 8846 10678 8902
rect 10764 8846 10820 8902
rect 10622 8704 10678 8760
rect 10764 8704 10820 8760
rect 10622 8562 10678 8618
rect 10764 8562 10820 8618
rect 10622 8420 10678 8476
rect 10764 8420 10820 8476
rect 10622 8278 10678 8334
rect 10764 8278 10820 8334
rect 10622 8136 10678 8192
rect 10764 8136 10820 8192
rect 10622 7994 10678 8050
rect 10764 7994 10820 8050
rect 10622 7852 10678 7908
rect 10764 7852 10820 7908
rect 10622 7710 10678 7766
rect 10764 7710 10820 7766
rect 10622 7568 10678 7624
rect 10764 7568 10820 7624
rect 10622 7426 10678 7482
rect 10764 7426 10820 7482
rect 10622 7284 10678 7340
rect 10764 7284 10820 7340
rect 10622 7142 10678 7198
rect 10764 7142 10820 7198
rect 10622 7000 10678 7056
rect 10764 7000 10820 7056
rect 10622 6858 10678 6914
rect 10764 6858 10820 6914
rect 10622 6716 10678 6772
rect 10764 6716 10820 6772
rect 10622 6574 10678 6630
rect 10764 6574 10820 6630
rect 10622 6432 10678 6488
rect 10764 6432 10820 6488
rect 10622 6290 10678 6346
rect 10764 6290 10820 6346
rect 10622 6148 10678 6204
rect 10764 6148 10820 6204
rect 10622 6006 10678 6062
rect 10764 6006 10820 6062
rect 10622 5864 10678 5920
rect 10764 5864 10820 5920
rect 10622 5722 10678 5778
rect 10764 5722 10820 5778
rect 10622 5580 10678 5636
rect 10764 5580 10820 5636
rect 10622 5438 10678 5494
rect 10764 5438 10820 5494
rect 10622 5296 10678 5352
rect 10764 5296 10820 5352
rect 10622 5154 10678 5210
rect 10764 5154 10820 5210
rect 10622 5012 10678 5068
rect 10764 5012 10820 5068
rect 10622 4870 10678 4926
rect 10764 4870 10820 4926
rect 10622 4728 10678 4784
rect 10764 4728 10820 4784
rect 10622 4586 10678 4642
rect 10764 4586 10820 4642
rect 10622 4444 10678 4500
rect 10764 4444 10820 4500
rect 10622 4302 10678 4358
rect 10764 4302 10820 4358
rect 10622 4160 10678 4216
rect 10764 4160 10820 4216
rect 10622 4018 10678 4074
rect 10764 4018 10820 4074
rect 10622 3876 10678 3932
rect 10764 3876 10820 3932
rect 10622 3734 10678 3790
rect 10764 3734 10820 3790
rect 10622 3592 10678 3648
rect 10764 3592 10820 3648
rect 10622 3450 10678 3506
rect 10764 3450 10820 3506
rect 10622 3308 10678 3364
rect 10764 3308 10820 3364
rect 10622 3166 10678 3222
rect 10764 3166 10820 3222
rect 10622 3024 10678 3080
rect 10764 3024 10820 3080
rect 10622 2882 10678 2938
rect 10764 2882 10820 2938
rect 10622 2740 10678 2796
rect 10764 2740 10820 2796
rect 10622 2598 10678 2654
rect 10764 2598 10820 2654
rect 10622 2456 10678 2512
rect 10764 2456 10820 2512
rect 10622 2314 10678 2370
rect 10764 2314 10820 2370
rect 10622 2172 10678 2228
rect 10764 2172 10820 2228
rect 10622 2030 10678 2086
rect 10764 2030 10820 2086
rect 10622 1888 10678 1944
rect 10764 1888 10820 1944
rect 10622 1746 10678 1802
rect 10764 1746 10820 1802
rect 10622 1604 10678 1660
rect 10764 1604 10820 1660
rect 10622 1462 10678 1518
rect 10764 1462 10820 1518
rect 10622 1320 10678 1376
rect 10764 1320 10820 1376
rect 10622 1178 10678 1234
rect 10764 1178 10820 1234
rect 10622 1036 10678 1092
rect 10764 1036 10820 1092
rect 10622 894 10678 950
rect 10764 894 10820 950
rect 10622 752 10678 808
rect 10764 752 10820 808
rect 10622 610 10678 666
rect 10764 610 10820 666
rect 10622 468 10678 524
rect 10764 468 10820 524
rect 11162 12254 11218 12310
rect 11304 12254 11360 12310
rect 11162 12112 11218 12168
rect 11304 12112 11360 12168
rect 11162 11970 11218 12026
rect 11304 11970 11360 12026
rect 11162 11828 11218 11884
rect 11304 11828 11360 11884
rect 11162 11686 11218 11742
rect 11304 11686 11360 11742
rect 11162 11544 11218 11600
rect 11304 11544 11360 11600
rect 11162 11402 11218 11458
rect 11304 11402 11360 11458
rect 11162 11260 11218 11316
rect 11304 11260 11360 11316
rect 11162 11118 11218 11174
rect 11304 11118 11360 11174
rect 11162 10976 11218 11032
rect 11304 10976 11360 11032
rect 11162 10834 11218 10890
rect 11304 10834 11360 10890
rect 11162 10692 11218 10748
rect 11304 10692 11360 10748
rect 11162 10550 11218 10606
rect 11304 10550 11360 10606
rect 11162 10408 11218 10464
rect 11304 10408 11360 10464
rect 11162 10266 11218 10322
rect 11304 10266 11360 10322
rect 11162 10124 11218 10180
rect 11304 10124 11360 10180
rect 11162 9982 11218 10038
rect 11304 9982 11360 10038
rect 11162 9840 11218 9896
rect 11304 9840 11360 9896
rect 11162 9698 11218 9754
rect 11304 9698 11360 9754
rect 11162 9556 11218 9612
rect 11304 9556 11360 9612
rect 11162 9414 11218 9470
rect 11304 9414 11360 9470
rect 11162 9272 11218 9328
rect 11304 9272 11360 9328
rect 11162 9130 11218 9186
rect 11304 9130 11360 9186
rect 11162 8988 11218 9044
rect 11304 8988 11360 9044
rect 11162 8846 11218 8902
rect 11304 8846 11360 8902
rect 11162 8704 11218 8760
rect 11304 8704 11360 8760
rect 11162 8562 11218 8618
rect 11304 8562 11360 8618
rect 11162 8420 11218 8476
rect 11304 8420 11360 8476
rect 11162 8278 11218 8334
rect 11304 8278 11360 8334
rect 11162 8136 11218 8192
rect 11304 8136 11360 8192
rect 11162 7994 11218 8050
rect 11304 7994 11360 8050
rect 11162 7852 11218 7908
rect 11304 7852 11360 7908
rect 11162 7710 11218 7766
rect 11304 7710 11360 7766
rect 11162 7568 11218 7624
rect 11304 7568 11360 7624
rect 11162 7426 11218 7482
rect 11304 7426 11360 7482
rect 11162 7284 11218 7340
rect 11304 7284 11360 7340
rect 11162 7142 11218 7198
rect 11304 7142 11360 7198
rect 11162 7000 11218 7056
rect 11304 7000 11360 7056
rect 11162 6858 11218 6914
rect 11304 6858 11360 6914
rect 11162 6716 11218 6772
rect 11304 6716 11360 6772
rect 11162 6574 11218 6630
rect 11304 6574 11360 6630
rect 11162 6432 11218 6488
rect 11304 6432 11360 6488
rect 11162 6290 11218 6346
rect 11304 6290 11360 6346
rect 11162 6148 11218 6204
rect 11304 6148 11360 6204
rect 11162 6006 11218 6062
rect 11304 6006 11360 6062
rect 11162 5864 11218 5920
rect 11304 5864 11360 5920
rect 11162 5722 11218 5778
rect 11304 5722 11360 5778
rect 11162 5580 11218 5636
rect 11304 5580 11360 5636
rect 11162 5438 11218 5494
rect 11304 5438 11360 5494
rect 11162 5296 11218 5352
rect 11304 5296 11360 5352
rect 11162 5154 11218 5210
rect 11304 5154 11360 5210
rect 11162 5012 11218 5068
rect 11304 5012 11360 5068
rect 11162 4870 11218 4926
rect 11304 4870 11360 4926
rect 11162 4728 11218 4784
rect 11304 4728 11360 4784
rect 11162 4586 11218 4642
rect 11304 4586 11360 4642
rect 11162 4444 11218 4500
rect 11304 4444 11360 4500
rect 11162 4302 11218 4358
rect 11304 4302 11360 4358
rect 11162 4160 11218 4216
rect 11304 4160 11360 4216
rect 11162 4018 11218 4074
rect 11304 4018 11360 4074
rect 11162 3876 11218 3932
rect 11304 3876 11360 3932
rect 11162 3734 11218 3790
rect 11304 3734 11360 3790
rect 11162 3592 11218 3648
rect 11304 3592 11360 3648
rect 11162 3450 11218 3506
rect 11304 3450 11360 3506
rect 11162 3308 11218 3364
rect 11304 3308 11360 3364
rect 11162 3166 11218 3222
rect 11304 3166 11360 3222
rect 11162 3024 11218 3080
rect 11304 3024 11360 3080
rect 11162 2882 11218 2938
rect 11304 2882 11360 2938
rect 11162 2740 11218 2796
rect 11304 2740 11360 2796
rect 11162 2598 11218 2654
rect 11304 2598 11360 2654
rect 11162 2456 11218 2512
rect 11304 2456 11360 2512
rect 11162 2314 11218 2370
rect 11304 2314 11360 2370
rect 11162 2172 11218 2228
rect 11304 2172 11360 2228
rect 11162 2030 11218 2086
rect 11304 2030 11360 2086
rect 11162 1888 11218 1944
rect 11304 1888 11360 1944
rect 11162 1746 11218 1802
rect 11304 1746 11360 1802
rect 11162 1604 11218 1660
rect 11304 1604 11360 1660
rect 11162 1462 11218 1518
rect 11304 1462 11360 1518
rect 11162 1320 11218 1376
rect 11304 1320 11360 1376
rect 11162 1178 11218 1234
rect 11304 1178 11360 1234
rect 11162 1036 11218 1092
rect 11304 1036 11360 1092
rect 11162 894 11218 950
rect 11304 894 11360 950
rect 11162 752 11218 808
rect 11304 752 11360 808
rect 11162 610 11218 666
rect 11304 610 11360 666
rect 11162 468 11218 524
rect 11304 468 11360 524
rect 11702 12254 11758 12310
rect 11844 12254 11900 12310
rect 11702 12112 11758 12168
rect 11844 12112 11900 12168
rect 11702 11970 11758 12026
rect 11844 11970 11900 12026
rect 11702 11828 11758 11884
rect 11844 11828 11900 11884
rect 11702 11686 11758 11742
rect 11844 11686 11900 11742
rect 11702 11544 11758 11600
rect 11844 11544 11900 11600
rect 11702 11402 11758 11458
rect 11844 11402 11900 11458
rect 11702 11260 11758 11316
rect 11844 11260 11900 11316
rect 11702 11118 11758 11174
rect 11844 11118 11900 11174
rect 11702 10976 11758 11032
rect 11844 10976 11900 11032
rect 11702 10834 11758 10890
rect 11844 10834 11900 10890
rect 11702 10692 11758 10748
rect 11844 10692 11900 10748
rect 11702 10550 11758 10606
rect 11844 10550 11900 10606
rect 11702 10408 11758 10464
rect 11844 10408 11900 10464
rect 11702 10266 11758 10322
rect 11844 10266 11900 10322
rect 11702 10124 11758 10180
rect 11844 10124 11900 10180
rect 11702 9982 11758 10038
rect 11844 9982 11900 10038
rect 11702 9840 11758 9896
rect 11844 9840 11900 9896
rect 11702 9698 11758 9754
rect 11844 9698 11900 9754
rect 11702 9556 11758 9612
rect 11844 9556 11900 9612
rect 11702 9414 11758 9470
rect 11844 9414 11900 9470
rect 11702 9272 11758 9328
rect 11844 9272 11900 9328
rect 11702 9130 11758 9186
rect 11844 9130 11900 9186
rect 11702 8988 11758 9044
rect 11844 8988 11900 9044
rect 11702 8846 11758 8902
rect 11844 8846 11900 8902
rect 11702 8704 11758 8760
rect 11844 8704 11900 8760
rect 11702 8562 11758 8618
rect 11844 8562 11900 8618
rect 11702 8420 11758 8476
rect 11844 8420 11900 8476
rect 11702 8278 11758 8334
rect 11844 8278 11900 8334
rect 11702 8136 11758 8192
rect 11844 8136 11900 8192
rect 11702 7994 11758 8050
rect 11844 7994 11900 8050
rect 11702 7852 11758 7908
rect 11844 7852 11900 7908
rect 11702 7710 11758 7766
rect 11844 7710 11900 7766
rect 11702 7568 11758 7624
rect 11844 7568 11900 7624
rect 11702 7426 11758 7482
rect 11844 7426 11900 7482
rect 11702 7284 11758 7340
rect 11844 7284 11900 7340
rect 11702 7142 11758 7198
rect 11844 7142 11900 7198
rect 11702 7000 11758 7056
rect 11844 7000 11900 7056
rect 11702 6858 11758 6914
rect 11844 6858 11900 6914
rect 11702 6716 11758 6772
rect 11844 6716 11900 6772
rect 11702 6574 11758 6630
rect 11844 6574 11900 6630
rect 11702 6432 11758 6488
rect 11844 6432 11900 6488
rect 11702 6290 11758 6346
rect 11844 6290 11900 6346
rect 11702 6148 11758 6204
rect 11844 6148 11900 6204
rect 11702 6006 11758 6062
rect 11844 6006 11900 6062
rect 11702 5864 11758 5920
rect 11844 5864 11900 5920
rect 11702 5722 11758 5778
rect 11844 5722 11900 5778
rect 11702 5580 11758 5636
rect 11844 5580 11900 5636
rect 11702 5438 11758 5494
rect 11844 5438 11900 5494
rect 11702 5296 11758 5352
rect 11844 5296 11900 5352
rect 11702 5154 11758 5210
rect 11844 5154 11900 5210
rect 11702 5012 11758 5068
rect 11844 5012 11900 5068
rect 11702 4870 11758 4926
rect 11844 4870 11900 4926
rect 11702 4728 11758 4784
rect 11844 4728 11900 4784
rect 11702 4586 11758 4642
rect 11844 4586 11900 4642
rect 11702 4444 11758 4500
rect 11844 4444 11900 4500
rect 11702 4302 11758 4358
rect 11844 4302 11900 4358
rect 11702 4160 11758 4216
rect 11844 4160 11900 4216
rect 11702 4018 11758 4074
rect 11844 4018 11900 4074
rect 11702 3876 11758 3932
rect 11844 3876 11900 3932
rect 11702 3734 11758 3790
rect 11844 3734 11900 3790
rect 11702 3592 11758 3648
rect 11844 3592 11900 3648
rect 11702 3450 11758 3506
rect 11844 3450 11900 3506
rect 11702 3308 11758 3364
rect 11844 3308 11900 3364
rect 11702 3166 11758 3222
rect 11844 3166 11900 3222
rect 11702 3024 11758 3080
rect 11844 3024 11900 3080
rect 11702 2882 11758 2938
rect 11844 2882 11900 2938
rect 11702 2740 11758 2796
rect 11844 2740 11900 2796
rect 11702 2598 11758 2654
rect 11844 2598 11900 2654
rect 11702 2456 11758 2512
rect 11844 2456 11900 2512
rect 11702 2314 11758 2370
rect 11844 2314 11900 2370
rect 11702 2172 11758 2228
rect 11844 2172 11900 2228
rect 11702 2030 11758 2086
rect 11844 2030 11900 2086
rect 11702 1888 11758 1944
rect 11844 1888 11900 1944
rect 11702 1746 11758 1802
rect 11844 1746 11900 1802
rect 11702 1604 11758 1660
rect 11844 1604 11900 1660
rect 11702 1462 11758 1518
rect 11844 1462 11900 1518
rect 11702 1320 11758 1376
rect 11844 1320 11900 1376
rect 11702 1178 11758 1234
rect 11844 1178 11900 1234
rect 11702 1036 11758 1092
rect 11844 1036 11900 1092
rect 11702 894 11758 950
rect 11844 894 11900 950
rect 11702 752 11758 808
rect 11844 752 11900 808
rect 11702 610 11758 666
rect 11844 610 11900 666
rect 11702 468 11758 524
rect 11844 468 11900 524
rect 12526 12302 12582 12358
rect 12650 12302 12706 12358
rect 12774 12302 12830 12358
rect 12898 12302 12954 12358
rect 13022 12302 13078 12358
rect 12526 12178 12582 12234
rect 12650 12178 12706 12234
rect 12774 12178 12830 12234
rect 12898 12178 12954 12234
rect 13022 12178 13078 12234
rect 12526 12054 12582 12110
rect 12650 12054 12706 12110
rect 12774 12054 12830 12110
rect 12898 12054 12954 12110
rect 13022 12054 13078 12110
rect 12526 11930 12582 11986
rect 12650 11930 12706 11986
rect 12774 11930 12830 11986
rect 12898 11930 12954 11986
rect 13022 11930 13078 11986
rect 12526 11806 12582 11862
rect 12650 11806 12706 11862
rect 12774 11806 12830 11862
rect 12898 11806 12954 11862
rect 13022 11806 13078 11862
rect 12526 11682 12582 11738
rect 12650 11682 12706 11738
rect 12774 11682 12830 11738
rect 12898 11682 12954 11738
rect 13022 11682 13078 11738
rect 12526 11558 12582 11614
rect 12650 11558 12706 11614
rect 12774 11558 12830 11614
rect 12898 11558 12954 11614
rect 13022 11558 13078 11614
rect 12526 11434 12582 11490
rect 12650 11434 12706 11490
rect 12774 11434 12830 11490
rect 12898 11434 12954 11490
rect 13022 11434 13078 11490
rect 12526 11310 12582 11366
rect 12650 11310 12706 11366
rect 12774 11310 12830 11366
rect 12898 11310 12954 11366
rect 13022 11310 13078 11366
rect 12526 11186 12582 11242
rect 12650 11186 12706 11242
rect 12774 11186 12830 11242
rect 12898 11186 12954 11242
rect 13022 11186 13078 11242
rect 12526 11062 12582 11118
rect 12650 11062 12706 11118
rect 12774 11062 12830 11118
rect 12898 11062 12954 11118
rect 13022 11062 13078 11118
rect 12526 10938 12582 10994
rect 12650 10938 12706 10994
rect 12774 10938 12830 10994
rect 12898 10938 12954 10994
rect 13022 10938 13078 10994
rect 12526 10814 12582 10870
rect 12650 10814 12706 10870
rect 12774 10814 12830 10870
rect 12898 10814 12954 10870
rect 13022 10814 13078 10870
rect 12526 10690 12582 10746
rect 12650 10690 12706 10746
rect 12774 10690 12830 10746
rect 12898 10690 12954 10746
rect 13022 10690 13078 10746
rect 12526 10566 12582 10622
rect 12650 10566 12706 10622
rect 12774 10566 12830 10622
rect 12898 10566 12954 10622
rect 13022 10566 13078 10622
rect 12526 10442 12582 10498
rect 12650 10442 12706 10498
rect 12774 10442 12830 10498
rect 12898 10442 12954 10498
rect 13022 10442 13078 10498
rect 12526 10318 12582 10374
rect 12650 10318 12706 10374
rect 12774 10318 12830 10374
rect 12898 10318 12954 10374
rect 13022 10318 13078 10374
rect 12526 10194 12582 10250
rect 12650 10194 12706 10250
rect 12774 10194 12830 10250
rect 12898 10194 12954 10250
rect 13022 10194 13078 10250
rect 12526 10070 12582 10126
rect 12650 10070 12706 10126
rect 12774 10070 12830 10126
rect 12898 10070 12954 10126
rect 13022 10070 13078 10126
rect 12526 9946 12582 10002
rect 12650 9946 12706 10002
rect 12774 9946 12830 10002
rect 12898 9946 12954 10002
rect 13022 9946 13078 10002
rect 12526 9822 12582 9878
rect 12650 9822 12706 9878
rect 12774 9822 12830 9878
rect 12898 9822 12954 9878
rect 13022 9822 13078 9878
rect 12526 9698 12582 9754
rect 12650 9698 12706 9754
rect 12774 9698 12830 9754
rect 12898 9698 12954 9754
rect 13022 9698 13078 9754
rect 12526 9574 12582 9630
rect 12650 9574 12706 9630
rect 12774 9574 12830 9630
rect 12898 9574 12954 9630
rect 13022 9574 13078 9630
rect 12526 9450 12582 9506
rect 12650 9450 12706 9506
rect 12774 9450 12830 9506
rect 12898 9450 12954 9506
rect 13022 9450 13078 9506
rect 12526 9326 12582 9382
rect 12650 9326 12706 9382
rect 12774 9326 12830 9382
rect 12898 9326 12954 9382
rect 13022 9326 13078 9382
rect 12526 9202 12582 9258
rect 12650 9202 12706 9258
rect 12774 9202 12830 9258
rect 12898 9202 12954 9258
rect 13022 9202 13078 9258
rect 12526 9078 12582 9134
rect 12650 9078 12706 9134
rect 12774 9078 12830 9134
rect 12898 9078 12954 9134
rect 13022 9078 13078 9134
rect 12526 8954 12582 9010
rect 12650 8954 12706 9010
rect 12774 8954 12830 9010
rect 12898 8954 12954 9010
rect 13022 8954 13078 9010
rect 12526 8830 12582 8886
rect 12650 8830 12706 8886
rect 12774 8830 12830 8886
rect 12898 8830 12954 8886
rect 13022 8830 13078 8886
rect 12526 8706 12582 8762
rect 12650 8706 12706 8762
rect 12774 8706 12830 8762
rect 12898 8706 12954 8762
rect 13022 8706 13078 8762
rect 12526 8582 12582 8638
rect 12650 8582 12706 8638
rect 12774 8582 12830 8638
rect 12898 8582 12954 8638
rect 13022 8582 13078 8638
rect 12526 8458 12582 8514
rect 12650 8458 12706 8514
rect 12774 8458 12830 8514
rect 12898 8458 12954 8514
rect 13022 8458 13078 8514
rect 12526 8334 12582 8390
rect 12650 8334 12706 8390
rect 12774 8334 12830 8390
rect 12898 8334 12954 8390
rect 13022 8334 13078 8390
rect 12526 8210 12582 8266
rect 12650 8210 12706 8266
rect 12774 8210 12830 8266
rect 12898 8210 12954 8266
rect 13022 8210 13078 8266
rect 12526 8086 12582 8142
rect 12650 8086 12706 8142
rect 12774 8086 12830 8142
rect 12898 8086 12954 8142
rect 13022 8086 13078 8142
rect 12526 7962 12582 8018
rect 12650 7962 12706 8018
rect 12774 7962 12830 8018
rect 12898 7962 12954 8018
rect 13022 7962 13078 8018
rect 12526 7838 12582 7894
rect 12650 7838 12706 7894
rect 12774 7838 12830 7894
rect 12898 7838 12954 7894
rect 13022 7838 13078 7894
rect 12526 7714 12582 7770
rect 12650 7714 12706 7770
rect 12774 7714 12830 7770
rect 12898 7714 12954 7770
rect 13022 7714 13078 7770
rect 12526 7590 12582 7646
rect 12650 7590 12706 7646
rect 12774 7590 12830 7646
rect 12898 7590 12954 7646
rect 13022 7590 13078 7646
rect 12526 7466 12582 7522
rect 12650 7466 12706 7522
rect 12774 7466 12830 7522
rect 12898 7466 12954 7522
rect 13022 7466 13078 7522
rect 12526 7342 12582 7398
rect 12650 7342 12706 7398
rect 12774 7342 12830 7398
rect 12898 7342 12954 7398
rect 13022 7342 13078 7398
rect 12526 7218 12582 7274
rect 12650 7218 12706 7274
rect 12774 7218 12830 7274
rect 12898 7218 12954 7274
rect 13022 7218 13078 7274
rect 12526 7094 12582 7150
rect 12650 7094 12706 7150
rect 12774 7094 12830 7150
rect 12898 7094 12954 7150
rect 13022 7094 13078 7150
rect 12526 6970 12582 7026
rect 12650 6970 12706 7026
rect 12774 6970 12830 7026
rect 12898 6970 12954 7026
rect 13022 6970 13078 7026
rect 12526 6846 12582 6902
rect 12650 6846 12706 6902
rect 12774 6846 12830 6902
rect 12898 6846 12954 6902
rect 13022 6846 13078 6902
rect 12526 6722 12582 6778
rect 12650 6722 12706 6778
rect 12774 6722 12830 6778
rect 12898 6722 12954 6778
rect 13022 6722 13078 6778
rect 12526 6598 12582 6654
rect 12650 6598 12706 6654
rect 12774 6598 12830 6654
rect 12898 6598 12954 6654
rect 13022 6598 13078 6654
rect 12526 6474 12582 6530
rect 12650 6474 12706 6530
rect 12774 6474 12830 6530
rect 12898 6474 12954 6530
rect 13022 6474 13078 6530
rect 12526 6350 12582 6406
rect 12650 6350 12706 6406
rect 12774 6350 12830 6406
rect 12898 6350 12954 6406
rect 13022 6350 13078 6406
rect 12526 6226 12582 6282
rect 12650 6226 12706 6282
rect 12774 6226 12830 6282
rect 12898 6226 12954 6282
rect 13022 6226 13078 6282
rect 12526 6102 12582 6158
rect 12650 6102 12706 6158
rect 12774 6102 12830 6158
rect 12898 6102 12954 6158
rect 13022 6102 13078 6158
rect 12526 5978 12582 6034
rect 12650 5978 12706 6034
rect 12774 5978 12830 6034
rect 12898 5978 12954 6034
rect 13022 5978 13078 6034
rect 12526 5854 12582 5910
rect 12650 5854 12706 5910
rect 12774 5854 12830 5910
rect 12898 5854 12954 5910
rect 13022 5854 13078 5910
rect 12526 5730 12582 5786
rect 12650 5730 12706 5786
rect 12774 5730 12830 5786
rect 12898 5730 12954 5786
rect 13022 5730 13078 5786
rect 12526 5606 12582 5662
rect 12650 5606 12706 5662
rect 12774 5606 12830 5662
rect 12898 5606 12954 5662
rect 13022 5606 13078 5662
rect 12526 5482 12582 5538
rect 12650 5482 12706 5538
rect 12774 5482 12830 5538
rect 12898 5482 12954 5538
rect 13022 5482 13078 5538
rect 12526 5358 12582 5414
rect 12650 5358 12706 5414
rect 12774 5358 12830 5414
rect 12898 5358 12954 5414
rect 13022 5358 13078 5414
rect 12526 5234 12582 5290
rect 12650 5234 12706 5290
rect 12774 5234 12830 5290
rect 12898 5234 12954 5290
rect 13022 5234 13078 5290
rect 12526 5110 12582 5166
rect 12650 5110 12706 5166
rect 12774 5110 12830 5166
rect 12898 5110 12954 5166
rect 13022 5110 13078 5166
rect 12526 4986 12582 5042
rect 12650 4986 12706 5042
rect 12774 4986 12830 5042
rect 12898 4986 12954 5042
rect 13022 4986 13078 5042
rect 12526 4862 12582 4918
rect 12650 4862 12706 4918
rect 12774 4862 12830 4918
rect 12898 4862 12954 4918
rect 13022 4862 13078 4918
rect 12526 4738 12582 4794
rect 12650 4738 12706 4794
rect 12774 4738 12830 4794
rect 12898 4738 12954 4794
rect 13022 4738 13078 4794
rect 12526 4614 12582 4670
rect 12650 4614 12706 4670
rect 12774 4614 12830 4670
rect 12898 4614 12954 4670
rect 13022 4614 13078 4670
rect 12526 4490 12582 4546
rect 12650 4490 12706 4546
rect 12774 4490 12830 4546
rect 12898 4490 12954 4546
rect 13022 4490 13078 4546
rect 12526 4366 12582 4422
rect 12650 4366 12706 4422
rect 12774 4366 12830 4422
rect 12898 4366 12954 4422
rect 13022 4366 13078 4422
rect 12526 4242 12582 4298
rect 12650 4242 12706 4298
rect 12774 4242 12830 4298
rect 12898 4242 12954 4298
rect 13022 4242 13078 4298
rect 12526 4118 12582 4174
rect 12650 4118 12706 4174
rect 12774 4118 12830 4174
rect 12898 4118 12954 4174
rect 13022 4118 13078 4174
rect 12526 3994 12582 4050
rect 12650 3994 12706 4050
rect 12774 3994 12830 4050
rect 12898 3994 12954 4050
rect 13022 3994 13078 4050
rect 12526 3870 12582 3926
rect 12650 3870 12706 3926
rect 12774 3870 12830 3926
rect 12898 3870 12954 3926
rect 13022 3870 13078 3926
rect 12526 3746 12582 3802
rect 12650 3746 12706 3802
rect 12774 3746 12830 3802
rect 12898 3746 12954 3802
rect 13022 3746 13078 3802
rect 12526 3622 12582 3678
rect 12650 3622 12706 3678
rect 12774 3622 12830 3678
rect 12898 3622 12954 3678
rect 13022 3622 13078 3678
rect 12526 3498 12582 3554
rect 12650 3498 12706 3554
rect 12774 3498 12830 3554
rect 12898 3498 12954 3554
rect 13022 3498 13078 3554
rect 12526 3374 12582 3430
rect 12650 3374 12706 3430
rect 12774 3374 12830 3430
rect 12898 3374 12954 3430
rect 13022 3374 13078 3430
rect 12526 3250 12582 3306
rect 12650 3250 12706 3306
rect 12774 3250 12830 3306
rect 12898 3250 12954 3306
rect 13022 3250 13078 3306
rect 12526 3126 12582 3182
rect 12650 3126 12706 3182
rect 12774 3126 12830 3182
rect 12898 3126 12954 3182
rect 13022 3126 13078 3182
rect 12526 3002 12582 3058
rect 12650 3002 12706 3058
rect 12774 3002 12830 3058
rect 12898 3002 12954 3058
rect 13022 3002 13078 3058
rect 12526 2878 12582 2934
rect 12650 2878 12706 2934
rect 12774 2878 12830 2934
rect 12898 2878 12954 2934
rect 13022 2878 13078 2934
rect 12526 2754 12582 2810
rect 12650 2754 12706 2810
rect 12774 2754 12830 2810
rect 12898 2754 12954 2810
rect 13022 2754 13078 2810
rect 12526 2630 12582 2686
rect 12650 2630 12706 2686
rect 12774 2630 12830 2686
rect 12898 2630 12954 2686
rect 13022 2630 13078 2686
rect 12526 2506 12582 2562
rect 12650 2506 12706 2562
rect 12774 2506 12830 2562
rect 12898 2506 12954 2562
rect 13022 2506 13078 2562
rect 12526 2382 12582 2438
rect 12650 2382 12706 2438
rect 12774 2382 12830 2438
rect 12898 2382 12954 2438
rect 13022 2382 13078 2438
rect 12526 2258 12582 2314
rect 12650 2258 12706 2314
rect 12774 2258 12830 2314
rect 12898 2258 12954 2314
rect 13022 2258 13078 2314
rect 12526 2134 12582 2190
rect 12650 2134 12706 2190
rect 12774 2134 12830 2190
rect 12898 2134 12954 2190
rect 13022 2134 13078 2190
rect 12526 2010 12582 2066
rect 12650 2010 12706 2066
rect 12774 2010 12830 2066
rect 12898 2010 12954 2066
rect 13022 2010 13078 2066
rect 12526 1886 12582 1942
rect 12650 1886 12706 1942
rect 12774 1886 12830 1942
rect 12898 1886 12954 1942
rect 13022 1886 13078 1942
rect 12526 1762 12582 1818
rect 12650 1762 12706 1818
rect 12774 1762 12830 1818
rect 12898 1762 12954 1818
rect 13022 1762 13078 1818
rect 12526 1638 12582 1694
rect 12650 1638 12706 1694
rect 12774 1638 12830 1694
rect 12898 1638 12954 1694
rect 13022 1638 13078 1694
rect 12526 1514 12582 1570
rect 12650 1514 12706 1570
rect 12774 1514 12830 1570
rect 12898 1514 12954 1570
rect 13022 1514 13078 1570
rect 12526 1390 12582 1446
rect 12650 1390 12706 1446
rect 12774 1390 12830 1446
rect 12898 1390 12954 1446
rect 13022 1390 13078 1446
rect 12526 1266 12582 1322
rect 12650 1266 12706 1322
rect 12774 1266 12830 1322
rect 12898 1266 12954 1322
rect 13022 1266 13078 1322
rect 12526 1142 12582 1198
rect 12650 1142 12706 1198
rect 12774 1142 12830 1198
rect 12898 1142 12954 1198
rect 13022 1142 13078 1198
rect 12526 1018 12582 1074
rect 12650 1018 12706 1074
rect 12774 1018 12830 1074
rect 12898 1018 12954 1074
rect 13022 1018 13078 1074
rect 12526 894 12582 950
rect 12650 894 12706 950
rect 12774 894 12830 950
rect 12898 894 12954 950
rect 13022 894 13078 950
rect 12526 770 12582 826
rect 12650 770 12706 826
rect 12774 770 12830 826
rect 12898 770 12954 826
rect 13022 770 13078 826
rect 12526 646 12582 702
rect 12650 646 12706 702
rect 12774 646 12830 702
rect 12898 646 12954 702
rect 13022 646 13078 702
rect 12526 522 12582 578
rect 12650 522 12706 578
rect 12774 522 12830 578
rect 12898 522 12954 578
rect 13022 522 13078 578
rect 12526 398 12582 454
rect 12650 398 12706 454
rect 12774 398 12830 454
rect 12898 398 12954 454
rect 13022 398 13078 454
rect -286 274 -230 330
rect -162 274 -106 330
rect -38 274 18 330
rect 86 274 142 330
rect 210 274 266 330
rect 415 246 471 302
rect 557 246 613 302
rect 699 246 755 302
rect 841 246 897 302
rect 983 246 1039 302
rect 1125 246 1181 302
rect 1267 246 1323 302
rect 1409 246 1465 302
rect 1551 246 1607 302
rect 1693 246 1749 302
rect 1835 246 1891 302
rect 1977 246 2033 302
rect 2119 246 2175 302
rect 2261 246 2317 302
rect 2403 246 2459 302
rect 2545 246 2601 302
rect 2687 246 2743 302
rect 2829 246 2885 302
rect 2971 246 3027 302
rect 3113 246 3169 302
rect 3255 246 3311 302
rect 3397 246 3453 302
rect 3539 246 3595 302
rect 3681 246 3737 302
rect 3823 246 3879 302
rect 3965 246 4021 302
rect 4107 246 4163 302
rect 4249 246 4305 302
rect 4391 246 4447 302
rect 4533 246 4589 302
rect 4675 246 4731 302
rect 4817 246 4873 302
rect 4959 246 5015 302
rect 5101 246 5157 302
rect 5243 246 5299 302
rect 5385 246 5441 302
rect 5527 246 5583 302
rect 5669 246 5725 302
rect 5811 246 5867 302
rect 5953 246 6009 302
rect 6095 246 6151 302
rect 6237 246 6293 302
rect 6379 246 6435 302
rect 6521 246 6577 302
rect 6663 246 6719 302
rect 6805 246 6861 302
rect 6947 246 7003 302
rect 7089 246 7145 302
rect 7231 246 7287 302
rect 7373 246 7429 302
rect 7515 246 7571 302
rect 7657 246 7713 302
rect 7799 246 7855 302
rect 7941 246 7997 302
rect 8083 246 8139 302
rect 8225 246 8281 302
rect 8367 246 8423 302
rect 8509 246 8565 302
rect 8651 246 8707 302
rect 8793 246 8849 302
rect 8935 246 8991 302
rect 9077 246 9133 302
rect 9219 246 9275 302
rect 9361 246 9417 302
rect 9503 246 9559 302
rect 9645 246 9701 302
rect 9787 246 9843 302
rect 9929 246 9985 302
rect 10071 246 10127 302
rect 10213 246 10269 302
rect 10355 246 10411 302
rect 10497 246 10553 302
rect 10639 246 10695 302
rect 10781 246 10837 302
rect 10923 246 10979 302
rect 11065 246 11121 302
rect 11207 246 11263 302
rect 11349 246 11405 302
rect 11491 246 11547 302
rect 11633 246 11689 302
rect 11775 246 11831 302
rect 11917 246 11973 302
rect 12059 246 12115 302
rect 12201 246 12257 302
rect 12343 246 12399 302
rect 12526 274 12582 330
rect 12650 274 12706 330
rect 12774 274 12830 330
rect 12898 274 12954 330
rect 13022 274 13078 330
rect -286 150 -230 206
rect -162 150 -106 206
rect -38 150 18 206
rect 86 150 142 206
rect 210 150 266 206
rect 415 104 471 160
rect 557 104 613 160
rect 699 104 755 160
rect 841 104 897 160
rect 983 104 1039 160
rect 1125 104 1181 160
rect 1267 104 1323 160
rect 1409 104 1465 160
rect 1551 104 1607 160
rect 1693 104 1749 160
rect 1835 104 1891 160
rect 1977 104 2033 160
rect 2119 104 2175 160
rect 2261 104 2317 160
rect 2403 104 2459 160
rect 2545 104 2601 160
rect 2687 104 2743 160
rect 2829 104 2885 160
rect 2971 104 3027 160
rect 3113 104 3169 160
rect 3255 104 3311 160
rect 3397 104 3453 160
rect 3539 104 3595 160
rect 3681 104 3737 160
rect 3823 104 3879 160
rect 3965 104 4021 160
rect 4107 104 4163 160
rect 4249 104 4305 160
rect 4391 104 4447 160
rect 4533 104 4589 160
rect 4675 104 4731 160
rect 4817 104 4873 160
rect 4959 104 5015 160
rect 5101 104 5157 160
rect 5243 104 5299 160
rect 5385 104 5441 160
rect 5527 104 5583 160
rect 5669 104 5725 160
rect 5811 104 5867 160
rect 5953 104 6009 160
rect 6095 104 6151 160
rect 6237 104 6293 160
rect 6379 104 6435 160
rect 6521 104 6577 160
rect 6663 104 6719 160
rect 6805 104 6861 160
rect 6947 104 7003 160
rect 7089 104 7145 160
rect 7231 104 7287 160
rect 7373 104 7429 160
rect 7515 104 7571 160
rect 7657 104 7713 160
rect 7799 104 7855 160
rect 7941 104 7997 160
rect 8083 104 8139 160
rect 8225 104 8281 160
rect 8367 104 8423 160
rect 8509 104 8565 160
rect 8651 104 8707 160
rect 8793 104 8849 160
rect 8935 104 8991 160
rect 9077 104 9133 160
rect 9219 104 9275 160
rect 9361 104 9417 160
rect 9503 104 9559 160
rect 9645 104 9701 160
rect 9787 104 9843 160
rect 9929 104 9985 160
rect 10071 104 10127 160
rect 10213 104 10269 160
rect 10355 104 10411 160
rect 10497 104 10553 160
rect 10639 104 10695 160
rect 10781 104 10837 160
rect 10923 104 10979 160
rect 11065 104 11121 160
rect 11207 104 11263 160
rect 11349 104 11405 160
rect 11491 104 11547 160
rect 11633 104 11689 160
rect 11775 104 11831 160
rect 11917 104 11973 160
rect 12059 104 12115 160
rect 12201 104 12257 160
rect 12343 104 12399 160
rect 12526 150 12582 206
rect 12650 150 12706 206
rect 12774 150 12830 206
rect 12898 150 12954 206
rect 13022 150 13078 206
<< metal3 >>
rect -400 12949 13200 13065
rect -400 12893 -254 12949
rect -198 12893 -130 12949
rect -74 12893 -6 12949
rect 50 12893 118 12949
rect 174 12893 242 12949
rect 298 12893 366 12949
rect 422 12893 490 12949
rect 546 12893 614 12949
rect 670 12893 738 12949
rect 794 12893 862 12949
rect 918 12893 986 12949
rect 1042 12893 1110 12949
rect 1166 12893 1234 12949
rect 1290 12893 1358 12949
rect 1414 12893 1482 12949
rect 1538 12893 1606 12949
rect 1662 12893 1730 12949
rect 1786 12893 1854 12949
rect 1910 12893 1978 12949
rect 2034 12893 2102 12949
rect 2158 12893 2226 12949
rect 2282 12893 2350 12949
rect 2406 12893 2474 12949
rect 2530 12893 2598 12949
rect 2654 12893 2722 12949
rect 2778 12893 2846 12949
rect 2902 12893 2970 12949
rect 3026 12893 3094 12949
rect 3150 12893 3218 12949
rect 3274 12893 3342 12949
rect 3398 12893 3466 12949
rect 3522 12893 3590 12949
rect 3646 12893 3714 12949
rect 3770 12893 3838 12949
rect 3894 12893 3962 12949
rect 4018 12893 4086 12949
rect 4142 12893 4210 12949
rect 4266 12893 4334 12949
rect 4390 12893 4458 12949
rect 4514 12893 4582 12949
rect 4638 12893 4706 12949
rect 4762 12893 4830 12949
rect 4886 12893 4954 12949
rect 5010 12893 5078 12949
rect 5134 12893 5202 12949
rect 5258 12893 5326 12949
rect 5382 12893 5450 12949
rect 5506 12893 5574 12949
rect 5630 12893 5698 12949
rect 5754 12893 5822 12949
rect 5878 12893 5946 12949
rect 6002 12893 6070 12949
rect 6126 12893 6194 12949
rect 6250 12893 6318 12949
rect 6374 12893 6442 12949
rect 6498 12893 6566 12949
rect 6622 12893 6690 12949
rect 6746 12893 6814 12949
rect 6870 12893 6938 12949
rect 6994 12893 7062 12949
rect 7118 12893 7186 12949
rect 7242 12893 7310 12949
rect 7366 12893 7434 12949
rect 7490 12893 7558 12949
rect 7614 12893 7682 12949
rect 7738 12893 7806 12949
rect 7862 12893 7930 12949
rect 7986 12893 8054 12949
rect 8110 12893 8178 12949
rect 8234 12893 8302 12949
rect 8358 12893 8426 12949
rect 8482 12893 8550 12949
rect 8606 12893 8674 12949
rect 8730 12893 8798 12949
rect 8854 12893 8922 12949
rect 8978 12893 9046 12949
rect 9102 12893 9170 12949
rect 9226 12893 9294 12949
rect 9350 12893 9418 12949
rect 9474 12893 9542 12949
rect 9598 12893 9666 12949
rect 9722 12893 9790 12949
rect 9846 12893 9914 12949
rect 9970 12893 10038 12949
rect 10094 12893 10162 12949
rect 10218 12893 10286 12949
rect 10342 12893 10410 12949
rect 10466 12893 10534 12949
rect 10590 12893 10658 12949
rect 10714 12893 10782 12949
rect 10838 12893 10906 12949
rect 10962 12893 11030 12949
rect 11086 12893 11154 12949
rect 11210 12893 11278 12949
rect 11334 12893 11402 12949
rect 11458 12893 11526 12949
rect 11582 12893 11650 12949
rect 11706 12893 11774 12949
rect 11830 12893 11898 12949
rect 11954 12893 12022 12949
rect 12078 12893 12146 12949
rect 12202 12893 12270 12949
rect 12326 12893 12394 12949
rect 12450 12893 12518 12949
rect 12574 12893 12642 12949
rect 12698 12893 12766 12949
rect 12822 12893 12890 12949
rect 12946 12893 13014 12949
rect 13070 12893 13200 12949
rect -400 12825 13200 12893
rect -400 12769 -254 12825
rect -198 12769 -130 12825
rect -74 12769 -6 12825
rect 50 12769 118 12825
rect 174 12769 242 12825
rect 298 12769 366 12825
rect 422 12769 490 12825
rect 546 12769 614 12825
rect 670 12769 738 12825
rect 794 12769 862 12825
rect 918 12769 986 12825
rect 1042 12769 1110 12825
rect 1166 12769 1234 12825
rect 1290 12769 1358 12825
rect 1414 12769 1482 12825
rect 1538 12769 1606 12825
rect 1662 12769 1730 12825
rect 1786 12769 1854 12825
rect 1910 12769 1978 12825
rect 2034 12769 2102 12825
rect 2158 12769 2226 12825
rect 2282 12769 2350 12825
rect 2406 12769 2474 12825
rect 2530 12769 2598 12825
rect 2654 12769 2722 12825
rect 2778 12769 2846 12825
rect 2902 12769 2970 12825
rect 3026 12769 3094 12825
rect 3150 12769 3218 12825
rect 3274 12769 3342 12825
rect 3398 12769 3466 12825
rect 3522 12769 3590 12825
rect 3646 12769 3714 12825
rect 3770 12769 3838 12825
rect 3894 12769 3962 12825
rect 4018 12769 4086 12825
rect 4142 12769 4210 12825
rect 4266 12769 4334 12825
rect 4390 12769 4458 12825
rect 4514 12769 4582 12825
rect 4638 12769 4706 12825
rect 4762 12769 4830 12825
rect 4886 12769 4954 12825
rect 5010 12769 5078 12825
rect 5134 12769 5202 12825
rect 5258 12769 5326 12825
rect 5382 12769 5450 12825
rect 5506 12769 5574 12825
rect 5630 12769 5698 12825
rect 5754 12769 5822 12825
rect 5878 12769 5946 12825
rect 6002 12769 6070 12825
rect 6126 12769 6194 12825
rect 6250 12769 6318 12825
rect 6374 12769 6442 12825
rect 6498 12769 6566 12825
rect 6622 12769 6690 12825
rect 6746 12769 6814 12825
rect 6870 12769 6938 12825
rect 6994 12769 7062 12825
rect 7118 12769 7186 12825
rect 7242 12769 7310 12825
rect 7366 12769 7434 12825
rect 7490 12769 7558 12825
rect 7614 12769 7682 12825
rect 7738 12769 7806 12825
rect 7862 12769 7930 12825
rect 7986 12769 8054 12825
rect 8110 12769 8178 12825
rect 8234 12769 8302 12825
rect 8358 12769 8426 12825
rect 8482 12769 8550 12825
rect 8606 12769 8674 12825
rect 8730 12769 8798 12825
rect 8854 12769 8922 12825
rect 8978 12769 9046 12825
rect 9102 12769 9170 12825
rect 9226 12769 9294 12825
rect 9350 12769 9418 12825
rect 9474 12769 9542 12825
rect 9598 12769 9666 12825
rect 9722 12769 9790 12825
rect 9846 12769 9914 12825
rect 9970 12769 10038 12825
rect 10094 12769 10162 12825
rect 10218 12769 10286 12825
rect 10342 12769 10410 12825
rect 10466 12769 10534 12825
rect 10590 12769 10658 12825
rect 10714 12769 10782 12825
rect 10838 12769 10906 12825
rect 10962 12769 11030 12825
rect 11086 12769 11154 12825
rect 11210 12769 11278 12825
rect 11334 12769 11402 12825
rect 11458 12769 11526 12825
rect 11582 12769 11650 12825
rect 11706 12769 11774 12825
rect 11830 12769 11898 12825
rect 11954 12769 12022 12825
rect 12078 12769 12146 12825
rect 12202 12769 12270 12825
rect 12326 12769 12394 12825
rect 12450 12769 12518 12825
rect 12574 12769 12642 12825
rect 12698 12769 12766 12825
rect 12822 12769 12890 12825
rect 12946 12769 13014 12825
rect 13070 12769 13200 12825
rect -400 12701 13200 12769
rect -400 12645 -254 12701
rect -198 12645 -130 12701
rect -74 12645 -6 12701
rect 50 12645 118 12701
rect 174 12645 242 12701
rect 298 12645 366 12701
rect 422 12645 490 12701
rect 546 12645 614 12701
rect 670 12645 738 12701
rect 794 12645 862 12701
rect 918 12645 986 12701
rect 1042 12645 1110 12701
rect 1166 12645 1234 12701
rect 1290 12645 1358 12701
rect 1414 12645 1482 12701
rect 1538 12645 1606 12701
rect 1662 12645 1730 12701
rect 1786 12645 1854 12701
rect 1910 12645 1978 12701
rect 2034 12645 2102 12701
rect 2158 12645 2226 12701
rect 2282 12645 2350 12701
rect 2406 12645 2474 12701
rect 2530 12645 2598 12701
rect 2654 12645 2722 12701
rect 2778 12645 2846 12701
rect 2902 12645 2970 12701
rect 3026 12645 3094 12701
rect 3150 12645 3218 12701
rect 3274 12645 3342 12701
rect 3398 12645 3466 12701
rect 3522 12645 3590 12701
rect 3646 12645 3714 12701
rect 3770 12645 3838 12701
rect 3894 12645 3962 12701
rect 4018 12645 4086 12701
rect 4142 12645 4210 12701
rect 4266 12645 4334 12701
rect 4390 12645 4458 12701
rect 4514 12645 4582 12701
rect 4638 12645 4706 12701
rect 4762 12645 4830 12701
rect 4886 12645 4954 12701
rect 5010 12645 5078 12701
rect 5134 12645 5202 12701
rect 5258 12645 5326 12701
rect 5382 12645 5450 12701
rect 5506 12645 5574 12701
rect 5630 12645 5698 12701
rect 5754 12645 5822 12701
rect 5878 12645 5946 12701
rect 6002 12645 6070 12701
rect 6126 12645 6194 12701
rect 6250 12645 6318 12701
rect 6374 12645 6442 12701
rect 6498 12645 6566 12701
rect 6622 12645 6690 12701
rect 6746 12645 6814 12701
rect 6870 12645 6938 12701
rect 6994 12645 7062 12701
rect 7118 12645 7186 12701
rect 7242 12645 7310 12701
rect 7366 12645 7434 12701
rect 7490 12645 7558 12701
rect 7614 12645 7682 12701
rect 7738 12645 7806 12701
rect 7862 12645 7930 12701
rect 7986 12645 8054 12701
rect 8110 12645 8178 12701
rect 8234 12645 8302 12701
rect 8358 12645 8426 12701
rect 8482 12645 8550 12701
rect 8606 12645 8674 12701
rect 8730 12645 8798 12701
rect 8854 12645 8922 12701
rect 8978 12645 9046 12701
rect 9102 12645 9170 12701
rect 9226 12645 9294 12701
rect 9350 12645 9418 12701
rect 9474 12645 9542 12701
rect 9598 12645 9666 12701
rect 9722 12645 9790 12701
rect 9846 12645 9914 12701
rect 9970 12645 10038 12701
rect 10094 12645 10162 12701
rect 10218 12645 10286 12701
rect 10342 12645 10410 12701
rect 10466 12645 10534 12701
rect 10590 12645 10658 12701
rect 10714 12645 10782 12701
rect 10838 12645 10906 12701
rect 10962 12645 11030 12701
rect 11086 12645 11154 12701
rect 11210 12645 11278 12701
rect 11334 12645 11402 12701
rect 11458 12645 11526 12701
rect 11582 12645 11650 12701
rect 11706 12645 11774 12701
rect 11830 12645 11898 12701
rect 11954 12645 12022 12701
rect 12078 12645 12146 12701
rect 12202 12645 12270 12701
rect 12326 12645 12394 12701
rect 12450 12645 12518 12701
rect 12574 12645 12642 12701
rect 12698 12645 12766 12701
rect 12822 12645 12890 12701
rect 12946 12645 13014 12701
rect 13070 12645 13200 12701
rect -400 12577 13200 12645
rect -400 12521 -254 12577
rect -198 12521 -130 12577
rect -74 12521 -6 12577
rect 50 12521 118 12577
rect 174 12521 242 12577
rect 298 12521 366 12577
rect 422 12521 490 12577
rect 546 12521 614 12577
rect 670 12521 738 12577
rect 794 12521 862 12577
rect 918 12521 986 12577
rect 1042 12521 1110 12577
rect 1166 12521 1234 12577
rect 1290 12521 1358 12577
rect 1414 12521 1482 12577
rect 1538 12521 1606 12577
rect 1662 12521 1730 12577
rect 1786 12521 1854 12577
rect 1910 12521 1978 12577
rect 2034 12521 2102 12577
rect 2158 12521 2226 12577
rect 2282 12521 2350 12577
rect 2406 12521 2474 12577
rect 2530 12521 2598 12577
rect 2654 12521 2722 12577
rect 2778 12521 2846 12577
rect 2902 12521 2970 12577
rect 3026 12521 3094 12577
rect 3150 12521 3218 12577
rect 3274 12521 3342 12577
rect 3398 12521 3466 12577
rect 3522 12521 3590 12577
rect 3646 12521 3714 12577
rect 3770 12521 3838 12577
rect 3894 12521 3962 12577
rect 4018 12521 4086 12577
rect 4142 12521 4210 12577
rect 4266 12521 4334 12577
rect 4390 12521 4458 12577
rect 4514 12521 4582 12577
rect 4638 12521 4706 12577
rect 4762 12521 4830 12577
rect 4886 12521 4954 12577
rect 5010 12521 5078 12577
rect 5134 12521 5202 12577
rect 5258 12521 5326 12577
rect 5382 12521 5450 12577
rect 5506 12521 5574 12577
rect 5630 12521 5698 12577
rect 5754 12521 5822 12577
rect 5878 12521 5946 12577
rect 6002 12521 6070 12577
rect 6126 12521 6194 12577
rect 6250 12521 6318 12577
rect 6374 12521 6442 12577
rect 6498 12521 6566 12577
rect 6622 12521 6690 12577
rect 6746 12521 6814 12577
rect 6870 12521 6938 12577
rect 6994 12521 7062 12577
rect 7118 12521 7186 12577
rect 7242 12521 7310 12577
rect 7366 12521 7434 12577
rect 7490 12521 7558 12577
rect 7614 12521 7682 12577
rect 7738 12521 7806 12577
rect 7862 12521 7930 12577
rect 7986 12521 8054 12577
rect 8110 12521 8178 12577
rect 8234 12521 8302 12577
rect 8358 12521 8426 12577
rect 8482 12521 8550 12577
rect 8606 12521 8674 12577
rect 8730 12521 8798 12577
rect 8854 12521 8922 12577
rect 8978 12521 9046 12577
rect 9102 12521 9170 12577
rect 9226 12521 9294 12577
rect 9350 12521 9418 12577
rect 9474 12521 9542 12577
rect 9598 12521 9666 12577
rect 9722 12521 9790 12577
rect 9846 12521 9914 12577
rect 9970 12521 10038 12577
rect 10094 12521 10162 12577
rect 10218 12521 10286 12577
rect 10342 12521 10410 12577
rect 10466 12521 10534 12577
rect 10590 12521 10658 12577
rect 10714 12521 10782 12577
rect 10838 12521 10906 12577
rect 10962 12521 11030 12577
rect 11086 12521 11154 12577
rect 11210 12521 11278 12577
rect 11334 12521 11402 12577
rect 11458 12521 11526 12577
rect 11582 12521 11650 12577
rect 11706 12521 11774 12577
rect 11830 12521 11898 12577
rect 11954 12521 12022 12577
rect 12078 12521 12146 12577
rect 12202 12521 12270 12577
rect 12326 12521 12394 12577
rect 12450 12521 12518 12577
rect 12574 12521 12642 12577
rect 12698 12521 12766 12577
rect 12822 12521 12890 12577
rect 12946 12521 13014 12577
rect 13070 12521 13200 12577
rect -400 12358 13200 12521
rect -400 12302 -286 12358
rect -230 12302 -162 12358
rect -106 12302 -38 12358
rect 18 12302 86 12358
rect 142 12302 210 12358
rect 266 12320 12526 12358
rect 266 12302 400 12320
rect -400 12234 400 12302
rect -400 12178 -286 12234
rect -230 12178 -162 12234
rect -106 12178 -38 12234
rect 18 12178 86 12234
rect 142 12178 210 12234
rect 266 12178 400 12234
rect -400 12110 400 12178
rect -400 12054 -286 12110
rect -230 12054 -162 12110
rect -106 12054 -38 12110
rect 18 12054 86 12110
rect 142 12054 210 12110
rect 266 12054 400 12110
rect -400 11986 400 12054
rect -400 11930 -286 11986
rect -230 11930 -162 11986
rect -106 11930 -38 11986
rect 18 11930 86 11986
rect 142 11930 210 11986
rect 266 11930 400 11986
rect -400 11862 400 11930
rect -400 11806 -286 11862
rect -230 11806 -162 11862
rect -106 11806 -38 11862
rect 18 11806 86 11862
rect 142 11806 210 11862
rect 266 11806 400 11862
rect -400 11738 400 11806
rect -400 11682 -286 11738
rect -230 11682 -162 11738
rect -106 11682 -38 11738
rect 18 11682 86 11738
rect 142 11682 210 11738
rect 266 11682 400 11738
rect -400 11614 400 11682
rect -400 11558 -286 11614
rect -230 11558 -162 11614
rect -106 11558 -38 11614
rect 18 11558 86 11614
rect 142 11558 210 11614
rect 266 11558 400 11614
rect -400 11490 400 11558
rect -400 11434 -286 11490
rect -230 11434 -162 11490
rect -106 11434 -38 11490
rect 18 11434 86 11490
rect 142 11434 210 11490
rect 266 11434 400 11490
rect -400 11366 400 11434
rect -400 11310 -286 11366
rect -230 11310 -162 11366
rect -106 11310 -38 11366
rect 18 11310 86 11366
rect 142 11310 210 11366
rect 266 11310 400 11366
rect -400 11242 400 11310
rect -400 11186 -286 11242
rect -230 11186 -162 11242
rect -106 11186 -38 11242
rect 18 11186 86 11242
rect 142 11186 210 11242
rect 266 11186 400 11242
rect -400 11118 400 11186
rect -400 11062 -286 11118
rect -230 11062 -162 11118
rect -106 11062 -38 11118
rect 18 11062 86 11118
rect 142 11062 210 11118
rect 266 11062 400 11118
rect -400 10994 400 11062
rect -400 10938 -286 10994
rect -230 10938 -162 10994
rect -106 10938 -38 10994
rect 18 10938 86 10994
rect 142 10938 210 10994
rect 266 10938 400 10994
rect -400 10870 400 10938
rect -400 10814 -286 10870
rect -230 10814 -162 10870
rect -106 10814 -38 10870
rect 18 10814 86 10870
rect 142 10814 210 10870
rect 266 10814 400 10870
rect -400 10746 400 10814
rect -400 10690 -286 10746
rect -230 10690 -162 10746
rect -106 10690 -38 10746
rect 18 10690 86 10746
rect 142 10690 210 10746
rect 266 10690 400 10746
rect -400 10622 400 10690
rect -400 10566 -286 10622
rect -230 10566 -162 10622
rect -106 10566 -38 10622
rect 18 10566 86 10622
rect 142 10566 210 10622
rect 266 10566 400 10622
rect -400 10498 400 10566
rect -400 10442 -286 10498
rect -230 10442 -162 10498
rect -106 10442 -38 10498
rect 18 10442 86 10498
rect 142 10442 210 10498
rect 266 10442 400 10498
rect -400 10374 400 10442
rect -400 10318 -286 10374
rect -230 10318 -162 10374
rect -106 10318 -38 10374
rect 18 10318 86 10374
rect 142 10318 210 10374
rect 266 10318 400 10374
rect -400 10250 400 10318
rect -400 10194 -286 10250
rect -230 10194 -162 10250
rect -106 10194 -38 10250
rect 18 10194 86 10250
rect 142 10194 210 10250
rect 266 10194 400 10250
rect -400 10126 400 10194
rect -400 10070 -286 10126
rect -230 10070 -162 10126
rect -106 10070 -38 10126
rect 18 10070 86 10126
rect 142 10070 210 10126
rect 266 10070 400 10126
rect -400 10002 400 10070
rect -400 9946 -286 10002
rect -230 9946 -162 10002
rect -106 9946 -38 10002
rect 18 9946 86 10002
rect 142 9946 210 10002
rect 266 9946 400 10002
rect -400 9878 400 9946
rect -400 9822 -286 9878
rect -230 9822 -162 9878
rect -106 9822 -38 9878
rect 18 9822 86 9878
rect 142 9822 210 9878
rect 266 9822 400 9878
rect -400 9754 400 9822
rect -400 9698 -286 9754
rect -230 9698 -162 9754
rect -106 9698 -38 9754
rect 18 9698 86 9754
rect 142 9698 210 9754
rect 266 9698 400 9754
rect -400 9630 400 9698
rect -400 9574 -286 9630
rect -230 9574 -162 9630
rect -106 9574 -38 9630
rect 18 9574 86 9630
rect 142 9574 210 9630
rect 266 9574 400 9630
rect -400 9506 400 9574
rect -400 9450 -286 9506
rect -230 9450 -162 9506
rect -106 9450 -38 9506
rect 18 9450 86 9506
rect 142 9450 210 9506
rect 266 9450 400 9506
rect -400 9382 400 9450
rect -400 9326 -286 9382
rect -230 9326 -162 9382
rect -106 9326 -38 9382
rect 18 9326 86 9382
rect 142 9326 210 9382
rect 266 9326 400 9382
rect -400 9258 400 9326
rect -400 9202 -286 9258
rect -230 9202 -162 9258
rect -106 9202 -38 9258
rect 18 9202 86 9258
rect 142 9202 210 9258
rect 266 9202 400 9258
rect -400 9134 400 9202
rect -400 9078 -286 9134
rect -230 9078 -162 9134
rect -106 9078 -38 9134
rect 18 9078 86 9134
rect 142 9078 210 9134
rect 266 9078 400 9134
rect -400 9010 400 9078
rect -400 8954 -286 9010
rect -230 8954 -162 9010
rect -106 8954 -38 9010
rect 18 8954 86 9010
rect 142 8954 210 9010
rect 266 8954 400 9010
rect -400 8886 400 8954
rect -400 8830 -286 8886
rect -230 8830 -162 8886
rect -106 8830 -38 8886
rect 18 8830 86 8886
rect 142 8830 210 8886
rect 266 8830 400 8886
rect -400 8762 400 8830
rect -400 8706 -286 8762
rect -230 8706 -162 8762
rect -106 8706 -38 8762
rect 18 8706 86 8762
rect 142 8706 210 8762
rect 266 8706 400 8762
rect -400 8638 400 8706
rect -400 8582 -286 8638
rect -230 8582 -162 8638
rect -106 8582 -38 8638
rect 18 8582 86 8638
rect 142 8582 210 8638
rect 266 8582 400 8638
rect -400 8514 400 8582
rect -400 8458 -286 8514
rect -230 8458 -162 8514
rect -106 8458 -38 8514
rect 18 8458 86 8514
rect 142 8458 210 8514
rect 266 8458 400 8514
rect -400 8390 400 8458
rect -400 8334 -286 8390
rect -230 8334 -162 8390
rect -106 8334 -38 8390
rect 18 8334 86 8390
rect 142 8334 210 8390
rect 266 8334 400 8390
rect -400 8266 400 8334
rect -400 8210 -286 8266
rect -230 8210 -162 8266
rect -106 8210 -38 8266
rect 18 8210 86 8266
rect 142 8210 210 8266
rect 266 8210 400 8266
rect -400 8142 400 8210
rect -400 8086 -286 8142
rect -230 8086 -162 8142
rect -106 8086 -38 8142
rect 18 8086 86 8142
rect 142 8086 210 8142
rect 266 8086 400 8142
rect -400 8018 400 8086
rect -400 7962 -286 8018
rect -230 7962 -162 8018
rect -106 7962 -38 8018
rect 18 7962 86 8018
rect 142 7962 210 8018
rect 266 7962 400 8018
rect -400 7894 400 7962
rect -400 7838 -286 7894
rect -230 7838 -162 7894
rect -106 7838 -38 7894
rect 18 7838 86 7894
rect 142 7838 210 7894
rect 266 7838 400 7894
rect -400 7770 400 7838
rect -400 7714 -286 7770
rect -230 7714 -162 7770
rect -106 7714 -38 7770
rect 18 7714 86 7770
rect 142 7714 210 7770
rect 266 7714 400 7770
rect -400 7646 400 7714
rect -400 7590 -286 7646
rect -230 7590 -162 7646
rect -106 7590 -38 7646
rect 18 7590 86 7646
rect 142 7590 210 7646
rect 266 7590 400 7646
rect -400 7522 400 7590
rect -400 7466 -286 7522
rect -230 7466 -162 7522
rect -106 7466 -38 7522
rect 18 7466 86 7522
rect 142 7466 210 7522
rect 266 7466 400 7522
rect -400 7398 400 7466
rect -400 7342 -286 7398
rect -230 7342 -162 7398
rect -106 7342 -38 7398
rect 18 7342 86 7398
rect 142 7342 210 7398
rect 266 7342 400 7398
rect -400 7274 400 7342
rect -400 7218 -286 7274
rect -230 7218 -162 7274
rect -106 7218 -38 7274
rect 18 7218 86 7274
rect 142 7218 210 7274
rect 266 7218 400 7274
rect -400 7150 400 7218
rect -400 7094 -286 7150
rect -230 7094 -162 7150
rect -106 7094 -38 7150
rect 18 7094 86 7150
rect 142 7094 210 7150
rect 266 7094 400 7150
rect -400 7026 400 7094
rect -400 6970 -286 7026
rect -230 6970 -162 7026
rect -106 6970 -38 7026
rect 18 6970 86 7026
rect 142 6970 210 7026
rect 266 6970 400 7026
rect -400 6902 400 6970
rect -400 6846 -286 6902
rect -230 6846 -162 6902
rect -106 6846 -38 6902
rect 18 6846 86 6902
rect 142 6846 210 6902
rect 266 6846 400 6902
rect -400 6778 400 6846
rect -400 6722 -286 6778
rect -230 6722 -162 6778
rect -106 6722 -38 6778
rect 18 6722 86 6778
rect 142 6722 210 6778
rect 266 6722 400 6778
rect -400 6654 400 6722
rect -400 6598 -286 6654
rect -230 6598 -162 6654
rect -106 6598 -38 6654
rect 18 6598 86 6654
rect 142 6598 210 6654
rect 266 6598 400 6654
rect -400 6530 400 6598
rect -400 6474 -286 6530
rect -230 6474 -162 6530
rect -106 6474 -38 6530
rect 18 6474 86 6530
rect 142 6474 210 6530
rect 266 6474 400 6530
rect -400 6406 400 6474
rect -400 6350 -286 6406
rect -230 6350 -162 6406
rect -106 6350 -38 6406
rect 18 6350 86 6406
rect 142 6350 210 6406
rect 266 6350 400 6406
rect -400 6282 400 6350
rect -400 6226 -286 6282
rect -230 6226 -162 6282
rect -106 6226 -38 6282
rect 18 6226 86 6282
rect 142 6226 210 6282
rect 266 6226 400 6282
rect -400 6158 400 6226
rect -400 6102 -286 6158
rect -230 6102 -162 6158
rect -106 6102 -38 6158
rect 18 6102 86 6158
rect 142 6102 210 6158
rect 266 6102 400 6158
rect -400 6034 400 6102
rect -400 5978 -286 6034
rect -230 5978 -162 6034
rect -106 5978 -38 6034
rect 18 5978 86 6034
rect 142 5978 210 6034
rect 266 5978 400 6034
rect -400 5910 400 5978
rect -400 5854 -286 5910
rect -230 5854 -162 5910
rect -106 5854 -38 5910
rect 18 5854 86 5910
rect 142 5854 210 5910
rect 266 5854 400 5910
rect -400 5786 400 5854
rect -400 5730 -286 5786
rect -230 5730 -162 5786
rect -106 5730 -38 5786
rect 18 5730 86 5786
rect 142 5730 210 5786
rect 266 5730 400 5786
rect -400 5662 400 5730
rect -400 5606 -286 5662
rect -230 5606 -162 5662
rect -106 5606 -38 5662
rect 18 5606 86 5662
rect 142 5606 210 5662
rect 266 5606 400 5662
rect -400 5538 400 5606
rect -400 5482 -286 5538
rect -230 5482 -162 5538
rect -106 5482 -38 5538
rect 18 5482 86 5538
rect 142 5482 210 5538
rect 266 5482 400 5538
rect -400 5414 400 5482
rect -400 5358 -286 5414
rect -230 5358 -162 5414
rect -106 5358 -38 5414
rect 18 5358 86 5414
rect 142 5358 210 5414
rect 266 5358 400 5414
rect -400 5290 400 5358
rect -400 5234 -286 5290
rect -230 5234 -162 5290
rect -106 5234 -38 5290
rect 18 5234 86 5290
rect 142 5234 210 5290
rect 266 5234 400 5290
rect -400 5166 400 5234
rect -400 5110 -286 5166
rect -230 5110 -162 5166
rect -106 5110 -38 5166
rect 18 5110 86 5166
rect 142 5110 210 5166
rect 266 5110 400 5166
rect -400 5042 400 5110
rect -400 4986 -286 5042
rect -230 4986 -162 5042
rect -106 4986 -38 5042
rect 18 4986 86 5042
rect 142 4986 210 5042
rect 266 4986 400 5042
rect -400 4918 400 4986
rect -400 4862 -286 4918
rect -230 4862 -162 4918
rect -106 4862 -38 4918
rect 18 4862 86 4918
rect 142 4862 210 4918
rect 266 4862 400 4918
rect -400 4794 400 4862
rect -400 4738 -286 4794
rect -230 4738 -162 4794
rect -106 4738 -38 4794
rect 18 4738 86 4794
rect 142 4738 210 4794
rect 266 4738 400 4794
rect -400 4670 400 4738
rect -400 4614 -286 4670
rect -230 4614 -162 4670
rect -106 4614 -38 4670
rect 18 4614 86 4670
rect 142 4614 210 4670
rect 266 4614 400 4670
rect -400 4546 400 4614
rect -400 4490 -286 4546
rect -230 4490 -162 4546
rect -106 4490 -38 4546
rect 18 4490 86 4546
rect 142 4490 210 4546
rect 266 4490 400 4546
rect -400 4422 400 4490
rect -400 4366 -286 4422
rect -230 4366 -162 4422
rect -106 4366 -38 4422
rect 18 4366 86 4422
rect 142 4366 210 4422
rect 266 4366 400 4422
rect -400 4298 400 4366
rect -400 4242 -286 4298
rect -230 4242 -162 4298
rect -106 4242 -38 4298
rect 18 4242 86 4298
rect 142 4242 210 4298
rect 266 4242 400 4298
rect -400 4174 400 4242
rect -400 4118 -286 4174
rect -230 4118 -162 4174
rect -106 4118 -38 4174
rect 18 4118 86 4174
rect 142 4118 210 4174
rect 266 4118 400 4174
rect -400 4050 400 4118
rect -400 3994 -286 4050
rect -230 3994 -162 4050
rect -106 3994 -38 4050
rect 18 3994 86 4050
rect 142 3994 210 4050
rect 266 3994 400 4050
rect -400 3926 400 3994
rect -400 3870 -286 3926
rect -230 3870 -162 3926
rect -106 3870 -38 3926
rect 18 3870 86 3926
rect 142 3870 210 3926
rect 266 3870 400 3926
rect -400 3802 400 3870
rect -400 3746 -286 3802
rect -230 3746 -162 3802
rect -106 3746 -38 3802
rect 18 3746 86 3802
rect 142 3746 210 3802
rect 266 3746 400 3802
rect -400 3678 400 3746
rect -400 3622 -286 3678
rect -230 3622 -162 3678
rect -106 3622 -38 3678
rect 18 3622 86 3678
rect 142 3622 210 3678
rect 266 3622 400 3678
rect -400 3554 400 3622
rect -400 3498 -286 3554
rect -230 3498 -162 3554
rect -106 3498 -38 3554
rect 18 3498 86 3554
rect 142 3498 210 3554
rect 266 3498 400 3554
rect -400 3430 400 3498
rect -400 3374 -286 3430
rect -230 3374 -162 3430
rect -106 3374 -38 3430
rect 18 3374 86 3430
rect 142 3374 210 3430
rect 266 3374 400 3430
rect -400 3306 400 3374
rect -400 3250 -286 3306
rect -230 3250 -162 3306
rect -106 3250 -38 3306
rect 18 3250 86 3306
rect 142 3250 210 3306
rect 266 3250 400 3306
rect -400 3182 400 3250
rect -400 3126 -286 3182
rect -230 3126 -162 3182
rect -106 3126 -38 3182
rect 18 3126 86 3182
rect 142 3126 210 3182
rect 266 3126 400 3182
rect -400 3058 400 3126
rect -400 3002 -286 3058
rect -230 3002 -162 3058
rect -106 3002 -38 3058
rect 18 3002 86 3058
rect 142 3002 210 3058
rect 266 3002 400 3058
rect -400 2934 400 3002
rect -400 2878 -286 2934
rect -230 2878 -162 2934
rect -106 2878 -38 2934
rect 18 2878 86 2934
rect 142 2878 210 2934
rect 266 2878 400 2934
rect -400 2810 400 2878
rect -400 2754 -286 2810
rect -230 2754 -162 2810
rect -106 2754 -38 2810
rect 18 2754 86 2810
rect 142 2754 210 2810
rect 266 2754 400 2810
rect -400 2686 400 2754
rect -400 2630 -286 2686
rect -230 2630 -162 2686
rect -106 2630 -38 2686
rect 18 2630 86 2686
rect 142 2630 210 2686
rect 266 2630 400 2686
rect -400 2562 400 2630
rect -400 2506 -286 2562
rect -230 2506 -162 2562
rect -106 2506 -38 2562
rect 18 2506 86 2562
rect 142 2506 210 2562
rect 266 2506 400 2562
rect -400 2438 400 2506
rect -400 2382 -286 2438
rect -230 2382 -162 2438
rect -106 2382 -38 2438
rect 18 2382 86 2438
rect 142 2382 210 2438
rect 266 2382 400 2438
rect -400 2314 400 2382
rect -400 2258 -286 2314
rect -230 2258 -162 2314
rect -106 2258 -38 2314
rect 18 2258 86 2314
rect 142 2258 210 2314
rect 266 2258 400 2314
rect -400 2190 400 2258
rect -400 2134 -286 2190
rect -230 2134 -162 2190
rect -106 2134 -38 2190
rect 18 2134 86 2190
rect 142 2134 210 2190
rect 266 2134 400 2190
rect -400 2066 400 2134
rect -400 2010 -286 2066
rect -230 2010 -162 2066
rect -106 2010 -38 2066
rect 18 2010 86 2066
rect 142 2010 210 2066
rect 266 2010 400 2066
rect -400 1942 400 2010
rect -400 1886 -286 1942
rect -230 1886 -162 1942
rect -106 1886 -38 1942
rect 18 1886 86 1942
rect 142 1886 210 1942
rect 266 1886 400 1942
rect -400 1818 400 1886
rect -400 1762 -286 1818
rect -230 1762 -162 1818
rect -106 1762 -38 1818
rect 18 1762 86 1818
rect 142 1762 210 1818
rect 266 1762 400 1818
rect -400 1694 400 1762
rect -400 1638 -286 1694
rect -230 1638 -162 1694
rect -106 1638 -38 1694
rect 18 1638 86 1694
rect 142 1638 210 1694
rect 266 1638 400 1694
rect -400 1570 400 1638
rect -400 1514 -286 1570
rect -230 1514 -162 1570
rect -106 1514 -38 1570
rect 18 1514 86 1570
rect 142 1514 210 1570
rect 266 1514 400 1570
rect -400 1446 400 1514
rect -400 1390 -286 1446
rect -230 1390 -162 1446
rect -106 1390 -38 1446
rect 18 1390 86 1446
rect 142 1390 210 1446
rect 266 1390 400 1446
rect -400 1322 400 1390
rect -400 1266 -286 1322
rect -230 1266 -162 1322
rect -106 1266 -38 1322
rect 18 1266 86 1322
rect 142 1266 210 1322
rect 266 1266 400 1322
rect -400 1198 400 1266
rect -400 1142 -286 1198
rect -230 1142 -162 1198
rect -106 1142 -38 1198
rect 18 1142 86 1198
rect 142 1142 210 1198
rect 266 1142 400 1198
rect -400 1074 400 1142
rect -400 1018 -286 1074
rect -230 1018 -162 1074
rect -106 1018 -38 1074
rect 18 1018 86 1074
rect 142 1018 210 1074
rect 266 1018 400 1074
rect -400 950 400 1018
rect -400 894 -286 950
rect -230 894 -162 950
rect -106 894 -38 950
rect 18 894 86 950
rect 142 894 210 950
rect 266 894 400 950
rect -400 826 400 894
rect -400 770 -286 826
rect -230 770 -162 826
rect -106 770 -38 826
rect 18 770 86 826
rect 142 770 210 826
rect 266 770 400 826
rect -400 702 400 770
rect -400 646 -286 702
rect -230 646 -162 702
rect -106 646 -38 702
rect 18 646 86 702
rect 142 646 210 702
rect 266 646 400 702
rect -400 578 400 646
rect -400 522 -286 578
rect -230 522 -162 578
rect -106 522 -38 578
rect 18 522 86 578
rect 142 522 210 578
rect 266 522 400 578
rect -400 458 400 522
rect 830 12310 1170 12320
rect 830 12254 903 12310
rect 959 12254 1045 12310
rect 1101 12254 1170 12310
rect 830 12168 1170 12254
rect 830 12112 903 12168
rect 959 12112 1045 12168
rect 1101 12112 1170 12168
rect 830 12026 1170 12112
rect 830 11970 903 12026
rect 959 11970 1045 12026
rect 1101 11970 1170 12026
rect 830 11884 1170 11970
rect 830 11828 903 11884
rect 959 11828 1045 11884
rect 1101 11828 1170 11884
rect 830 11742 1170 11828
rect 830 11686 903 11742
rect 959 11686 1045 11742
rect 1101 11686 1170 11742
rect 830 11600 1170 11686
rect 830 11544 903 11600
rect 959 11544 1045 11600
rect 1101 11544 1170 11600
rect 830 11458 1170 11544
rect 830 11402 903 11458
rect 959 11402 1045 11458
rect 1101 11402 1170 11458
rect 830 11316 1170 11402
rect 830 11260 903 11316
rect 959 11260 1045 11316
rect 1101 11260 1170 11316
rect 830 11174 1170 11260
rect 830 11118 903 11174
rect 959 11118 1045 11174
rect 1101 11118 1170 11174
rect 830 11032 1170 11118
rect 830 10976 903 11032
rect 959 10976 1045 11032
rect 1101 10976 1170 11032
rect 830 10890 1170 10976
rect 830 10834 903 10890
rect 959 10834 1045 10890
rect 1101 10834 1170 10890
rect 830 10748 1170 10834
rect 830 10692 903 10748
rect 959 10692 1045 10748
rect 1101 10692 1170 10748
rect 830 10606 1170 10692
rect 830 10550 903 10606
rect 959 10550 1045 10606
rect 1101 10550 1170 10606
rect 830 10464 1170 10550
rect 830 10408 903 10464
rect 959 10408 1045 10464
rect 1101 10408 1170 10464
rect 830 10322 1170 10408
rect 830 10266 903 10322
rect 959 10266 1045 10322
rect 1101 10266 1170 10322
rect 830 10180 1170 10266
rect 830 10124 903 10180
rect 959 10124 1045 10180
rect 1101 10124 1170 10180
rect 830 10038 1170 10124
rect 830 9982 903 10038
rect 959 9982 1045 10038
rect 1101 9982 1170 10038
rect 830 9896 1170 9982
rect 830 9840 903 9896
rect 959 9840 1045 9896
rect 1101 9840 1170 9896
rect 830 9754 1170 9840
rect 830 9698 903 9754
rect 959 9698 1045 9754
rect 1101 9698 1170 9754
rect 830 9612 1170 9698
rect 830 9556 903 9612
rect 959 9556 1045 9612
rect 1101 9556 1170 9612
rect 830 9470 1170 9556
rect 830 9414 903 9470
rect 959 9414 1045 9470
rect 1101 9414 1170 9470
rect 830 9328 1170 9414
rect 830 9272 903 9328
rect 959 9272 1045 9328
rect 1101 9272 1170 9328
rect 830 9186 1170 9272
rect 830 9130 903 9186
rect 959 9130 1045 9186
rect 1101 9130 1170 9186
rect 830 9044 1170 9130
rect 830 8988 903 9044
rect 959 8988 1045 9044
rect 1101 8988 1170 9044
rect 830 8902 1170 8988
rect 830 8846 903 8902
rect 959 8846 1045 8902
rect 1101 8846 1170 8902
rect 830 8760 1170 8846
rect 830 8704 903 8760
rect 959 8704 1045 8760
rect 1101 8704 1170 8760
rect 830 8618 1170 8704
rect 830 8562 903 8618
rect 959 8562 1045 8618
rect 1101 8562 1170 8618
rect 830 8476 1170 8562
rect 830 8420 903 8476
rect 959 8420 1045 8476
rect 1101 8420 1170 8476
rect 830 8334 1170 8420
rect 830 8278 903 8334
rect 959 8278 1045 8334
rect 1101 8278 1170 8334
rect 830 8192 1170 8278
rect 830 8136 903 8192
rect 959 8136 1045 8192
rect 1101 8136 1170 8192
rect 830 8050 1170 8136
rect 830 7994 903 8050
rect 959 7994 1045 8050
rect 1101 7994 1170 8050
rect 830 7908 1170 7994
rect 830 7852 903 7908
rect 959 7852 1045 7908
rect 1101 7852 1170 7908
rect 830 7766 1170 7852
rect 830 7710 903 7766
rect 959 7710 1045 7766
rect 1101 7710 1170 7766
rect 830 7624 1170 7710
rect 830 7568 903 7624
rect 959 7568 1045 7624
rect 1101 7568 1170 7624
rect 830 7482 1170 7568
rect 830 7426 903 7482
rect 959 7426 1045 7482
rect 1101 7426 1170 7482
rect 830 7340 1170 7426
rect 830 7284 903 7340
rect 959 7284 1045 7340
rect 1101 7284 1170 7340
rect 830 7198 1170 7284
rect 830 7142 903 7198
rect 959 7142 1045 7198
rect 1101 7142 1170 7198
rect 830 7056 1170 7142
rect 830 7000 903 7056
rect 959 7000 1045 7056
rect 1101 7000 1170 7056
rect 830 6914 1170 7000
rect 830 6858 903 6914
rect 959 6858 1045 6914
rect 1101 6858 1170 6914
rect 830 6772 1170 6858
rect 830 6716 903 6772
rect 959 6716 1045 6772
rect 1101 6716 1170 6772
rect 830 6630 1170 6716
rect 830 6574 903 6630
rect 959 6574 1045 6630
rect 1101 6574 1170 6630
rect 830 6488 1170 6574
rect 830 6432 903 6488
rect 959 6432 1045 6488
rect 1101 6432 1170 6488
rect 830 6346 1170 6432
rect 830 6290 903 6346
rect 959 6290 1045 6346
rect 1101 6290 1170 6346
rect 830 6204 1170 6290
rect 830 6148 903 6204
rect 959 6148 1045 6204
rect 1101 6148 1170 6204
rect 830 6062 1170 6148
rect 830 6006 903 6062
rect 959 6006 1045 6062
rect 1101 6006 1170 6062
rect 830 5920 1170 6006
rect 830 5864 903 5920
rect 959 5864 1045 5920
rect 1101 5864 1170 5920
rect 830 5778 1170 5864
rect 830 5722 903 5778
rect 959 5722 1045 5778
rect 1101 5722 1170 5778
rect 830 5636 1170 5722
rect 830 5580 903 5636
rect 959 5580 1045 5636
rect 1101 5580 1170 5636
rect 830 5494 1170 5580
rect 830 5438 903 5494
rect 959 5438 1045 5494
rect 1101 5438 1170 5494
rect 830 5352 1170 5438
rect 830 5296 903 5352
rect 959 5296 1045 5352
rect 1101 5296 1170 5352
rect 830 5210 1170 5296
rect 830 5154 903 5210
rect 959 5154 1045 5210
rect 1101 5154 1170 5210
rect 830 5068 1170 5154
rect 830 5012 903 5068
rect 959 5012 1045 5068
rect 1101 5012 1170 5068
rect 830 4926 1170 5012
rect 830 4870 903 4926
rect 959 4870 1045 4926
rect 1101 4870 1170 4926
rect 830 4784 1170 4870
rect 830 4728 903 4784
rect 959 4728 1045 4784
rect 1101 4728 1170 4784
rect 830 4642 1170 4728
rect 830 4586 903 4642
rect 959 4586 1045 4642
rect 1101 4586 1170 4642
rect 830 4500 1170 4586
rect 830 4444 903 4500
rect 959 4444 1045 4500
rect 1101 4444 1170 4500
rect 830 4358 1170 4444
rect 830 4302 903 4358
rect 959 4302 1045 4358
rect 1101 4302 1170 4358
rect 830 4216 1170 4302
rect 830 4160 903 4216
rect 959 4160 1045 4216
rect 1101 4160 1170 4216
rect 830 4074 1170 4160
rect 830 4018 903 4074
rect 959 4018 1045 4074
rect 1101 4018 1170 4074
rect 830 3932 1170 4018
rect 830 3876 903 3932
rect 959 3876 1045 3932
rect 1101 3876 1170 3932
rect 830 3790 1170 3876
rect 830 3734 903 3790
rect 959 3734 1045 3790
rect 1101 3734 1170 3790
rect 830 3648 1170 3734
rect 830 3592 903 3648
rect 959 3592 1045 3648
rect 1101 3592 1170 3648
rect 830 3506 1170 3592
rect 830 3450 903 3506
rect 959 3450 1045 3506
rect 1101 3450 1170 3506
rect 830 3364 1170 3450
rect 830 3308 903 3364
rect 959 3308 1045 3364
rect 1101 3308 1170 3364
rect 830 3222 1170 3308
rect 830 3166 903 3222
rect 959 3166 1045 3222
rect 1101 3166 1170 3222
rect 830 3080 1170 3166
rect 830 3024 903 3080
rect 959 3024 1045 3080
rect 1101 3024 1170 3080
rect 830 2938 1170 3024
rect 830 2882 903 2938
rect 959 2882 1045 2938
rect 1101 2882 1170 2938
rect 830 2796 1170 2882
rect 830 2740 903 2796
rect 959 2740 1045 2796
rect 1101 2740 1170 2796
rect 830 2654 1170 2740
rect 830 2598 903 2654
rect 959 2598 1045 2654
rect 1101 2598 1170 2654
rect 830 2512 1170 2598
rect 830 2456 903 2512
rect 959 2456 1045 2512
rect 1101 2456 1170 2512
rect 830 2370 1170 2456
rect 830 2314 903 2370
rect 959 2314 1045 2370
rect 1101 2314 1170 2370
rect 830 2228 1170 2314
rect 830 2172 903 2228
rect 959 2172 1045 2228
rect 1101 2172 1170 2228
rect 830 2086 1170 2172
rect 830 2030 903 2086
rect 959 2030 1045 2086
rect 1101 2030 1170 2086
rect 830 1944 1170 2030
rect 830 1888 903 1944
rect 959 1888 1045 1944
rect 1101 1888 1170 1944
rect 830 1802 1170 1888
rect 830 1746 903 1802
rect 959 1746 1045 1802
rect 1101 1746 1170 1802
rect 830 1660 1170 1746
rect 830 1604 903 1660
rect 959 1604 1045 1660
rect 1101 1604 1170 1660
rect 830 1518 1170 1604
rect 830 1462 903 1518
rect 959 1462 1045 1518
rect 1101 1462 1170 1518
rect 830 1376 1170 1462
rect 830 1320 903 1376
rect 959 1320 1045 1376
rect 1101 1320 1170 1376
rect 830 1234 1170 1320
rect 830 1178 903 1234
rect 959 1178 1045 1234
rect 1101 1178 1170 1234
rect 830 1092 1170 1178
rect 830 1036 903 1092
rect 959 1036 1045 1092
rect 1101 1036 1170 1092
rect 830 950 1170 1036
rect 830 894 903 950
rect 959 894 1045 950
rect 1101 894 1170 950
rect 830 808 1170 894
rect 830 752 903 808
rect 959 752 1045 808
rect 1101 752 1170 808
rect 830 666 1170 752
rect 830 610 903 666
rect 959 610 1045 666
rect 1101 610 1170 666
rect 830 524 1170 610
rect 830 468 903 524
rect 959 468 1045 524
rect 1101 468 1170 524
rect 830 458 1170 468
rect 1370 12310 1710 12320
rect 1370 12254 1444 12310
rect 1500 12254 1586 12310
rect 1642 12254 1710 12310
rect 1370 12168 1710 12254
rect 1370 12112 1444 12168
rect 1500 12112 1586 12168
rect 1642 12112 1710 12168
rect 1370 12026 1710 12112
rect 1370 11970 1444 12026
rect 1500 11970 1586 12026
rect 1642 11970 1710 12026
rect 1370 11884 1710 11970
rect 1370 11828 1444 11884
rect 1500 11828 1586 11884
rect 1642 11828 1710 11884
rect 1370 11742 1710 11828
rect 1370 11686 1444 11742
rect 1500 11686 1586 11742
rect 1642 11686 1710 11742
rect 1370 11600 1710 11686
rect 1370 11544 1444 11600
rect 1500 11544 1586 11600
rect 1642 11544 1710 11600
rect 1370 11458 1710 11544
rect 1370 11402 1444 11458
rect 1500 11402 1586 11458
rect 1642 11402 1710 11458
rect 1370 11316 1710 11402
rect 1370 11260 1444 11316
rect 1500 11260 1586 11316
rect 1642 11260 1710 11316
rect 1370 11174 1710 11260
rect 1370 11118 1444 11174
rect 1500 11118 1586 11174
rect 1642 11118 1710 11174
rect 1370 11032 1710 11118
rect 1370 10976 1444 11032
rect 1500 10976 1586 11032
rect 1642 10976 1710 11032
rect 1370 10890 1710 10976
rect 1370 10834 1444 10890
rect 1500 10834 1586 10890
rect 1642 10834 1710 10890
rect 1370 10748 1710 10834
rect 1370 10692 1444 10748
rect 1500 10692 1586 10748
rect 1642 10692 1710 10748
rect 1370 10606 1710 10692
rect 1370 10550 1444 10606
rect 1500 10550 1586 10606
rect 1642 10550 1710 10606
rect 1370 10464 1710 10550
rect 1370 10408 1444 10464
rect 1500 10408 1586 10464
rect 1642 10408 1710 10464
rect 1370 10322 1710 10408
rect 1370 10266 1444 10322
rect 1500 10266 1586 10322
rect 1642 10266 1710 10322
rect 1370 10180 1710 10266
rect 1370 10124 1444 10180
rect 1500 10124 1586 10180
rect 1642 10124 1710 10180
rect 1370 10038 1710 10124
rect 1370 9982 1444 10038
rect 1500 9982 1586 10038
rect 1642 9982 1710 10038
rect 1370 9896 1710 9982
rect 1370 9840 1444 9896
rect 1500 9840 1586 9896
rect 1642 9840 1710 9896
rect 1370 9754 1710 9840
rect 1370 9698 1444 9754
rect 1500 9698 1586 9754
rect 1642 9698 1710 9754
rect 1370 9612 1710 9698
rect 1370 9556 1444 9612
rect 1500 9556 1586 9612
rect 1642 9556 1710 9612
rect 1370 9470 1710 9556
rect 1370 9414 1444 9470
rect 1500 9414 1586 9470
rect 1642 9414 1710 9470
rect 1370 9328 1710 9414
rect 1370 9272 1444 9328
rect 1500 9272 1586 9328
rect 1642 9272 1710 9328
rect 1370 9186 1710 9272
rect 1370 9130 1444 9186
rect 1500 9130 1586 9186
rect 1642 9130 1710 9186
rect 1370 9044 1710 9130
rect 1370 8988 1444 9044
rect 1500 8988 1586 9044
rect 1642 8988 1710 9044
rect 1370 8902 1710 8988
rect 1370 8846 1444 8902
rect 1500 8846 1586 8902
rect 1642 8846 1710 8902
rect 1370 8760 1710 8846
rect 1370 8704 1444 8760
rect 1500 8704 1586 8760
rect 1642 8704 1710 8760
rect 1370 8618 1710 8704
rect 1370 8562 1444 8618
rect 1500 8562 1586 8618
rect 1642 8562 1710 8618
rect 1370 8476 1710 8562
rect 1370 8420 1444 8476
rect 1500 8420 1586 8476
rect 1642 8420 1710 8476
rect 1370 8334 1710 8420
rect 1370 8278 1444 8334
rect 1500 8278 1586 8334
rect 1642 8278 1710 8334
rect 1370 8192 1710 8278
rect 1370 8136 1444 8192
rect 1500 8136 1586 8192
rect 1642 8136 1710 8192
rect 1370 8050 1710 8136
rect 1370 7994 1444 8050
rect 1500 7994 1586 8050
rect 1642 7994 1710 8050
rect 1370 7908 1710 7994
rect 1370 7852 1444 7908
rect 1500 7852 1586 7908
rect 1642 7852 1710 7908
rect 1370 7766 1710 7852
rect 1370 7710 1444 7766
rect 1500 7710 1586 7766
rect 1642 7710 1710 7766
rect 1370 7624 1710 7710
rect 1370 7568 1444 7624
rect 1500 7568 1586 7624
rect 1642 7568 1710 7624
rect 1370 7482 1710 7568
rect 1370 7426 1444 7482
rect 1500 7426 1586 7482
rect 1642 7426 1710 7482
rect 1370 7340 1710 7426
rect 1370 7284 1444 7340
rect 1500 7284 1586 7340
rect 1642 7284 1710 7340
rect 1370 7198 1710 7284
rect 1370 7142 1444 7198
rect 1500 7142 1586 7198
rect 1642 7142 1710 7198
rect 1370 7056 1710 7142
rect 1370 7000 1444 7056
rect 1500 7000 1586 7056
rect 1642 7000 1710 7056
rect 1370 6914 1710 7000
rect 1370 6858 1444 6914
rect 1500 6858 1586 6914
rect 1642 6858 1710 6914
rect 1370 6772 1710 6858
rect 1370 6716 1444 6772
rect 1500 6716 1586 6772
rect 1642 6716 1710 6772
rect 1370 6630 1710 6716
rect 1370 6574 1444 6630
rect 1500 6574 1586 6630
rect 1642 6574 1710 6630
rect 1370 6488 1710 6574
rect 1370 6432 1444 6488
rect 1500 6432 1586 6488
rect 1642 6432 1710 6488
rect 1370 6346 1710 6432
rect 1370 6290 1444 6346
rect 1500 6290 1586 6346
rect 1642 6290 1710 6346
rect 1370 6204 1710 6290
rect 1370 6148 1444 6204
rect 1500 6148 1586 6204
rect 1642 6148 1710 6204
rect 1370 6062 1710 6148
rect 1370 6006 1444 6062
rect 1500 6006 1586 6062
rect 1642 6006 1710 6062
rect 1370 5920 1710 6006
rect 1370 5864 1444 5920
rect 1500 5864 1586 5920
rect 1642 5864 1710 5920
rect 1370 5778 1710 5864
rect 1370 5722 1444 5778
rect 1500 5722 1586 5778
rect 1642 5722 1710 5778
rect 1370 5636 1710 5722
rect 1370 5580 1444 5636
rect 1500 5580 1586 5636
rect 1642 5580 1710 5636
rect 1370 5494 1710 5580
rect 1370 5438 1444 5494
rect 1500 5438 1586 5494
rect 1642 5438 1710 5494
rect 1370 5352 1710 5438
rect 1370 5296 1444 5352
rect 1500 5296 1586 5352
rect 1642 5296 1710 5352
rect 1370 5210 1710 5296
rect 1370 5154 1444 5210
rect 1500 5154 1586 5210
rect 1642 5154 1710 5210
rect 1370 5068 1710 5154
rect 1370 5012 1444 5068
rect 1500 5012 1586 5068
rect 1642 5012 1710 5068
rect 1370 4926 1710 5012
rect 1370 4870 1444 4926
rect 1500 4870 1586 4926
rect 1642 4870 1710 4926
rect 1370 4784 1710 4870
rect 1370 4728 1444 4784
rect 1500 4728 1586 4784
rect 1642 4728 1710 4784
rect 1370 4642 1710 4728
rect 1370 4586 1444 4642
rect 1500 4586 1586 4642
rect 1642 4586 1710 4642
rect 1370 4500 1710 4586
rect 1370 4444 1444 4500
rect 1500 4444 1586 4500
rect 1642 4444 1710 4500
rect 1370 4358 1710 4444
rect 1370 4302 1444 4358
rect 1500 4302 1586 4358
rect 1642 4302 1710 4358
rect 1370 4216 1710 4302
rect 1370 4160 1444 4216
rect 1500 4160 1586 4216
rect 1642 4160 1710 4216
rect 1370 4074 1710 4160
rect 1370 4018 1444 4074
rect 1500 4018 1586 4074
rect 1642 4018 1710 4074
rect 1370 3932 1710 4018
rect 1370 3876 1444 3932
rect 1500 3876 1586 3932
rect 1642 3876 1710 3932
rect 1370 3790 1710 3876
rect 1370 3734 1444 3790
rect 1500 3734 1586 3790
rect 1642 3734 1710 3790
rect 1370 3648 1710 3734
rect 1370 3592 1444 3648
rect 1500 3592 1586 3648
rect 1642 3592 1710 3648
rect 1370 3506 1710 3592
rect 1370 3450 1444 3506
rect 1500 3450 1586 3506
rect 1642 3450 1710 3506
rect 1370 3364 1710 3450
rect 1370 3308 1444 3364
rect 1500 3308 1586 3364
rect 1642 3308 1710 3364
rect 1370 3222 1710 3308
rect 1370 3166 1444 3222
rect 1500 3166 1586 3222
rect 1642 3166 1710 3222
rect 1370 3080 1710 3166
rect 1370 3024 1444 3080
rect 1500 3024 1586 3080
rect 1642 3024 1710 3080
rect 1370 2938 1710 3024
rect 1370 2882 1444 2938
rect 1500 2882 1586 2938
rect 1642 2882 1710 2938
rect 1370 2796 1710 2882
rect 1370 2740 1444 2796
rect 1500 2740 1586 2796
rect 1642 2740 1710 2796
rect 1370 2654 1710 2740
rect 1370 2598 1444 2654
rect 1500 2598 1586 2654
rect 1642 2598 1710 2654
rect 1370 2512 1710 2598
rect 1370 2456 1444 2512
rect 1500 2456 1586 2512
rect 1642 2456 1710 2512
rect 1370 2370 1710 2456
rect 1370 2314 1444 2370
rect 1500 2314 1586 2370
rect 1642 2314 1710 2370
rect 1370 2228 1710 2314
rect 1370 2172 1444 2228
rect 1500 2172 1586 2228
rect 1642 2172 1710 2228
rect 1370 2086 1710 2172
rect 1370 2030 1444 2086
rect 1500 2030 1586 2086
rect 1642 2030 1710 2086
rect 1370 1944 1710 2030
rect 1370 1888 1444 1944
rect 1500 1888 1586 1944
rect 1642 1888 1710 1944
rect 1370 1802 1710 1888
rect 1370 1746 1444 1802
rect 1500 1746 1586 1802
rect 1642 1746 1710 1802
rect 1370 1660 1710 1746
rect 1370 1604 1444 1660
rect 1500 1604 1586 1660
rect 1642 1604 1710 1660
rect 1370 1518 1710 1604
rect 1370 1462 1444 1518
rect 1500 1462 1586 1518
rect 1642 1462 1710 1518
rect 1370 1376 1710 1462
rect 1370 1320 1444 1376
rect 1500 1320 1586 1376
rect 1642 1320 1710 1376
rect 1370 1234 1710 1320
rect 1370 1178 1444 1234
rect 1500 1178 1586 1234
rect 1642 1178 1710 1234
rect 1370 1092 1710 1178
rect 1370 1036 1444 1092
rect 1500 1036 1586 1092
rect 1642 1036 1710 1092
rect 1370 950 1710 1036
rect 1370 894 1444 950
rect 1500 894 1586 950
rect 1642 894 1710 950
rect 1370 808 1710 894
rect 1370 752 1444 808
rect 1500 752 1586 808
rect 1642 752 1710 808
rect 1370 666 1710 752
rect 1370 610 1444 666
rect 1500 610 1586 666
rect 1642 610 1710 666
rect 1370 524 1710 610
rect 1370 468 1444 524
rect 1500 468 1586 524
rect 1642 468 1710 524
rect 1370 458 1710 468
rect 1910 12310 2250 12320
rect 1910 12254 1984 12310
rect 2040 12254 2126 12310
rect 2182 12254 2250 12310
rect 1910 12168 2250 12254
rect 1910 12112 1984 12168
rect 2040 12112 2126 12168
rect 2182 12112 2250 12168
rect 1910 12026 2250 12112
rect 1910 11970 1984 12026
rect 2040 11970 2126 12026
rect 2182 11970 2250 12026
rect 1910 11884 2250 11970
rect 1910 11828 1984 11884
rect 2040 11828 2126 11884
rect 2182 11828 2250 11884
rect 1910 11742 2250 11828
rect 1910 11686 1984 11742
rect 2040 11686 2126 11742
rect 2182 11686 2250 11742
rect 1910 11600 2250 11686
rect 1910 11544 1984 11600
rect 2040 11544 2126 11600
rect 2182 11544 2250 11600
rect 1910 11458 2250 11544
rect 1910 11402 1984 11458
rect 2040 11402 2126 11458
rect 2182 11402 2250 11458
rect 1910 11316 2250 11402
rect 1910 11260 1984 11316
rect 2040 11260 2126 11316
rect 2182 11260 2250 11316
rect 1910 11174 2250 11260
rect 1910 11118 1984 11174
rect 2040 11118 2126 11174
rect 2182 11118 2250 11174
rect 1910 11032 2250 11118
rect 1910 10976 1984 11032
rect 2040 10976 2126 11032
rect 2182 10976 2250 11032
rect 1910 10890 2250 10976
rect 1910 10834 1984 10890
rect 2040 10834 2126 10890
rect 2182 10834 2250 10890
rect 1910 10748 2250 10834
rect 1910 10692 1984 10748
rect 2040 10692 2126 10748
rect 2182 10692 2250 10748
rect 1910 10606 2250 10692
rect 1910 10550 1984 10606
rect 2040 10550 2126 10606
rect 2182 10550 2250 10606
rect 1910 10464 2250 10550
rect 1910 10408 1984 10464
rect 2040 10408 2126 10464
rect 2182 10408 2250 10464
rect 1910 10322 2250 10408
rect 1910 10266 1984 10322
rect 2040 10266 2126 10322
rect 2182 10266 2250 10322
rect 1910 10180 2250 10266
rect 1910 10124 1984 10180
rect 2040 10124 2126 10180
rect 2182 10124 2250 10180
rect 1910 10038 2250 10124
rect 1910 9982 1984 10038
rect 2040 9982 2126 10038
rect 2182 9982 2250 10038
rect 1910 9896 2250 9982
rect 1910 9840 1984 9896
rect 2040 9840 2126 9896
rect 2182 9840 2250 9896
rect 1910 9754 2250 9840
rect 1910 9698 1984 9754
rect 2040 9698 2126 9754
rect 2182 9698 2250 9754
rect 1910 9612 2250 9698
rect 1910 9556 1984 9612
rect 2040 9556 2126 9612
rect 2182 9556 2250 9612
rect 1910 9470 2250 9556
rect 1910 9414 1984 9470
rect 2040 9414 2126 9470
rect 2182 9414 2250 9470
rect 1910 9328 2250 9414
rect 1910 9272 1984 9328
rect 2040 9272 2126 9328
rect 2182 9272 2250 9328
rect 1910 9186 2250 9272
rect 1910 9130 1984 9186
rect 2040 9130 2126 9186
rect 2182 9130 2250 9186
rect 1910 9044 2250 9130
rect 1910 8988 1984 9044
rect 2040 8988 2126 9044
rect 2182 8988 2250 9044
rect 1910 8902 2250 8988
rect 1910 8846 1984 8902
rect 2040 8846 2126 8902
rect 2182 8846 2250 8902
rect 1910 8760 2250 8846
rect 1910 8704 1984 8760
rect 2040 8704 2126 8760
rect 2182 8704 2250 8760
rect 1910 8618 2250 8704
rect 1910 8562 1984 8618
rect 2040 8562 2126 8618
rect 2182 8562 2250 8618
rect 1910 8476 2250 8562
rect 1910 8420 1984 8476
rect 2040 8420 2126 8476
rect 2182 8420 2250 8476
rect 1910 8334 2250 8420
rect 1910 8278 1984 8334
rect 2040 8278 2126 8334
rect 2182 8278 2250 8334
rect 1910 8192 2250 8278
rect 1910 8136 1984 8192
rect 2040 8136 2126 8192
rect 2182 8136 2250 8192
rect 1910 8050 2250 8136
rect 1910 7994 1984 8050
rect 2040 7994 2126 8050
rect 2182 7994 2250 8050
rect 1910 7908 2250 7994
rect 1910 7852 1984 7908
rect 2040 7852 2126 7908
rect 2182 7852 2250 7908
rect 1910 7766 2250 7852
rect 1910 7710 1984 7766
rect 2040 7710 2126 7766
rect 2182 7710 2250 7766
rect 1910 7624 2250 7710
rect 1910 7568 1984 7624
rect 2040 7568 2126 7624
rect 2182 7568 2250 7624
rect 1910 7482 2250 7568
rect 1910 7426 1984 7482
rect 2040 7426 2126 7482
rect 2182 7426 2250 7482
rect 1910 7340 2250 7426
rect 1910 7284 1984 7340
rect 2040 7284 2126 7340
rect 2182 7284 2250 7340
rect 1910 7198 2250 7284
rect 1910 7142 1984 7198
rect 2040 7142 2126 7198
rect 2182 7142 2250 7198
rect 1910 7056 2250 7142
rect 1910 7000 1984 7056
rect 2040 7000 2126 7056
rect 2182 7000 2250 7056
rect 1910 6914 2250 7000
rect 1910 6858 1984 6914
rect 2040 6858 2126 6914
rect 2182 6858 2250 6914
rect 1910 6772 2250 6858
rect 1910 6716 1984 6772
rect 2040 6716 2126 6772
rect 2182 6716 2250 6772
rect 1910 6630 2250 6716
rect 1910 6574 1984 6630
rect 2040 6574 2126 6630
rect 2182 6574 2250 6630
rect 1910 6488 2250 6574
rect 1910 6432 1984 6488
rect 2040 6432 2126 6488
rect 2182 6432 2250 6488
rect 1910 6346 2250 6432
rect 1910 6290 1984 6346
rect 2040 6290 2126 6346
rect 2182 6290 2250 6346
rect 1910 6204 2250 6290
rect 1910 6148 1984 6204
rect 2040 6148 2126 6204
rect 2182 6148 2250 6204
rect 1910 6062 2250 6148
rect 1910 6006 1984 6062
rect 2040 6006 2126 6062
rect 2182 6006 2250 6062
rect 1910 5920 2250 6006
rect 1910 5864 1984 5920
rect 2040 5864 2126 5920
rect 2182 5864 2250 5920
rect 1910 5778 2250 5864
rect 1910 5722 1984 5778
rect 2040 5722 2126 5778
rect 2182 5722 2250 5778
rect 1910 5636 2250 5722
rect 1910 5580 1984 5636
rect 2040 5580 2126 5636
rect 2182 5580 2250 5636
rect 1910 5494 2250 5580
rect 1910 5438 1984 5494
rect 2040 5438 2126 5494
rect 2182 5438 2250 5494
rect 1910 5352 2250 5438
rect 1910 5296 1984 5352
rect 2040 5296 2126 5352
rect 2182 5296 2250 5352
rect 1910 5210 2250 5296
rect 1910 5154 1984 5210
rect 2040 5154 2126 5210
rect 2182 5154 2250 5210
rect 1910 5068 2250 5154
rect 1910 5012 1984 5068
rect 2040 5012 2126 5068
rect 2182 5012 2250 5068
rect 1910 4926 2250 5012
rect 1910 4870 1984 4926
rect 2040 4870 2126 4926
rect 2182 4870 2250 4926
rect 1910 4784 2250 4870
rect 1910 4728 1984 4784
rect 2040 4728 2126 4784
rect 2182 4728 2250 4784
rect 1910 4642 2250 4728
rect 1910 4586 1984 4642
rect 2040 4586 2126 4642
rect 2182 4586 2250 4642
rect 1910 4500 2250 4586
rect 1910 4444 1984 4500
rect 2040 4444 2126 4500
rect 2182 4444 2250 4500
rect 1910 4358 2250 4444
rect 1910 4302 1984 4358
rect 2040 4302 2126 4358
rect 2182 4302 2250 4358
rect 1910 4216 2250 4302
rect 1910 4160 1984 4216
rect 2040 4160 2126 4216
rect 2182 4160 2250 4216
rect 1910 4074 2250 4160
rect 1910 4018 1984 4074
rect 2040 4018 2126 4074
rect 2182 4018 2250 4074
rect 1910 3932 2250 4018
rect 1910 3876 1984 3932
rect 2040 3876 2126 3932
rect 2182 3876 2250 3932
rect 1910 3790 2250 3876
rect 1910 3734 1984 3790
rect 2040 3734 2126 3790
rect 2182 3734 2250 3790
rect 1910 3648 2250 3734
rect 1910 3592 1984 3648
rect 2040 3592 2126 3648
rect 2182 3592 2250 3648
rect 1910 3506 2250 3592
rect 1910 3450 1984 3506
rect 2040 3450 2126 3506
rect 2182 3450 2250 3506
rect 1910 3364 2250 3450
rect 1910 3308 1984 3364
rect 2040 3308 2126 3364
rect 2182 3308 2250 3364
rect 1910 3222 2250 3308
rect 1910 3166 1984 3222
rect 2040 3166 2126 3222
rect 2182 3166 2250 3222
rect 1910 3080 2250 3166
rect 1910 3024 1984 3080
rect 2040 3024 2126 3080
rect 2182 3024 2250 3080
rect 1910 2938 2250 3024
rect 1910 2882 1984 2938
rect 2040 2882 2126 2938
rect 2182 2882 2250 2938
rect 1910 2796 2250 2882
rect 1910 2740 1984 2796
rect 2040 2740 2126 2796
rect 2182 2740 2250 2796
rect 1910 2654 2250 2740
rect 1910 2598 1984 2654
rect 2040 2598 2126 2654
rect 2182 2598 2250 2654
rect 1910 2512 2250 2598
rect 1910 2456 1984 2512
rect 2040 2456 2126 2512
rect 2182 2456 2250 2512
rect 1910 2370 2250 2456
rect 1910 2314 1984 2370
rect 2040 2314 2126 2370
rect 2182 2314 2250 2370
rect 1910 2228 2250 2314
rect 1910 2172 1984 2228
rect 2040 2172 2126 2228
rect 2182 2172 2250 2228
rect 1910 2086 2250 2172
rect 1910 2030 1984 2086
rect 2040 2030 2126 2086
rect 2182 2030 2250 2086
rect 1910 1944 2250 2030
rect 1910 1888 1984 1944
rect 2040 1888 2126 1944
rect 2182 1888 2250 1944
rect 1910 1802 2250 1888
rect 1910 1746 1984 1802
rect 2040 1746 2126 1802
rect 2182 1746 2250 1802
rect 1910 1660 2250 1746
rect 1910 1604 1984 1660
rect 2040 1604 2126 1660
rect 2182 1604 2250 1660
rect 1910 1518 2250 1604
rect 1910 1462 1984 1518
rect 2040 1462 2126 1518
rect 2182 1462 2250 1518
rect 1910 1376 2250 1462
rect 1910 1320 1984 1376
rect 2040 1320 2126 1376
rect 2182 1320 2250 1376
rect 1910 1234 2250 1320
rect 1910 1178 1984 1234
rect 2040 1178 2126 1234
rect 2182 1178 2250 1234
rect 1910 1092 2250 1178
rect 1910 1036 1984 1092
rect 2040 1036 2126 1092
rect 2182 1036 2250 1092
rect 1910 950 2250 1036
rect 1910 894 1984 950
rect 2040 894 2126 950
rect 2182 894 2250 950
rect 1910 808 2250 894
rect 1910 752 1984 808
rect 2040 752 2126 808
rect 2182 752 2250 808
rect 1910 666 2250 752
rect 1910 610 1984 666
rect 2040 610 2126 666
rect 2182 610 2250 666
rect 1910 524 2250 610
rect 1910 468 1984 524
rect 2040 468 2126 524
rect 2182 468 2250 524
rect 1910 458 2250 468
rect 2450 12310 2790 12320
rect 2450 12254 2521 12310
rect 2577 12254 2663 12310
rect 2719 12254 2790 12310
rect 2450 12168 2790 12254
rect 2450 12112 2521 12168
rect 2577 12112 2663 12168
rect 2719 12112 2790 12168
rect 2450 12026 2790 12112
rect 2450 11970 2521 12026
rect 2577 11970 2663 12026
rect 2719 11970 2790 12026
rect 2450 11884 2790 11970
rect 2450 11828 2521 11884
rect 2577 11828 2663 11884
rect 2719 11828 2790 11884
rect 2450 11742 2790 11828
rect 2450 11686 2521 11742
rect 2577 11686 2663 11742
rect 2719 11686 2790 11742
rect 2450 11600 2790 11686
rect 2450 11544 2521 11600
rect 2577 11544 2663 11600
rect 2719 11544 2790 11600
rect 2450 11458 2790 11544
rect 2450 11402 2521 11458
rect 2577 11402 2663 11458
rect 2719 11402 2790 11458
rect 2450 11316 2790 11402
rect 2450 11260 2521 11316
rect 2577 11260 2663 11316
rect 2719 11260 2790 11316
rect 2450 11174 2790 11260
rect 2450 11118 2521 11174
rect 2577 11118 2663 11174
rect 2719 11118 2790 11174
rect 2450 11032 2790 11118
rect 2450 10976 2521 11032
rect 2577 10976 2663 11032
rect 2719 10976 2790 11032
rect 2450 10890 2790 10976
rect 2450 10834 2521 10890
rect 2577 10834 2663 10890
rect 2719 10834 2790 10890
rect 2450 10748 2790 10834
rect 2450 10692 2521 10748
rect 2577 10692 2663 10748
rect 2719 10692 2790 10748
rect 2450 10606 2790 10692
rect 2450 10550 2521 10606
rect 2577 10550 2663 10606
rect 2719 10550 2790 10606
rect 2450 10464 2790 10550
rect 2450 10408 2521 10464
rect 2577 10408 2663 10464
rect 2719 10408 2790 10464
rect 2450 10322 2790 10408
rect 2450 10266 2521 10322
rect 2577 10266 2663 10322
rect 2719 10266 2790 10322
rect 2450 10180 2790 10266
rect 2450 10124 2521 10180
rect 2577 10124 2663 10180
rect 2719 10124 2790 10180
rect 2450 10038 2790 10124
rect 2450 9982 2521 10038
rect 2577 9982 2663 10038
rect 2719 9982 2790 10038
rect 2450 9896 2790 9982
rect 2450 9840 2521 9896
rect 2577 9840 2663 9896
rect 2719 9840 2790 9896
rect 2450 9754 2790 9840
rect 2450 9698 2521 9754
rect 2577 9698 2663 9754
rect 2719 9698 2790 9754
rect 2450 9612 2790 9698
rect 2450 9556 2521 9612
rect 2577 9556 2663 9612
rect 2719 9556 2790 9612
rect 2450 9470 2790 9556
rect 2450 9414 2521 9470
rect 2577 9414 2663 9470
rect 2719 9414 2790 9470
rect 2450 9328 2790 9414
rect 2450 9272 2521 9328
rect 2577 9272 2663 9328
rect 2719 9272 2790 9328
rect 2450 9186 2790 9272
rect 2450 9130 2521 9186
rect 2577 9130 2663 9186
rect 2719 9130 2790 9186
rect 2450 9044 2790 9130
rect 2450 8988 2521 9044
rect 2577 8988 2663 9044
rect 2719 8988 2790 9044
rect 2450 8902 2790 8988
rect 2450 8846 2521 8902
rect 2577 8846 2663 8902
rect 2719 8846 2790 8902
rect 2450 8760 2790 8846
rect 2450 8704 2521 8760
rect 2577 8704 2663 8760
rect 2719 8704 2790 8760
rect 2450 8618 2790 8704
rect 2450 8562 2521 8618
rect 2577 8562 2663 8618
rect 2719 8562 2790 8618
rect 2450 8476 2790 8562
rect 2450 8420 2521 8476
rect 2577 8420 2663 8476
rect 2719 8420 2790 8476
rect 2450 8334 2790 8420
rect 2450 8278 2521 8334
rect 2577 8278 2663 8334
rect 2719 8278 2790 8334
rect 2450 8192 2790 8278
rect 2450 8136 2521 8192
rect 2577 8136 2663 8192
rect 2719 8136 2790 8192
rect 2450 8050 2790 8136
rect 2450 7994 2521 8050
rect 2577 7994 2663 8050
rect 2719 7994 2790 8050
rect 2450 7908 2790 7994
rect 2450 7852 2521 7908
rect 2577 7852 2663 7908
rect 2719 7852 2790 7908
rect 2450 7766 2790 7852
rect 2450 7710 2521 7766
rect 2577 7710 2663 7766
rect 2719 7710 2790 7766
rect 2450 7624 2790 7710
rect 2450 7568 2521 7624
rect 2577 7568 2663 7624
rect 2719 7568 2790 7624
rect 2450 7482 2790 7568
rect 2450 7426 2521 7482
rect 2577 7426 2663 7482
rect 2719 7426 2790 7482
rect 2450 7340 2790 7426
rect 2450 7284 2521 7340
rect 2577 7284 2663 7340
rect 2719 7284 2790 7340
rect 2450 7198 2790 7284
rect 2450 7142 2521 7198
rect 2577 7142 2663 7198
rect 2719 7142 2790 7198
rect 2450 7056 2790 7142
rect 2450 7000 2521 7056
rect 2577 7000 2663 7056
rect 2719 7000 2790 7056
rect 2450 6914 2790 7000
rect 2450 6858 2521 6914
rect 2577 6858 2663 6914
rect 2719 6858 2790 6914
rect 2450 6772 2790 6858
rect 2450 6716 2521 6772
rect 2577 6716 2663 6772
rect 2719 6716 2790 6772
rect 2450 6630 2790 6716
rect 2450 6574 2521 6630
rect 2577 6574 2663 6630
rect 2719 6574 2790 6630
rect 2450 6488 2790 6574
rect 2450 6432 2521 6488
rect 2577 6432 2663 6488
rect 2719 6432 2790 6488
rect 2450 6346 2790 6432
rect 2450 6290 2521 6346
rect 2577 6290 2663 6346
rect 2719 6290 2790 6346
rect 2450 6204 2790 6290
rect 2450 6148 2521 6204
rect 2577 6148 2663 6204
rect 2719 6148 2790 6204
rect 2450 6062 2790 6148
rect 2450 6006 2521 6062
rect 2577 6006 2663 6062
rect 2719 6006 2790 6062
rect 2450 5920 2790 6006
rect 2450 5864 2521 5920
rect 2577 5864 2663 5920
rect 2719 5864 2790 5920
rect 2450 5778 2790 5864
rect 2450 5722 2521 5778
rect 2577 5722 2663 5778
rect 2719 5722 2790 5778
rect 2450 5636 2790 5722
rect 2450 5580 2521 5636
rect 2577 5580 2663 5636
rect 2719 5580 2790 5636
rect 2450 5494 2790 5580
rect 2450 5438 2521 5494
rect 2577 5438 2663 5494
rect 2719 5438 2790 5494
rect 2450 5352 2790 5438
rect 2450 5296 2521 5352
rect 2577 5296 2663 5352
rect 2719 5296 2790 5352
rect 2450 5210 2790 5296
rect 2450 5154 2521 5210
rect 2577 5154 2663 5210
rect 2719 5154 2790 5210
rect 2450 5068 2790 5154
rect 2450 5012 2521 5068
rect 2577 5012 2663 5068
rect 2719 5012 2790 5068
rect 2450 4926 2790 5012
rect 2450 4870 2521 4926
rect 2577 4870 2663 4926
rect 2719 4870 2790 4926
rect 2450 4784 2790 4870
rect 2450 4728 2521 4784
rect 2577 4728 2663 4784
rect 2719 4728 2790 4784
rect 2450 4642 2790 4728
rect 2450 4586 2521 4642
rect 2577 4586 2663 4642
rect 2719 4586 2790 4642
rect 2450 4500 2790 4586
rect 2450 4444 2521 4500
rect 2577 4444 2663 4500
rect 2719 4444 2790 4500
rect 2450 4358 2790 4444
rect 2450 4302 2521 4358
rect 2577 4302 2663 4358
rect 2719 4302 2790 4358
rect 2450 4216 2790 4302
rect 2450 4160 2521 4216
rect 2577 4160 2663 4216
rect 2719 4160 2790 4216
rect 2450 4074 2790 4160
rect 2450 4018 2521 4074
rect 2577 4018 2663 4074
rect 2719 4018 2790 4074
rect 2450 3932 2790 4018
rect 2450 3876 2521 3932
rect 2577 3876 2663 3932
rect 2719 3876 2790 3932
rect 2450 3790 2790 3876
rect 2450 3734 2521 3790
rect 2577 3734 2663 3790
rect 2719 3734 2790 3790
rect 2450 3648 2790 3734
rect 2450 3592 2521 3648
rect 2577 3592 2663 3648
rect 2719 3592 2790 3648
rect 2450 3506 2790 3592
rect 2450 3450 2521 3506
rect 2577 3450 2663 3506
rect 2719 3450 2790 3506
rect 2450 3364 2790 3450
rect 2450 3308 2521 3364
rect 2577 3308 2663 3364
rect 2719 3308 2790 3364
rect 2450 3222 2790 3308
rect 2450 3166 2521 3222
rect 2577 3166 2663 3222
rect 2719 3166 2790 3222
rect 2450 3080 2790 3166
rect 2450 3024 2521 3080
rect 2577 3024 2663 3080
rect 2719 3024 2790 3080
rect 2450 2938 2790 3024
rect 2450 2882 2521 2938
rect 2577 2882 2663 2938
rect 2719 2882 2790 2938
rect 2450 2796 2790 2882
rect 2450 2740 2521 2796
rect 2577 2740 2663 2796
rect 2719 2740 2790 2796
rect 2450 2654 2790 2740
rect 2450 2598 2521 2654
rect 2577 2598 2663 2654
rect 2719 2598 2790 2654
rect 2450 2512 2790 2598
rect 2450 2456 2521 2512
rect 2577 2456 2663 2512
rect 2719 2456 2790 2512
rect 2450 2370 2790 2456
rect 2450 2314 2521 2370
rect 2577 2314 2663 2370
rect 2719 2314 2790 2370
rect 2450 2228 2790 2314
rect 2450 2172 2521 2228
rect 2577 2172 2663 2228
rect 2719 2172 2790 2228
rect 2450 2086 2790 2172
rect 2450 2030 2521 2086
rect 2577 2030 2663 2086
rect 2719 2030 2790 2086
rect 2450 1944 2790 2030
rect 2450 1888 2521 1944
rect 2577 1888 2663 1944
rect 2719 1888 2790 1944
rect 2450 1802 2790 1888
rect 2450 1746 2521 1802
rect 2577 1746 2663 1802
rect 2719 1746 2790 1802
rect 2450 1660 2790 1746
rect 2450 1604 2521 1660
rect 2577 1604 2663 1660
rect 2719 1604 2790 1660
rect 2450 1518 2790 1604
rect 2450 1462 2521 1518
rect 2577 1462 2663 1518
rect 2719 1462 2790 1518
rect 2450 1376 2790 1462
rect 2450 1320 2521 1376
rect 2577 1320 2663 1376
rect 2719 1320 2790 1376
rect 2450 1234 2790 1320
rect 2450 1178 2521 1234
rect 2577 1178 2663 1234
rect 2719 1178 2790 1234
rect 2450 1092 2790 1178
rect 2450 1036 2521 1092
rect 2577 1036 2663 1092
rect 2719 1036 2790 1092
rect 2450 950 2790 1036
rect 2450 894 2521 950
rect 2577 894 2663 950
rect 2719 894 2790 950
rect 2450 808 2790 894
rect 2450 752 2521 808
rect 2577 752 2663 808
rect 2719 752 2790 808
rect 2450 666 2790 752
rect 2450 610 2521 666
rect 2577 610 2663 666
rect 2719 610 2790 666
rect 2450 524 2790 610
rect 2450 468 2521 524
rect 2577 468 2663 524
rect 2719 468 2790 524
rect 2450 458 2790 468
rect 2990 12310 3330 12320
rect 2990 12254 3058 12310
rect 3114 12254 3200 12310
rect 3256 12254 3330 12310
rect 2990 12168 3330 12254
rect 2990 12112 3058 12168
rect 3114 12112 3200 12168
rect 3256 12112 3330 12168
rect 2990 12026 3330 12112
rect 2990 11970 3058 12026
rect 3114 11970 3200 12026
rect 3256 11970 3330 12026
rect 2990 11884 3330 11970
rect 2990 11828 3058 11884
rect 3114 11828 3200 11884
rect 3256 11828 3330 11884
rect 2990 11742 3330 11828
rect 2990 11686 3058 11742
rect 3114 11686 3200 11742
rect 3256 11686 3330 11742
rect 2990 11600 3330 11686
rect 2990 11544 3058 11600
rect 3114 11544 3200 11600
rect 3256 11544 3330 11600
rect 2990 11458 3330 11544
rect 2990 11402 3058 11458
rect 3114 11402 3200 11458
rect 3256 11402 3330 11458
rect 2990 11316 3330 11402
rect 2990 11260 3058 11316
rect 3114 11260 3200 11316
rect 3256 11260 3330 11316
rect 2990 11174 3330 11260
rect 2990 11118 3058 11174
rect 3114 11118 3200 11174
rect 3256 11118 3330 11174
rect 2990 11032 3330 11118
rect 2990 10976 3058 11032
rect 3114 10976 3200 11032
rect 3256 10976 3330 11032
rect 2990 10890 3330 10976
rect 2990 10834 3058 10890
rect 3114 10834 3200 10890
rect 3256 10834 3330 10890
rect 2990 10748 3330 10834
rect 2990 10692 3058 10748
rect 3114 10692 3200 10748
rect 3256 10692 3330 10748
rect 2990 10606 3330 10692
rect 2990 10550 3058 10606
rect 3114 10550 3200 10606
rect 3256 10550 3330 10606
rect 2990 10464 3330 10550
rect 2990 10408 3058 10464
rect 3114 10408 3200 10464
rect 3256 10408 3330 10464
rect 2990 10322 3330 10408
rect 2990 10266 3058 10322
rect 3114 10266 3200 10322
rect 3256 10266 3330 10322
rect 2990 10180 3330 10266
rect 2990 10124 3058 10180
rect 3114 10124 3200 10180
rect 3256 10124 3330 10180
rect 2990 10038 3330 10124
rect 2990 9982 3058 10038
rect 3114 9982 3200 10038
rect 3256 9982 3330 10038
rect 2990 9896 3330 9982
rect 2990 9840 3058 9896
rect 3114 9840 3200 9896
rect 3256 9840 3330 9896
rect 2990 9754 3330 9840
rect 2990 9698 3058 9754
rect 3114 9698 3200 9754
rect 3256 9698 3330 9754
rect 2990 9612 3330 9698
rect 2990 9556 3058 9612
rect 3114 9556 3200 9612
rect 3256 9556 3330 9612
rect 2990 9470 3330 9556
rect 2990 9414 3058 9470
rect 3114 9414 3200 9470
rect 3256 9414 3330 9470
rect 2990 9328 3330 9414
rect 2990 9272 3058 9328
rect 3114 9272 3200 9328
rect 3256 9272 3330 9328
rect 2990 9186 3330 9272
rect 2990 9130 3058 9186
rect 3114 9130 3200 9186
rect 3256 9130 3330 9186
rect 2990 9044 3330 9130
rect 2990 8988 3058 9044
rect 3114 8988 3200 9044
rect 3256 8988 3330 9044
rect 2990 8902 3330 8988
rect 2990 8846 3058 8902
rect 3114 8846 3200 8902
rect 3256 8846 3330 8902
rect 2990 8760 3330 8846
rect 2990 8704 3058 8760
rect 3114 8704 3200 8760
rect 3256 8704 3330 8760
rect 2990 8618 3330 8704
rect 2990 8562 3058 8618
rect 3114 8562 3200 8618
rect 3256 8562 3330 8618
rect 2990 8476 3330 8562
rect 2990 8420 3058 8476
rect 3114 8420 3200 8476
rect 3256 8420 3330 8476
rect 2990 8334 3330 8420
rect 2990 8278 3058 8334
rect 3114 8278 3200 8334
rect 3256 8278 3330 8334
rect 2990 8192 3330 8278
rect 2990 8136 3058 8192
rect 3114 8136 3200 8192
rect 3256 8136 3330 8192
rect 2990 8050 3330 8136
rect 2990 7994 3058 8050
rect 3114 7994 3200 8050
rect 3256 7994 3330 8050
rect 2990 7908 3330 7994
rect 2990 7852 3058 7908
rect 3114 7852 3200 7908
rect 3256 7852 3330 7908
rect 2990 7766 3330 7852
rect 2990 7710 3058 7766
rect 3114 7710 3200 7766
rect 3256 7710 3330 7766
rect 2990 7624 3330 7710
rect 2990 7568 3058 7624
rect 3114 7568 3200 7624
rect 3256 7568 3330 7624
rect 2990 7482 3330 7568
rect 2990 7426 3058 7482
rect 3114 7426 3200 7482
rect 3256 7426 3330 7482
rect 2990 7340 3330 7426
rect 2990 7284 3058 7340
rect 3114 7284 3200 7340
rect 3256 7284 3330 7340
rect 2990 7198 3330 7284
rect 2990 7142 3058 7198
rect 3114 7142 3200 7198
rect 3256 7142 3330 7198
rect 2990 7056 3330 7142
rect 2990 7000 3058 7056
rect 3114 7000 3200 7056
rect 3256 7000 3330 7056
rect 2990 6914 3330 7000
rect 2990 6858 3058 6914
rect 3114 6858 3200 6914
rect 3256 6858 3330 6914
rect 2990 6772 3330 6858
rect 2990 6716 3058 6772
rect 3114 6716 3200 6772
rect 3256 6716 3330 6772
rect 2990 6630 3330 6716
rect 2990 6574 3058 6630
rect 3114 6574 3200 6630
rect 3256 6574 3330 6630
rect 2990 6488 3330 6574
rect 2990 6432 3058 6488
rect 3114 6432 3200 6488
rect 3256 6432 3330 6488
rect 2990 6346 3330 6432
rect 2990 6290 3058 6346
rect 3114 6290 3200 6346
rect 3256 6290 3330 6346
rect 2990 6204 3330 6290
rect 2990 6148 3058 6204
rect 3114 6148 3200 6204
rect 3256 6148 3330 6204
rect 2990 6062 3330 6148
rect 2990 6006 3058 6062
rect 3114 6006 3200 6062
rect 3256 6006 3330 6062
rect 2990 5920 3330 6006
rect 2990 5864 3058 5920
rect 3114 5864 3200 5920
rect 3256 5864 3330 5920
rect 2990 5778 3330 5864
rect 2990 5722 3058 5778
rect 3114 5722 3200 5778
rect 3256 5722 3330 5778
rect 2990 5636 3330 5722
rect 2990 5580 3058 5636
rect 3114 5580 3200 5636
rect 3256 5580 3330 5636
rect 2990 5494 3330 5580
rect 2990 5438 3058 5494
rect 3114 5438 3200 5494
rect 3256 5438 3330 5494
rect 2990 5352 3330 5438
rect 2990 5296 3058 5352
rect 3114 5296 3200 5352
rect 3256 5296 3330 5352
rect 2990 5210 3330 5296
rect 2990 5154 3058 5210
rect 3114 5154 3200 5210
rect 3256 5154 3330 5210
rect 2990 5068 3330 5154
rect 2990 5012 3058 5068
rect 3114 5012 3200 5068
rect 3256 5012 3330 5068
rect 2990 4926 3330 5012
rect 2990 4870 3058 4926
rect 3114 4870 3200 4926
rect 3256 4870 3330 4926
rect 2990 4784 3330 4870
rect 2990 4728 3058 4784
rect 3114 4728 3200 4784
rect 3256 4728 3330 4784
rect 2990 4642 3330 4728
rect 2990 4586 3058 4642
rect 3114 4586 3200 4642
rect 3256 4586 3330 4642
rect 2990 4500 3330 4586
rect 2990 4444 3058 4500
rect 3114 4444 3200 4500
rect 3256 4444 3330 4500
rect 2990 4358 3330 4444
rect 2990 4302 3058 4358
rect 3114 4302 3200 4358
rect 3256 4302 3330 4358
rect 2990 4216 3330 4302
rect 2990 4160 3058 4216
rect 3114 4160 3200 4216
rect 3256 4160 3330 4216
rect 2990 4074 3330 4160
rect 2990 4018 3058 4074
rect 3114 4018 3200 4074
rect 3256 4018 3330 4074
rect 2990 3932 3330 4018
rect 2990 3876 3058 3932
rect 3114 3876 3200 3932
rect 3256 3876 3330 3932
rect 2990 3790 3330 3876
rect 2990 3734 3058 3790
rect 3114 3734 3200 3790
rect 3256 3734 3330 3790
rect 2990 3648 3330 3734
rect 2990 3592 3058 3648
rect 3114 3592 3200 3648
rect 3256 3592 3330 3648
rect 2990 3506 3330 3592
rect 2990 3450 3058 3506
rect 3114 3450 3200 3506
rect 3256 3450 3330 3506
rect 2990 3364 3330 3450
rect 2990 3308 3058 3364
rect 3114 3308 3200 3364
rect 3256 3308 3330 3364
rect 2990 3222 3330 3308
rect 2990 3166 3058 3222
rect 3114 3166 3200 3222
rect 3256 3166 3330 3222
rect 2990 3080 3330 3166
rect 2990 3024 3058 3080
rect 3114 3024 3200 3080
rect 3256 3024 3330 3080
rect 2990 2938 3330 3024
rect 2990 2882 3058 2938
rect 3114 2882 3200 2938
rect 3256 2882 3330 2938
rect 2990 2796 3330 2882
rect 2990 2740 3058 2796
rect 3114 2740 3200 2796
rect 3256 2740 3330 2796
rect 2990 2654 3330 2740
rect 2990 2598 3058 2654
rect 3114 2598 3200 2654
rect 3256 2598 3330 2654
rect 2990 2512 3330 2598
rect 2990 2456 3058 2512
rect 3114 2456 3200 2512
rect 3256 2456 3330 2512
rect 2990 2370 3330 2456
rect 2990 2314 3058 2370
rect 3114 2314 3200 2370
rect 3256 2314 3330 2370
rect 2990 2228 3330 2314
rect 2990 2172 3058 2228
rect 3114 2172 3200 2228
rect 3256 2172 3330 2228
rect 2990 2086 3330 2172
rect 2990 2030 3058 2086
rect 3114 2030 3200 2086
rect 3256 2030 3330 2086
rect 2990 1944 3330 2030
rect 2990 1888 3058 1944
rect 3114 1888 3200 1944
rect 3256 1888 3330 1944
rect 2990 1802 3330 1888
rect 2990 1746 3058 1802
rect 3114 1746 3200 1802
rect 3256 1746 3330 1802
rect 2990 1660 3330 1746
rect 2990 1604 3058 1660
rect 3114 1604 3200 1660
rect 3256 1604 3330 1660
rect 2990 1518 3330 1604
rect 2990 1462 3058 1518
rect 3114 1462 3200 1518
rect 3256 1462 3330 1518
rect 2990 1376 3330 1462
rect 2990 1320 3058 1376
rect 3114 1320 3200 1376
rect 3256 1320 3330 1376
rect 2990 1234 3330 1320
rect 2990 1178 3058 1234
rect 3114 1178 3200 1234
rect 3256 1178 3330 1234
rect 2990 1092 3330 1178
rect 2990 1036 3058 1092
rect 3114 1036 3200 1092
rect 3256 1036 3330 1092
rect 2990 950 3330 1036
rect 2990 894 3058 950
rect 3114 894 3200 950
rect 3256 894 3330 950
rect 2990 808 3330 894
rect 2990 752 3058 808
rect 3114 752 3200 808
rect 3256 752 3330 808
rect 2990 666 3330 752
rect 2990 610 3058 666
rect 3114 610 3200 666
rect 3256 610 3330 666
rect 2990 524 3330 610
rect 2990 468 3058 524
rect 3114 468 3200 524
rect 3256 468 3330 524
rect 2990 458 3330 468
rect 3530 12310 3870 12320
rect 3530 12254 3602 12310
rect 3658 12254 3744 12310
rect 3800 12254 3870 12310
rect 3530 12168 3870 12254
rect 3530 12112 3602 12168
rect 3658 12112 3744 12168
rect 3800 12112 3870 12168
rect 3530 12026 3870 12112
rect 3530 11970 3602 12026
rect 3658 11970 3744 12026
rect 3800 11970 3870 12026
rect 3530 11884 3870 11970
rect 3530 11828 3602 11884
rect 3658 11828 3744 11884
rect 3800 11828 3870 11884
rect 3530 11742 3870 11828
rect 3530 11686 3602 11742
rect 3658 11686 3744 11742
rect 3800 11686 3870 11742
rect 3530 11600 3870 11686
rect 3530 11544 3602 11600
rect 3658 11544 3744 11600
rect 3800 11544 3870 11600
rect 3530 11458 3870 11544
rect 3530 11402 3602 11458
rect 3658 11402 3744 11458
rect 3800 11402 3870 11458
rect 3530 11316 3870 11402
rect 3530 11260 3602 11316
rect 3658 11260 3744 11316
rect 3800 11260 3870 11316
rect 3530 11174 3870 11260
rect 3530 11118 3602 11174
rect 3658 11118 3744 11174
rect 3800 11118 3870 11174
rect 3530 11032 3870 11118
rect 3530 10976 3602 11032
rect 3658 10976 3744 11032
rect 3800 10976 3870 11032
rect 3530 10890 3870 10976
rect 3530 10834 3602 10890
rect 3658 10834 3744 10890
rect 3800 10834 3870 10890
rect 3530 10748 3870 10834
rect 3530 10692 3602 10748
rect 3658 10692 3744 10748
rect 3800 10692 3870 10748
rect 3530 10606 3870 10692
rect 3530 10550 3602 10606
rect 3658 10550 3744 10606
rect 3800 10550 3870 10606
rect 3530 10464 3870 10550
rect 3530 10408 3602 10464
rect 3658 10408 3744 10464
rect 3800 10408 3870 10464
rect 3530 10322 3870 10408
rect 3530 10266 3602 10322
rect 3658 10266 3744 10322
rect 3800 10266 3870 10322
rect 3530 10180 3870 10266
rect 3530 10124 3602 10180
rect 3658 10124 3744 10180
rect 3800 10124 3870 10180
rect 3530 10038 3870 10124
rect 3530 9982 3602 10038
rect 3658 9982 3744 10038
rect 3800 9982 3870 10038
rect 3530 9896 3870 9982
rect 3530 9840 3602 9896
rect 3658 9840 3744 9896
rect 3800 9840 3870 9896
rect 3530 9754 3870 9840
rect 3530 9698 3602 9754
rect 3658 9698 3744 9754
rect 3800 9698 3870 9754
rect 3530 9612 3870 9698
rect 3530 9556 3602 9612
rect 3658 9556 3744 9612
rect 3800 9556 3870 9612
rect 3530 9470 3870 9556
rect 3530 9414 3602 9470
rect 3658 9414 3744 9470
rect 3800 9414 3870 9470
rect 3530 9328 3870 9414
rect 3530 9272 3602 9328
rect 3658 9272 3744 9328
rect 3800 9272 3870 9328
rect 3530 9186 3870 9272
rect 3530 9130 3602 9186
rect 3658 9130 3744 9186
rect 3800 9130 3870 9186
rect 3530 9044 3870 9130
rect 3530 8988 3602 9044
rect 3658 8988 3744 9044
rect 3800 8988 3870 9044
rect 3530 8902 3870 8988
rect 3530 8846 3602 8902
rect 3658 8846 3744 8902
rect 3800 8846 3870 8902
rect 3530 8760 3870 8846
rect 3530 8704 3602 8760
rect 3658 8704 3744 8760
rect 3800 8704 3870 8760
rect 3530 8618 3870 8704
rect 3530 8562 3602 8618
rect 3658 8562 3744 8618
rect 3800 8562 3870 8618
rect 3530 8476 3870 8562
rect 3530 8420 3602 8476
rect 3658 8420 3744 8476
rect 3800 8420 3870 8476
rect 3530 8334 3870 8420
rect 3530 8278 3602 8334
rect 3658 8278 3744 8334
rect 3800 8278 3870 8334
rect 3530 8192 3870 8278
rect 3530 8136 3602 8192
rect 3658 8136 3744 8192
rect 3800 8136 3870 8192
rect 3530 8050 3870 8136
rect 3530 7994 3602 8050
rect 3658 7994 3744 8050
rect 3800 7994 3870 8050
rect 3530 7908 3870 7994
rect 3530 7852 3602 7908
rect 3658 7852 3744 7908
rect 3800 7852 3870 7908
rect 3530 7766 3870 7852
rect 3530 7710 3602 7766
rect 3658 7710 3744 7766
rect 3800 7710 3870 7766
rect 3530 7624 3870 7710
rect 3530 7568 3602 7624
rect 3658 7568 3744 7624
rect 3800 7568 3870 7624
rect 3530 7482 3870 7568
rect 3530 7426 3602 7482
rect 3658 7426 3744 7482
rect 3800 7426 3870 7482
rect 3530 7340 3870 7426
rect 3530 7284 3602 7340
rect 3658 7284 3744 7340
rect 3800 7284 3870 7340
rect 3530 7198 3870 7284
rect 3530 7142 3602 7198
rect 3658 7142 3744 7198
rect 3800 7142 3870 7198
rect 3530 7056 3870 7142
rect 3530 7000 3602 7056
rect 3658 7000 3744 7056
rect 3800 7000 3870 7056
rect 3530 6914 3870 7000
rect 3530 6858 3602 6914
rect 3658 6858 3744 6914
rect 3800 6858 3870 6914
rect 3530 6772 3870 6858
rect 3530 6716 3602 6772
rect 3658 6716 3744 6772
rect 3800 6716 3870 6772
rect 3530 6630 3870 6716
rect 3530 6574 3602 6630
rect 3658 6574 3744 6630
rect 3800 6574 3870 6630
rect 3530 6488 3870 6574
rect 3530 6432 3602 6488
rect 3658 6432 3744 6488
rect 3800 6432 3870 6488
rect 3530 6346 3870 6432
rect 3530 6290 3602 6346
rect 3658 6290 3744 6346
rect 3800 6290 3870 6346
rect 3530 6204 3870 6290
rect 3530 6148 3602 6204
rect 3658 6148 3744 6204
rect 3800 6148 3870 6204
rect 3530 6062 3870 6148
rect 3530 6006 3602 6062
rect 3658 6006 3744 6062
rect 3800 6006 3870 6062
rect 3530 5920 3870 6006
rect 3530 5864 3602 5920
rect 3658 5864 3744 5920
rect 3800 5864 3870 5920
rect 3530 5778 3870 5864
rect 3530 5722 3602 5778
rect 3658 5722 3744 5778
rect 3800 5722 3870 5778
rect 3530 5636 3870 5722
rect 3530 5580 3602 5636
rect 3658 5580 3744 5636
rect 3800 5580 3870 5636
rect 3530 5494 3870 5580
rect 3530 5438 3602 5494
rect 3658 5438 3744 5494
rect 3800 5438 3870 5494
rect 3530 5352 3870 5438
rect 3530 5296 3602 5352
rect 3658 5296 3744 5352
rect 3800 5296 3870 5352
rect 3530 5210 3870 5296
rect 3530 5154 3602 5210
rect 3658 5154 3744 5210
rect 3800 5154 3870 5210
rect 3530 5068 3870 5154
rect 3530 5012 3602 5068
rect 3658 5012 3744 5068
rect 3800 5012 3870 5068
rect 3530 4926 3870 5012
rect 3530 4870 3602 4926
rect 3658 4870 3744 4926
rect 3800 4870 3870 4926
rect 3530 4784 3870 4870
rect 3530 4728 3602 4784
rect 3658 4728 3744 4784
rect 3800 4728 3870 4784
rect 3530 4642 3870 4728
rect 3530 4586 3602 4642
rect 3658 4586 3744 4642
rect 3800 4586 3870 4642
rect 3530 4500 3870 4586
rect 3530 4444 3602 4500
rect 3658 4444 3744 4500
rect 3800 4444 3870 4500
rect 3530 4358 3870 4444
rect 3530 4302 3602 4358
rect 3658 4302 3744 4358
rect 3800 4302 3870 4358
rect 3530 4216 3870 4302
rect 3530 4160 3602 4216
rect 3658 4160 3744 4216
rect 3800 4160 3870 4216
rect 3530 4074 3870 4160
rect 3530 4018 3602 4074
rect 3658 4018 3744 4074
rect 3800 4018 3870 4074
rect 3530 3932 3870 4018
rect 3530 3876 3602 3932
rect 3658 3876 3744 3932
rect 3800 3876 3870 3932
rect 3530 3790 3870 3876
rect 3530 3734 3602 3790
rect 3658 3734 3744 3790
rect 3800 3734 3870 3790
rect 3530 3648 3870 3734
rect 3530 3592 3602 3648
rect 3658 3592 3744 3648
rect 3800 3592 3870 3648
rect 3530 3506 3870 3592
rect 3530 3450 3602 3506
rect 3658 3450 3744 3506
rect 3800 3450 3870 3506
rect 3530 3364 3870 3450
rect 3530 3308 3602 3364
rect 3658 3308 3744 3364
rect 3800 3308 3870 3364
rect 3530 3222 3870 3308
rect 3530 3166 3602 3222
rect 3658 3166 3744 3222
rect 3800 3166 3870 3222
rect 3530 3080 3870 3166
rect 3530 3024 3602 3080
rect 3658 3024 3744 3080
rect 3800 3024 3870 3080
rect 3530 2938 3870 3024
rect 3530 2882 3602 2938
rect 3658 2882 3744 2938
rect 3800 2882 3870 2938
rect 3530 2796 3870 2882
rect 3530 2740 3602 2796
rect 3658 2740 3744 2796
rect 3800 2740 3870 2796
rect 3530 2654 3870 2740
rect 3530 2598 3602 2654
rect 3658 2598 3744 2654
rect 3800 2598 3870 2654
rect 3530 2512 3870 2598
rect 3530 2456 3602 2512
rect 3658 2456 3744 2512
rect 3800 2456 3870 2512
rect 3530 2370 3870 2456
rect 3530 2314 3602 2370
rect 3658 2314 3744 2370
rect 3800 2314 3870 2370
rect 3530 2228 3870 2314
rect 3530 2172 3602 2228
rect 3658 2172 3744 2228
rect 3800 2172 3870 2228
rect 3530 2086 3870 2172
rect 3530 2030 3602 2086
rect 3658 2030 3744 2086
rect 3800 2030 3870 2086
rect 3530 1944 3870 2030
rect 3530 1888 3602 1944
rect 3658 1888 3744 1944
rect 3800 1888 3870 1944
rect 3530 1802 3870 1888
rect 3530 1746 3602 1802
rect 3658 1746 3744 1802
rect 3800 1746 3870 1802
rect 3530 1660 3870 1746
rect 3530 1604 3602 1660
rect 3658 1604 3744 1660
rect 3800 1604 3870 1660
rect 3530 1518 3870 1604
rect 3530 1462 3602 1518
rect 3658 1462 3744 1518
rect 3800 1462 3870 1518
rect 3530 1376 3870 1462
rect 3530 1320 3602 1376
rect 3658 1320 3744 1376
rect 3800 1320 3870 1376
rect 3530 1234 3870 1320
rect 3530 1178 3602 1234
rect 3658 1178 3744 1234
rect 3800 1178 3870 1234
rect 3530 1092 3870 1178
rect 3530 1036 3602 1092
rect 3658 1036 3744 1092
rect 3800 1036 3870 1092
rect 3530 950 3870 1036
rect 3530 894 3602 950
rect 3658 894 3744 950
rect 3800 894 3870 950
rect 3530 808 3870 894
rect 3530 752 3602 808
rect 3658 752 3744 808
rect 3800 752 3870 808
rect 3530 666 3870 752
rect 3530 610 3602 666
rect 3658 610 3744 666
rect 3800 610 3870 666
rect 3530 524 3870 610
rect 3530 468 3602 524
rect 3658 468 3744 524
rect 3800 468 3870 524
rect 3530 458 3870 468
rect 4070 12310 4410 12320
rect 4070 12254 4138 12310
rect 4194 12254 4280 12310
rect 4336 12254 4410 12310
rect 4070 12168 4410 12254
rect 4070 12112 4138 12168
rect 4194 12112 4280 12168
rect 4336 12112 4410 12168
rect 4070 12026 4410 12112
rect 4070 11970 4138 12026
rect 4194 11970 4280 12026
rect 4336 11970 4410 12026
rect 4070 11884 4410 11970
rect 4070 11828 4138 11884
rect 4194 11828 4280 11884
rect 4336 11828 4410 11884
rect 4070 11742 4410 11828
rect 4070 11686 4138 11742
rect 4194 11686 4280 11742
rect 4336 11686 4410 11742
rect 4070 11600 4410 11686
rect 4070 11544 4138 11600
rect 4194 11544 4280 11600
rect 4336 11544 4410 11600
rect 4070 11458 4410 11544
rect 4070 11402 4138 11458
rect 4194 11402 4280 11458
rect 4336 11402 4410 11458
rect 4070 11316 4410 11402
rect 4070 11260 4138 11316
rect 4194 11260 4280 11316
rect 4336 11260 4410 11316
rect 4070 11174 4410 11260
rect 4070 11118 4138 11174
rect 4194 11118 4280 11174
rect 4336 11118 4410 11174
rect 4070 11032 4410 11118
rect 4070 10976 4138 11032
rect 4194 10976 4280 11032
rect 4336 10976 4410 11032
rect 4070 10890 4410 10976
rect 4070 10834 4138 10890
rect 4194 10834 4280 10890
rect 4336 10834 4410 10890
rect 4070 10748 4410 10834
rect 4070 10692 4138 10748
rect 4194 10692 4280 10748
rect 4336 10692 4410 10748
rect 4070 10606 4410 10692
rect 4070 10550 4138 10606
rect 4194 10550 4280 10606
rect 4336 10550 4410 10606
rect 4070 10464 4410 10550
rect 4070 10408 4138 10464
rect 4194 10408 4280 10464
rect 4336 10408 4410 10464
rect 4070 10322 4410 10408
rect 4070 10266 4138 10322
rect 4194 10266 4280 10322
rect 4336 10266 4410 10322
rect 4070 10180 4410 10266
rect 4070 10124 4138 10180
rect 4194 10124 4280 10180
rect 4336 10124 4410 10180
rect 4070 10038 4410 10124
rect 4070 9982 4138 10038
rect 4194 9982 4280 10038
rect 4336 9982 4410 10038
rect 4070 9896 4410 9982
rect 4070 9840 4138 9896
rect 4194 9840 4280 9896
rect 4336 9840 4410 9896
rect 4070 9754 4410 9840
rect 4070 9698 4138 9754
rect 4194 9698 4280 9754
rect 4336 9698 4410 9754
rect 4070 9612 4410 9698
rect 4070 9556 4138 9612
rect 4194 9556 4280 9612
rect 4336 9556 4410 9612
rect 4070 9470 4410 9556
rect 4070 9414 4138 9470
rect 4194 9414 4280 9470
rect 4336 9414 4410 9470
rect 4070 9328 4410 9414
rect 4070 9272 4138 9328
rect 4194 9272 4280 9328
rect 4336 9272 4410 9328
rect 4070 9186 4410 9272
rect 4070 9130 4138 9186
rect 4194 9130 4280 9186
rect 4336 9130 4410 9186
rect 4070 9044 4410 9130
rect 4070 8988 4138 9044
rect 4194 8988 4280 9044
rect 4336 8988 4410 9044
rect 4070 8902 4410 8988
rect 4070 8846 4138 8902
rect 4194 8846 4280 8902
rect 4336 8846 4410 8902
rect 4070 8760 4410 8846
rect 4070 8704 4138 8760
rect 4194 8704 4280 8760
rect 4336 8704 4410 8760
rect 4070 8618 4410 8704
rect 4070 8562 4138 8618
rect 4194 8562 4280 8618
rect 4336 8562 4410 8618
rect 4070 8476 4410 8562
rect 4070 8420 4138 8476
rect 4194 8420 4280 8476
rect 4336 8420 4410 8476
rect 4070 8334 4410 8420
rect 4070 8278 4138 8334
rect 4194 8278 4280 8334
rect 4336 8278 4410 8334
rect 4070 8192 4410 8278
rect 4070 8136 4138 8192
rect 4194 8136 4280 8192
rect 4336 8136 4410 8192
rect 4070 8050 4410 8136
rect 4070 7994 4138 8050
rect 4194 7994 4280 8050
rect 4336 7994 4410 8050
rect 4070 7908 4410 7994
rect 4070 7852 4138 7908
rect 4194 7852 4280 7908
rect 4336 7852 4410 7908
rect 4070 7766 4410 7852
rect 4070 7710 4138 7766
rect 4194 7710 4280 7766
rect 4336 7710 4410 7766
rect 4070 7624 4410 7710
rect 4070 7568 4138 7624
rect 4194 7568 4280 7624
rect 4336 7568 4410 7624
rect 4070 7482 4410 7568
rect 4070 7426 4138 7482
rect 4194 7426 4280 7482
rect 4336 7426 4410 7482
rect 4070 7340 4410 7426
rect 4070 7284 4138 7340
rect 4194 7284 4280 7340
rect 4336 7284 4410 7340
rect 4070 7198 4410 7284
rect 4070 7142 4138 7198
rect 4194 7142 4280 7198
rect 4336 7142 4410 7198
rect 4070 7056 4410 7142
rect 4070 7000 4138 7056
rect 4194 7000 4280 7056
rect 4336 7000 4410 7056
rect 4070 6914 4410 7000
rect 4070 6858 4138 6914
rect 4194 6858 4280 6914
rect 4336 6858 4410 6914
rect 4070 6772 4410 6858
rect 4070 6716 4138 6772
rect 4194 6716 4280 6772
rect 4336 6716 4410 6772
rect 4070 6630 4410 6716
rect 4070 6574 4138 6630
rect 4194 6574 4280 6630
rect 4336 6574 4410 6630
rect 4070 6488 4410 6574
rect 4070 6432 4138 6488
rect 4194 6432 4280 6488
rect 4336 6432 4410 6488
rect 4070 6346 4410 6432
rect 4070 6290 4138 6346
rect 4194 6290 4280 6346
rect 4336 6290 4410 6346
rect 4070 6204 4410 6290
rect 4070 6148 4138 6204
rect 4194 6148 4280 6204
rect 4336 6148 4410 6204
rect 4070 6062 4410 6148
rect 4070 6006 4138 6062
rect 4194 6006 4280 6062
rect 4336 6006 4410 6062
rect 4070 5920 4410 6006
rect 4070 5864 4138 5920
rect 4194 5864 4280 5920
rect 4336 5864 4410 5920
rect 4070 5778 4410 5864
rect 4070 5722 4138 5778
rect 4194 5722 4280 5778
rect 4336 5722 4410 5778
rect 4070 5636 4410 5722
rect 4070 5580 4138 5636
rect 4194 5580 4280 5636
rect 4336 5580 4410 5636
rect 4070 5494 4410 5580
rect 4070 5438 4138 5494
rect 4194 5438 4280 5494
rect 4336 5438 4410 5494
rect 4070 5352 4410 5438
rect 4070 5296 4138 5352
rect 4194 5296 4280 5352
rect 4336 5296 4410 5352
rect 4070 5210 4410 5296
rect 4070 5154 4138 5210
rect 4194 5154 4280 5210
rect 4336 5154 4410 5210
rect 4070 5068 4410 5154
rect 4070 5012 4138 5068
rect 4194 5012 4280 5068
rect 4336 5012 4410 5068
rect 4070 4926 4410 5012
rect 4070 4870 4138 4926
rect 4194 4870 4280 4926
rect 4336 4870 4410 4926
rect 4070 4784 4410 4870
rect 4070 4728 4138 4784
rect 4194 4728 4280 4784
rect 4336 4728 4410 4784
rect 4070 4642 4410 4728
rect 4070 4586 4138 4642
rect 4194 4586 4280 4642
rect 4336 4586 4410 4642
rect 4070 4500 4410 4586
rect 4070 4444 4138 4500
rect 4194 4444 4280 4500
rect 4336 4444 4410 4500
rect 4070 4358 4410 4444
rect 4070 4302 4138 4358
rect 4194 4302 4280 4358
rect 4336 4302 4410 4358
rect 4070 4216 4410 4302
rect 4070 4160 4138 4216
rect 4194 4160 4280 4216
rect 4336 4160 4410 4216
rect 4070 4074 4410 4160
rect 4070 4018 4138 4074
rect 4194 4018 4280 4074
rect 4336 4018 4410 4074
rect 4070 3932 4410 4018
rect 4070 3876 4138 3932
rect 4194 3876 4280 3932
rect 4336 3876 4410 3932
rect 4070 3790 4410 3876
rect 4070 3734 4138 3790
rect 4194 3734 4280 3790
rect 4336 3734 4410 3790
rect 4070 3648 4410 3734
rect 4070 3592 4138 3648
rect 4194 3592 4280 3648
rect 4336 3592 4410 3648
rect 4070 3506 4410 3592
rect 4070 3450 4138 3506
rect 4194 3450 4280 3506
rect 4336 3450 4410 3506
rect 4070 3364 4410 3450
rect 4070 3308 4138 3364
rect 4194 3308 4280 3364
rect 4336 3308 4410 3364
rect 4070 3222 4410 3308
rect 4070 3166 4138 3222
rect 4194 3166 4280 3222
rect 4336 3166 4410 3222
rect 4070 3080 4410 3166
rect 4070 3024 4138 3080
rect 4194 3024 4280 3080
rect 4336 3024 4410 3080
rect 4070 2938 4410 3024
rect 4070 2882 4138 2938
rect 4194 2882 4280 2938
rect 4336 2882 4410 2938
rect 4070 2796 4410 2882
rect 4070 2740 4138 2796
rect 4194 2740 4280 2796
rect 4336 2740 4410 2796
rect 4070 2654 4410 2740
rect 4070 2598 4138 2654
rect 4194 2598 4280 2654
rect 4336 2598 4410 2654
rect 4070 2512 4410 2598
rect 4070 2456 4138 2512
rect 4194 2456 4280 2512
rect 4336 2456 4410 2512
rect 4070 2370 4410 2456
rect 4070 2314 4138 2370
rect 4194 2314 4280 2370
rect 4336 2314 4410 2370
rect 4070 2228 4410 2314
rect 4070 2172 4138 2228
rect 4194 2172 4280 2228
rect 4336 2172 4410 2228
rect 4070 2086 4410 2172
rect 4070 2030 4138 2086
rect 4194 2030 4280 2086
rect 4336 2030 4410 2086
rect 4070 1944 4410 2030
rect 4070 1888 4138 1944
rect 4194 1888 4280 1944
rect 4336 1888 4410 1944
rect 4070 1802 4410 1888
rect 4070 1746 4138 1802
rect 4194 1746 4280 1802
rect 4336 1746 4410 1802
rect 4070 1660 4410 1746
rect 4070 1604 4138 1660
rect 4194 1604 4280 1660
rect 4336 1604 4410 1660
rect 4070 1518 4410 1604
rect 4070 1462 4138 1518
rect 4194 1462 4280 1518
rect 4336 1462 4410 1518
rect 4070 1376 4410 1462
rect 4070 1320 4138 1376
rect 4194 1320 4280 1376
rect 4336 1320 4410 1376
rect 4070 1234 4410 1320
rect 4070 1178 4138 1234
rect 4194 1178 4280 1234
rect 4336 1178 4410 1234
rect 4070 1092 4410 1178
rect 4070 1036 4138 1092
rect 4194 1036 4280 1092
rect 4336 1036 4410 1092
rect 4070 950 4410 1036
rect 4070 894 4138 950
rect 4194 894 4280 950
rect 4336 894 4410 950
rect 4070 808 4410 894
rect 4070 752 4138 808
rect 4194 752 4280 808
rect 4336 752 4410 808
rect 4070 666 4410 752
rect 4070 610 4138 666
rect 4194 610 4280 666
rect 4336 610 4410 666
rect 4070 524 4410 610
rect 4070 468 4138 524
rect 4194 468 4280 524
rect 4336 468 4410 524
rect 4070 458 4410 468
rect 4610 12310 4950 12320
rect 4610 12254 4678 12310
rect 4734 12254 4820 12310
rect 4876 12254 4950 12310
rect 4610 12168 4950 12254
rect 4610 12112 4678 12168
rect 4734 12112 4820 12168
rect 4876 12112 4950 12168
rect 4610 12026 4950 12112
rect 4610 11970 4678 12026
rect 4734 11970 4820 12026
rect 4876 11970 4950 12026
rect 4610 11884 4950 11970
rect 4610 11828 4678 11884
rect 4734 11828 4820 11884
rect 4876 11828 4950 11884
rect 4610 11742 4950 11828
rect 4610 11686 4678 11742
rect 4734 11686 4820 11742
rect 4876 11686 4950 11742
rect 4610 11600 4950 11686
rect 4610 11544 4678 11600
rect 4734 11544 4820 11600
rect 4876 11544 4950 11600
rect 4610 11458 4950 11544
rect 4610 11402 4678 11458
rect 4734 11402 4820 11458
rect 4876 11402 4950 11458
rect 4610 11316 4950 11402
rect 4610 11260 4678 11316
rect 4734 11260 4820 11316
rect 4876 11260 4950 11316
rect 4610 11174 4950 11260
rect 4610 11118 4678 11174
rect 4734 11118 4820 11174
rect 4876 11118 4950 11174
rect 4610 11032 4950 11118
rect 4610 10976 4678 11032
rect 4734 10976 4820 11032
rect 4876 10976 4950 11032
rect 4610 10890 4950 10976
rect 4610 10834 4678 10890
rect 4734 10834 4820 10890
rect 4876 10834 4950 10890
rect 4610 10748 4950 10834
rect 4610 10692 4678 10748
rect 4734 10692 4820 10748
rect 4876 10692 4950 10748
rect 4610 10606 4950 10692
rect 4610 10550 4678 10606
rect 4734 10550 4820 10606
rect 4876 10550 4950 10606
rect 4610 10464 4950 10550
rect 4610 10408 4678 10464
rect 4734 10408 4820 10464
rect 4876 10408 4950 10464
rect 4610 10322 4950 10408
rect 4610 10266 4678 10322
rect 4734 10266 4820 10322
rect 4876 10266 4950 10322
rect 4610 10180 4950 10266
rect 4610 10124 4678 10180
rect 4734 10124 4820 10180
rect 4876 10124 4950 10180
rect 4610 10038 4950 10124
rect 4610 9982 4678 10038
rect 4734 9982 4820 10038
rect 4876 9982 4950 10038
rect 4610 9896 4950 9982
rect 4610 9840 4678 9896
rect 4734 9840 4820 9896
rect 4876 9840 4950 9896
rect 4610 9754 4950 9840
rect 4610 9698 4678 9754
rect 4734 9698 4820 9754
rect 4876 9698 4950 9754
rect 4610 9612 4950 9698
rect 4610 9556 4678 9612
rect 4734 9556 4820 9612
rect 4876 9556 4950 9612
rect 4610 9470 4950 9556
rect 4610 9414 4678 9470
rect 4734 9414 4820 9470
rect 4876 9414 4950 9470
rect 4610 9328 4950 9414
rect 4610 9272 4678 9328
rect 4734 9272 4820 9328
rect 4876 9272 4950 9328
rect 4610 9186 4950 9272
rect 4610 9130 4678 9186
rect 4734 9130 4820 9186
rect 4876 9130 4950 9186
rect 4610 9044 4950 9130
rect 4610 8988 4678 9044
rect 4734 8988 4820 9044
rect 4876 8988 4950 9044
rect 4610 8902 4950 8988
rect 4610 8846 4678 8902
rect 4734 8846 4820 8902
rect 4876 8846 4950 8902
rect 4610 8760 4950 8846
rect 4610 8704 4678 8760
rect 4734 8704 4820 8760
rect 4876 8704 4950 8760
rect 4610 8618 4950 8704
rect 4610 8562 4678 8618
rect 4734 8562 4820 8618
rect 4876 8562 4950 8618
rect 4610 8476 4950 8562
rect 4610 8420 4678 8476
rect 4734 8420 4820 8476
rect 4876 8420 4950 8476
rect 4610 8334 4950 8420
rect 4610 8278 4678 8334
rect 4734 8278 4820 8334
rect 4876 8278 4950 8334
rect 4610 8192 4950 8278
rect 4610 8136 4678 8192
rect 4734 8136 4820 8192
rect 4876 8136 4950 8192
rect 4610 8050 4950 8136
rect 4610 7994 4678 8050
rect 4734 7994 4820 8050
rect 4876 7994 4950 8050
rect 4610 7908 4950 7994
rect 4610 7852 4678 7908
rect 4734 7852 4820 7908
rect 4876 7852 4950 7908
rect 4610 7766 4950 7852
rect 4610 7710 4678 7766
rect 4734 7710 4820 7766
rect 4876 7710 4950 7766
rect 4610 7624 4950 7710
rect 4610 7568 4678 7624
rect 4734 7568 4820 7624
rect 4876 7568 4950 7624
rect 4610 7482 4950 7568
rect 4610 7426 4678 7482
rect 4734 7426 4820 7482
rect 4876 7426 4950 7482
rect 4610 7340 4950 7426
rect 4610 7284 4678 7340
rect 4734 7284 4820 7340
rect 4876 7284 4950 7340
rect 4610 7198 4950 7284
rect 4610 7142 4678 7198
rect 4734 7142 4820 7198
rect 4876 7142 4950 7198
rect 4610 7056 4950 7142
rect 4610 7000 4678 7056
rect 4734 7000 4820 7056
rect 4876 7000 4950 7056
rect 4610 6914 4950 7000
rect 4610 6858 4678 6914
rect 4734 6858 4820 6914
rect 4876 6858 4950 6914
rect 4610 6772 4950 6858
rect 4610 6716 4678 6772
rect 4734 6716 4820 6772
rect 4876 6716 4950 6772
rect 4610 6630 4950 6716
rect 4610 6574 4678 6630
rect 4734 6574 4820 6630
rect 4876 6574 4950 6630
rect 4610 6488 4950 6574
rect 4610 6432 4678 6488
rect 4734 6432 4820 6488
rect 4876 6432 4950 6488
rect 4610 6346 4950 6432
rect 4610 6290 4678 6346
rect 4734 6290 4820 6346
rect 4876 6290 4950 6346
rect 4610 6204 4950 6290
rect 4610 6148 4678 6204
rect 4734 6148 4820 6204
rect 4876 6148 4950 6204
rect 4610 6062 4950 6148
rect 4610 6006 4678 6062
rect 4734 6006 4820 6062
rect 4876 6006 4950 6062
rect 4610 5920 4950 6006
rect 4610 5864 4678 5920
rect 4734 5864 4820 5920
rect 4876 5864 4950 5920
rect 4610 5778 4950 5864
rect 4610 5722 4678 5778
rect 4734 5722 4820 5778
rect 4876 5722 4950 5778
rect 4610 5636 4950 5722
rect 4610 5580 4678 5636
rect 4734 5580 4820 5636
rect 4876 5580 4950 5636
rect 4610 5494 4950 5580
rect 4610 5438 4678 5494
rect 4734 5438 4820 5494
rect 4876 5438 4950 5494
rect 4610 5352 4950 5438
rect 4610 5296 4678 5352
rect 4734 5296 4820 5352
rect 4876 5296 4950 5352
rect 4610 5210 4950 5296
rect 4610 5154 4678 5210
rect 4734 5154 4820 5210
rect 4876 5154 4950 5210
rect 4610 5068 4950 5154
rect 4610 5012 4678 5068
rect 4734 5012 4820 5068
rect 4876 5012 4950 5068
rect 4610 4926 4950 5012
rect 4610 4870 4678 4926
rect 4734 4870 4820 4926
rect 4876 4870 4950 4926
rect 4610 4784 4950 4870
rect 4610 4728 4678 4784
rect 4734 4728 4820 4784
rect 4876 4728 4950 4784
rect 4610 4642 4950 4728
rect 4610 4586 4678 4642
rect 4734 4586 4820 4642
rect 4876 4586 4950 4642
rect 4610 4500 4950 4586
rect 4610 4444 4678 4500
rect 4734 4444 4820 4500
rect 4876 4444 4950 4500
rect 4610 4358 4950 4444
rect 4610 4302 4678 4358
rect 4734 4302 4820 4358
rect 4876 4302 4950 4358
rect 4610 4216 4950 4302
rect 4610 4160 4678 4216
rect 4734 4160 4820 4216
rect 4876 4160 4950 4216
rect 4610 4074 4950 4160
rect 4610 4018 4678 4074
rect 4734 4018 4820 4074
rect 4876 4018 4950 4074
rect 4610 3932 4950 4018
rect 4610 3876 4678 3932
rect 4734 3876 4820 3932
rect 4876 3876 4950 3932
rect 4610 3790 4950 3876
rect 4610 3734 4678 3790
rect 4734 3734 4820 3790
rect 4876 3734 4950 3790
rect 4610 3648 4950 3734
rect 4610 3592 4678 3648
rect 4734 3592 4820 3648
rect 4876 3592 4950 3648
rect 4610 3506 4950 3592
rect 4610 3450 4678 3506
rect 4734 3450 4820 3506
rect 4876 3450 4950 3506
rect 4610 3364 4950 3450
rect 4610 3308 4678 3364
rect 4734 3308 4820 3364
rect 4876 3308 4950 3364
rect 4610 3222 4950 3308
rect 4610 3166 4678 3222
rect 4734 3166 4820 3222
rect 4876 3166 4950 3222
rect 4610 3080 4950 3166
rect 4610 3024 4678 3080
rect 4734 3024 4820 3080
rect 4876 3024 4950 3080
rect 4610 2938 4950 3024
rect 4610 2882 4678 2938
rect 4734 2882 4820 2938
rect 4876 2882 4950 2938
rect 4610 2796 4950 2882
rect 4610 2740 4678 2796
rect 4734 2740 4820 2796
rect 4876 2740 4950 2796
rect 4610 2654 4950 2740
rect 4610 2598 4678 2654
rect 4734 2598 4820 2654
rect 4876 2598 4950 2654
rect 4610 2512 4950 2598
rect 4610 2456 4678 2512
rect 4734 2456 4820 2512
rect 4876 2456 4950 2512
rect 4610 2370 4950 2456
rect 4610 2314 4678 2370
rect 4734 2314 4820 2370
rect 4876 2314 4950 2370
rect 4610 2228 4950 2314
rect 4610 2172 4678 2228
rect 4734 2172 4820 2228
rect 4876 2172 4950 2228
rect 4610 2086 4950 2172
rect 4610 2030 4678 2086
rect 4734 2030 4820 2086
rect 4876 2030 4950 2086
rect 4610 1944 4950 2030
rect 4610 1888 4678 1944
rect 4734 1888 4820 1944
rect 4876 1888 4950 1944
rect 4610 1802 4950 1888
rect 4610 1746 4678 1802
rect 4734 1746 4820 1802
rect 4876 1746 4950 1802
rect 4610 1660 4950 1746
rect 4610 1604 4678 1660
rect 4734 1604 4820 1660
rect 4876 1604 4950 1660
rect 4610 1518 4950 1604
rect 4610 1462 4678 1518
rect 4734 1462 4820 1518
rect 4876 1462 4950 1518
rect 4610 1376 4950 1462
rect 4610 1320 4678 1376
rect 4734 1320 4820 1376
rect 4876 1320 4950 1376
rect 4610 1234 4950 1320
rect 4610 1178 4678 1234
rect 4734 1178 4820 1234
rect 4876 1178 4950 1234
rect 4610 1092 4950 1178
rect 4610 1036 4678 1092
rect 4734 1036 4820 1092
rect 4876 1036 4950 1092
rect 4610 950 4950 1036
rect 4610 894 4678 950
rect 4734 894 4820 950
rect 4876 894 4950 950
rect 4610 808 4950 894
rect 4610 752 4678 808
rect 4734 752 4820 808
rect 4876 752 4950 808
rect 4610 666 4950 752
rect 4610 610 4678 666
rect 4734 610 4820 666
rect 4876 610 4950 666
rect 4610 524 4950 610
rect 4610 468 4678 524
rect 4734 468 4820 524
rect 4876 468 4950 524
rect 4610 458 4950 468
rect 5150 12310 5490 12320
rect 5150 12254 5215 12310
rect 5271 12254 5357 12310
rect 5413 12254 5490 12310
rect 5150 12168 5490 12254
rect 5150 12112 5215 12168
rect 5271 12112 5357 12168
rect 5413 12112 5490 12168
rect 5150 12026 5490 12112
rect 5150 11970 5215 12026
rect 5271 11970 5357 12026
rect 5413 11970 5490 12026
rect 5150 11884 5490 11970
rect 5150 11828 5215 11884
rect 5271 11828 5357 11884
rect 5413 11828 5490 11884
rect 5150 11742 5490 11828
rect 5150 11686 5215 11742
rect 5271 11686 5357 11742
rect 5413 11686 5490 11742
rect 5150 11600 5490 11686
rect 5150 11544 5215 11600
rect 5271 11544 5357 11600
rect 5413 11544 5490 11600
rect 5150 11458 5490 11544
rect 5150 11402 5215 11458
rect 5271 11402 5357 11458
rect 5413 11402 5490 11458
rect 5150 11316 5490 11402
rect 5150 11260 5215 11316
rect 5271 11260 5357 11316
rect 5413 11260 5490 11316
rect 5150 11174 5490 11260
rect 5150 11118 5215 11174
rect 5271 11118 5357 11174
rect 5413 11118 5490 11174
rect 5150 11032 5490 11118
rect 5150 10976 5215 11032
rect 5271 10976 5357 11032
rect 5413 10976 5490 11032
rect 5150 10890 5490 10976
rect 5150 10834 5215 10890
rect 5271 10834 5357 10890
rect 5413 10834 5490 10890
rect 5150 10748 5490 10834
rect 5150 10692 5215 10748
rect 5271 10692 5357 10748
rect 5413 10692 5490 10748
rect 5150 10606 5490 10692
rect 5150 10550 5215 10606
rect 5271 10550 5357 10606
rect 5413 10550 5490 10606
rect 5150 10464 5490 10550
rect 5150 10408 5215 10464
rect 5271 10408 5357 10464
rect 5413 10408 5490 10464
rect 5150 10322 5490 10408
rect 5150 10266 5215 10322
rect 5271 10266 5357 10322
rect 5413 10266 5490 10322
rect 5150 10180 5490 10266
rect 5150 10124 5215 10180
rect 5271 10124 5357 10180
rect 5413 10124 5490 10180
rect 5150 10038 5490 10124
rect 5150 9982 5215 10038
rect 5271 9982 5357 10038
rect 5413 9982 5490 10038
rect 5150 9896 5490 9982
rect 5150 9840 5215 9896
rect 5271 9840 5357 9896
rect 5413 9840 5490 9896
rect 5150 9754 5490 9840
rect 5150 9698 5215 9754
rect 5271 9698 5357 9754
rect 5413 9698 5490 9754
rect 5150 9612 5490 9698
rect 5150 9556 5215 9612
rect 5271 9556 5357 9612
rect 5413 9556 5490 9612
rect 5150 9470 5490 9556
rect 5150 9414 5215 9470
rect 5271 9414 5357 9470
rect 5413 9414 5490 9470
rect 5150 9328 5490 9414
rect 5150 9272 5215 9328
rect 5271 9272 5357 9328
rect 5413 9272 5490 9328
rect 5150 9186 5490 9272
rect 5150 9130 5215 9186
rect 5271 9130 5357 9186
rect 5413 9130 5490 9186
rect 5150 9044 5490 9130
rect 5150 8988 5215 9044
rect 5271 8988 5357 9044
rect 5413 8988 5490 9044
rect 5150 8902 5490 8988
rect 5150 8846 5215 8902
rect 5271 8846 5357 8902
rect 5413 8846 5490 8902
rect 5150 8760 5490 8846
rect 5150 8704 5215 8760
rect 5271 8704 5357 8760
rect 5413 8704 5490 8760
rect 5150 8618 5490 8704
rect 5150 8562 5215 8618
rect 5271 8562 5357 8618
rect 5413 8562 5490 8618
rect 5150 8476 5490 8562
rect 5150 8420 5215 8476
rect 5271 8420 5357 8476
rect 5413 8420 5490 8476
rect 5150 8334 5490 8420
rect 5150 8278 5215 8334
rect 5271 8278 5357 8334
rect 5413 8278 5490 8334
rect 5150 8192 5490 8278
rect 5150 8136 5215 8192
rect 5271 8136 5357 8192
rect 5413 8136 5490 8192
rect 5150 8050 5490 8136
rect 5150 7994 5215 8050
rect 5271 7994 5357 8050
rect 5413 7994 5490 8050
rect 5150 7908 5490 7994
rect 5150 7852 5215 7908
rect 5271 7852 5357 7908
rect 5413 7852 5490 7908
rect 5150 7766 5490 7852
rect 5150 7710 5215 7766
rect 5271 7710 5357 7766
rect 5413 7710 5490 7766
rect 5150 7624 5490 7710
rect 5150 7568 5215 7624
rect 5271 7568 5357 7624
rect 5413 7568 5490 7624
rect 5150 7482 5490 7568
rect 5150 7426 5215 7482
rect 5271 7426 5357 7482
rect 5413 7426 5490 7482
rect 5150 7340 5490 7426
rect 5150 7284 5215 7340
rect 5271 7284 5357 7340
rect 5413 7284 5490 7340
rect 5150 7198 5490 7284
rect 5150 7142 5215 7198
rect 5271 7142 5357 7198
rect 5413 7142 5490 7198
rect 5150 7056 5490 7142
rect 5150 7000 5215 7056
rect 5271 7000 5357 7056
rect 5413 7000 5490 7056
rect 5150 6914 5490 7000
rect 5150 6858 5215 6914
rect 5271 6858 5357 6914
rect 5413 6858 5490 6914
rect 5150 6772 5490 6858
rect 5150 6716 5215 6772
rect 5271 6716 5357 6772
rect 5413 6716 5490 6772
rect 5150 6630 5490 6716
rect 5150 6574 5215 6630
rect 5271 6574 5357 6630
rect 5413 6574 5490 6630
rect 5150 6488 5490 6574
rect 5150 6432 5215 6488
rect 5271 6432 5357 6488
rect 5413 6432 5490 6488
rect 5150 6346 5490 6432
rect 5150 6290 5215 6346
rect 5271 6290 5357 6346
rect 5413 6290 5490 6346
rect 5150 6204 5490 6290
rect 5150 6148 5215 6204
rect 5271 6148 5357 6204
rect 5413 6148 5490 6204
rect 5150 6062 5490 6148
rect 5150 6006 5215 6062
rect 5271 6006 5357 6062
rect 5413 6006 5490 6062
rect 5150 5920 5490 6006
rect 5150 5864 5215 5920
rect 5271 5864 5357 5920
rect 5413 5864 5490 5920
rect 5150 5778 5490 5864
rect 5150 5722 5215 5778
rect 5271 5722 5357 5778
rect 5413 5722 5490 5778
rect 5150 5636 5490 5722
rect 5150 5580 5215 5636
rect 5271 5580 5357 5636
rect 5413 5580 5490 5636
rect 5150 5494 5490 5580
rect 5150 5438 5215 5494
rect 5271 5438 5357 5494
rect 5413 5438 5490 5494
rect 5150 5352 5490 5438
rect 5150 5296 5215 5352
rect 5271 5296 5357 5352
rect 5413 5296 5490 5352
rect 5150 5210 5490 5296
rect 5150 5154 5215 5210
rect 5271 5154 5357 5210
rect 5413 5154 5490 5210
rect 5150 5068 5490 5154
rect 5150 5012 5215 5068
rect 5271 5012 5357 5068
rect 5413 5012 5490 5068
rect 5150 4926 5490 5012
rect 5150 4870 5215 4926
rect 5271 4870 5357 4926
rect 5413 4870 5490 4926
rect 5150 4784 5490 4870
rect 5150 4728 5215 4784
rect 5271 4728 5357 4784
rect 5413 4728 5490 4784
rect 5150 4642 5490 4728
rect 5150 4586 5215 4642
rect 5271 4586 5357 4642
rect 5413 4586 5490 4642
rect 5150 4500 5490 4586
rect 5150 4444 5215 4500
rect 5271 4444 5357 4500
rect 5413 4444 5490 4500
rect 5150 4358 5490 4444
rect 5150 4302 5215 4358
rect 5271 4302 5357 4358
rect 5413 4302 5490 4358
rect 5150 4216 5490 4302
rect 5150 4160 5215 4216
rect 5271 4160 5357 4216
rect 5413 4160 5490 4216
rect 5150 4074 5490 4160
rect 5150 4018 5215 4074
rect 5271 4018 5357 4074
rect 5413 4018 5490 4074
rect 5150 3932 5490 4018
rect 5150 3876 5215 3932
rect 5271 3876 5357 3932
rect 5413 3876 5490 3932
rect 5150 3790 5490 3876
rect 5150 3734 5215 3790
rect 5271 3734 5357 3790
rect 5413 3734 5490 3790
rect 5150 3648 5490 3734
rect 5150 3592 5215 3648
rect 5271 3592 5357 3648
rect 5413 3592 5490 3648
rect 5150 3506 5490 3592
rect 5150 3450 5215 3506
rect 5271 3450 5357 3506
rect 5413 3450 5490 3506
rect 5150 3364 5490 3450
rect 5150 3308 5215 3364
rect 5271 3308 5357 3364
rect 5413 3308 5490 3364
rect 5150 3222 5490 3308
rect 5150 3166 5215 3222
rect 5271 3166 5357 3222
rect 5413 3166 5490 3222
rect 5150 3080 5490 3166
rect 5150 3024 5215 3080
rect 5271 3024 5357 3080
rect 5413 3024 5490 3080
rect 5150 2938 5490 3024
rect 5150 2882 5215 2938
rect 5271 2882 5357 2938
rect 5413 2882 5490 2938
rect 5150 2796 5490 2882
rect 5150 2740 5215 2796
rect 5271 2740 5357 2796
rect 5413 2740 5490 2796
rect 5150 2654 5490 2740
rect 5150 2598 5215 2654
rect 5271 2598 5357 2654
rect 5413 2598 5490 2654
rect 5150 2512 5490 2598
rect 5150 2456 5215 2512
rect 5271 2456 5357 2512
rect 5413 2456 5490 2512
rect 5150 2370 5490 2456
rect 5150 2314 5215 2370
rect 5271 2314 5357 2370
rect 5413 2314 5490 2370
rect 5150 2228 5490 2314
rect 5150 2172 5215 2228
rect 5271 2172 5357 2228
rect 5413 2172 5490 2228
rect 5150 2086 5490 2172
rect 5150 2030 5215 2086
rect 5271 2030 5357 2086
rect 5413 2030 5490 2086
rect 5150 1944 5490 2030
rect 5150 1888 5215 1944
rect 5271 1888 5357 1944
rect 5413 1888 5490 1944
rect 5150 1802 5490 1888
rect 5150 1746 5215 1802
rect 5271 1746 5357 1802
rect 5413 1746 5490 1802
rect 5150 1660 5490 1746
rect 5150 1604 5215 1660
rect 5271 1604 5357 1660
rect 5413 1604 5490 1660
rect 5150 1518 5490 1604
rect 5150 1462 5215 1518
rect 5271 1462 5357 1518
rect 5413 1462 5490 1518
rect 5150 1376 5490 1462
rect 5150 1320 5215 1376
rect 5271 1320 5357 1376
rect 5413 1320 5490 1376
rect 5150 1234 5490 1320
rect 5150 1178 5215 1234
rect 5271 1178 5357 1234
rect 5413 1178 5490 1234
rect 5150 1092 5490 1178
rect 5150 1036 5215 1092
rect 5271 1036 5357 1092
rect 5413 1036 5490 1092
rect 5150 950 5490 1036
rect 5150 894 5215 950
rect 5271 894 5357 950
rect 5413 894 5490 950
rect 5150 808 5490 894
rect 5150 752 5215 808
rect 5271 752 5357 808
rect 5413 752 5490 808
rect 5150 666 5490 752
rect 5150 610 5215 666
rect 5271 610 5357 666
rect 5413 610 5490 666
rect 5150 524 5490 610
rect 5150 468 5215 524
rect 5271 468 5357 524
rect 5413 468 5490 524
rect 5150 458 5490 468
rect 5690 12310 6030 12320
rect 5690 12254 5760 12310
rect 5816 12254 5902 12310
rect 5958 12254 6030 12310
rect 5690 12168 6030 12254
rect 5690 12112 5760 12168
rect 5816 12112 5902 12168
rect 5958 12112 6030 12168
rect 5690 12026 6030 12112
rect 5690 11970 5760 12026
rect 5816 11970 5902 12026
rect 5958 11970 6030 12026
rect 5690 11884 6030 11970
rect 5690 11828 5760 11884
rect 5816 11828 5902 11884
rect 5958 11828 6030 11884
rect 5690 11742 6030 11828
rect 5690 11686 5760 11742
rect 5816 11686 5902 11742
rect 5958 11686 6030 11742
rect 5690 11600 6030 11686
rect 5690 11544 5760 11600
rect 5816 11544 5902 11600
rect 5958 11544 6030 11600
rect 5690 11458 6030 11544
rect 5690 11402 5760 11458
rect 5816 11402 5902 11458
rect 5958 11402 6030 11458
rect 5690 11316 6030 11402
rect 5690 11260 5760 11316
rect 5816 11260 5902 11316
rect 5958 11260 6030 11316
rect 5690 11174 6030 11260
rect 5690 11118 5760 11174
rect 5816 11118 5902 11174
rect 5958 11118 6030 11174
rect 5690 11032 6030 11118
rect 5690 10976 5760 11032
rect 5816 10976 5902 11032
rect 5958 10976 6030 11032
rect 5690 10890 6030 10976
rect 5690 10834 5760 10890
rect 5816 10834 5902 10890
rect 5958 10834 6030 10890
rect 5690 10748 6030 10834
rect 5690 10692 5760 10748
rect 5816 10692 5902 10748
rect 5958 10692 6030 10748
rect 5690 10606 6030 10692
rect 5690 10550 5760 10606
rect 5816 10550 5902 10606
rect 5958 10550 6030 10606
rect 5690 10464 6030 10550
rect 5690 10408 5760 10464
rect 5816 10408 5902 10464
rect 5958 10408 6030 10464
rect 5690 10322 6030 10408
rect 5690 10266 5760 10322
rect 5816 10266 5902 10322
rect 5958 10266 6030 10322
rect 5690 10180 6030 10266
rect 5690 10124 5760 10180
rect 5816 10124 5902 10180
rect 5958 10124 6030 10180
rect 5690 10038 6030 10124
rect 5690 9982 5760 10038
rect 5816 9982 5902 10038
rect 5958 9982 6030 10038
rect 5690 9896 6030 9982
rect 5690 9840 5760 9896
rect 5816 9840 5902 9896
rect 5958 9840 6030 9896
rect 5690 9754 6030 9840
rect 5690 9698 5760 9754
rect 5816 9698 5902 9754
rect 5958 9698 6030 9754
rect 5690 9612 6030 9698
rect 5690 9556 5760 9612
rect 5816 9556 5902 9612
rect 5958 9556 6030 9612
rect 5690 9470 6030 9556
rect 5690 9414 5760 9470
rect 5816 9414 5902 9470
rect 5958 9414 6030 9470
rect 5690 9328 6030 9414
rect 5690 9272 5760 9328
rect 5816 9272 5902 9328
rect 5958 9272 6030 9328
rect 5690 9186 6030 9272
rect 5690 9130 5760 9186
rect 5816 9130 5902 9186
rect 5958 9130 6030 9186
rect 5690 9044 6030 9130
rect 5690 8988 5760 9044
rect 5816 8988 5902 9044
rect 5958 8988 6030 9044
rect 5690 8902 6030 8988
rect 5690 8846 5760 8902
rect 5816 8846 5902 8902
rect 5958 8846 6030 8902
rect 5690 8760 6030 8846
rect 5690 8704 5760 8760
rect 5816 8704 5902 8760
rect 5958 8704 6030 8760
rect 5690 8618 6030 8704
rect 5690 8562 5760 8618
rect 5816 8562 5902 8618
rect 5958 8562 6030 8618
rect 5690 8476 6030 8562
rect 5690 8420 5760 8476
rect 5816 8420 5902 8476
rect 5958 8420 6030 8476
rect 5690 8334 6030 8420
rect 5690 8278 5760 8334
rect 5816 8278 5902 8334
rect 5958 8278 6030 8334
rect 5690 8192 6030 8278
rect 5690 8136 5760 8192
rect 5816 8136 5902 8192
rect 5958 8136 6030 8192
rect 5690 8050 6030 8136
rect 5690 7994 5760 8050
rect 5816 7994 5902 8050
rect 5958 7994 6030 8050
rect 5690 7908 6030 7994
rect 5690 7852 5760 7908
rect 5816 7852 5902 7908
rect 5958 7852 6030 7908
rect 5690 7766 6030 7852
rect 5690 7710 5760 7766
rect 5816 7710 5902 7766
rect 5958 7710 6030 7766
rect 5690 7624 6030 7710
rect 5690 7568 5760 7624
rect 5816 7568 5902 7624
rect 5958 7568 6030 7624
rect 5690 7482 6030 7568
rect 5690 7426 5760 7482
rect 5816 7426 5902 7482
rect 5958 7426 6030 7482
rect 5690 7340 6030 7426
rect 5690 7284 5760 7340
rect 5816 7284 5902 7340
rect 5958 7284 6030 7340
rect 5690 7198 6030 7284
rect 5690 7142 5760 7198
rect 5816 7142 5902 7198
rect 5958 7142 6030 7198
rect 5690 7056 6030 7142
rect 5690 7000 5760 7056
rect 5816 7000 5902 7056
rect 5958 7000 6030 7056
rect 5690 6914 6030 7000
rect 5690 6858 5760 6914
rect 5816 6858 5902 6914
rect 5958 6858 6030 6914
rect 5690 6772 6030 6858
rect 5690 6716 5760 6772
rect 5816 6716 5902 6772
rect 5958 6716 6030 6772
rect 5690 6630 6030 6716
rect 5690 6574 5760 6630
rect 5816 6574 5902 6630
rect 5958 6574 6030 6630
rect 5690 6488 6030 6574
rect 5690 6432 5760 6488
rect 5816 6432 5902 6488
rect 5958 6432 6030 6488
rect 5690 6346 6030 6432
rect 5690 6290 5760 6346
rect 5816 6290 5902 6346
rect 5958 6290 6030 6346
rect 5690 6204 6030 6290
rect 5690 6148 5760 6204
rect 5816 6148 5902 6204
rect 5958 6148 6030 6204
rect 5690 6062 6030 6148
rect 5690 6006 5760 6062
rect 5816 6006 5902 6062
rect 5958 6006 6030 6062
rect 5690 5920 6030 6006
rect 5690 5864 5760 5920
rect 5816 5864 5902 5920
rect 5958 5864 6030 5920
rect 5690 5778 6030 5864
rect 5690 5722 5760 5778
rect 5816 5722 5902 5778
rect 5958 5722 6030 5778
rect 5690 5636 6030 5722
rect 5690 5580 5760 5636
rect 5816 5580 5902 5636
rect 5958 5580 6030 5636
rect 5690 5494 6030 5580
rect 5690 5438 5760 5494
rect 5816 5438 5902 5494
rect 5958 5438 6030 5494
rect 5690 5352 6030 5438
rect 5690 5296 5760 5352
rect 5816 5296 5902 5352
rect 5958 5296 6030 5352
rect 5690 5210 6030 5296
rect 5690 5154 5760 5210
rect 5816 5154 5902 5210
rect 5958 5154 6030 5210
rect 5690 5068 6030 5154
rect 5690 5012 5760 5068
rect 5816 5012 5902 5068
rect 5958 5012 6030 5068
rect 5690 4926 6030 5012
rect 5690 4870 5760 4926
rect 5816 4870 5902 4926
rect 5958 4870 6030 4926
rect 5690 4784 6030 4870
rect 5690 4728 5760 4784
rect 5816 4728 5902 4784
rect 5958 4728 6030 4784
rect 5690 4642 6030 4728
rect 5690 4586 5760 4642
rect 5816 4586 5902 4642
rect 5958 4586 6030 4642
rect 5690 4500 6030 4586
rect 5690 4444 5760 4500
rect 5816 4444 5902 4500
rect 5958 4444 6030 4500
rect 5690 4358 6030 4444
rect 5690 4302 5760 4358
rect 5816 4302 5902 4358
rect 5958 4302 6030 4358
rect 5690 4216 6030 4302
rect 5690 4160 5760 4216
rect 5816 4160 5902 4216
rect 5958 4160 6030 4216
rect 5690 4074 6030 4160
rect 5690 4018 5760 4074
rect 5816 4018 5902 4074
rect 5958 4018 6030 4074
rect 5690 3932 6030 4018
rect 5690 3876 5760 3932
rect 5816 3876 5902 3932
rect 5958 3876 6030 3932
rect 5690 3790 6030 3876
rect 5690 3734 5760 3790
rect 5816 3734 5902 3790
rect 5958 3734 6030 3790
rect 5690 3648 6030 3734
rect 5690 3592 5760 3648
rect 5816 3592 5902 3648
rect 5958 3592 6030 3648
rect 5690 3506 6030 3592
rect 5690 3450 5760 3506
rect 5816 3450 5902 3506
rect 5958 3450 6030 3506
rect 5690 3364 6030 3450
rect 5690 3308 5760 3364
rect 5816 3308 5902 3364
rect 5958 3308 6030 3364
rect 5690 3222 6030 3308
rect 5690 3166 5760 3222
rect 5816 3166 5902 3222
rect 5958 3166 6030 3222
rect 5690 3080 6030 3166
rect 5690 3024 5760 3080
rect 5816 3024 5902 3080
rect 5958 3024 6030 3080
rect 5690 2938 6030 3024
rect 5690 2882 5760 2938
rect 5816 2882 5902 2938
rect 5958 2882 6030 2938
rect 5690 2796 6030 2882
rect 5690 2740 5760 2796
rect 5816 2740 5902 2796
rect 5958 2740 6030 2796
rect 5690 2654 6030 2740
rect 5690 2598 5760 2654
rect 5816 2598 5902 2654
rect 5958 2598 6030 2654
rect 5690 2512 6030 2598
rect 5690 2456 5760 2512
rect 5816 2456 5902 2512
rect 5958 2456 6030 2512
rect 5690 2370 6030 2456
rect 5690 2314 5760 2370
rect 5816 2314 5902 2370
rect 5958 2314 6030 2370
rect 5690 2228 6030 2314
rect 5690 2172 5760 2228
rect 5816 2172 5902 2228
rect 5958 2172 6030 2228
rect 5690 2086 6030 2172
rect 5690 2030 5760 2086
rect 5816 2030 5902 2086
rect 5958 2030 6030 2086
rect 5690 1944 6030 2030
rect 5690 1888 5760 1944
rect 5816 1888 5902 1944
rect 5958 1888 6030 1944
rect 5690 1802 6030 1888
rect 5690 1746 5760 1802
rect 5816 1746 5902 1802
rect 5958 1746 6030 1802
rect 5690 1660 6030 1746
rect 5690 1604 5760 1660
rect 5816 1604 5902 1660
rect 5958 1604 6030 1660
rect 5690 1518 6030 1604
rect 5690 1462 5760 1518
rect 5816 1462 5902 1518
rect 5958 1462 6030 1518
rect 5690 1376 6030 1462
rect 5690 1320 5760 1376
rect 5816 1320 5902 1376
rect 5958 1320 6030 1376
rect 5690 1234 6030 1320
rect 5690 1178 5760 1234
rect 5816 1178 5902 1234
rect 5958 1178 6030 1234
rect 5690 1092 6030 1178
rect 5690 1036 5760 1092
rect 5816 1036 5902 1092
rect 5958 1036 6030 1092
rect 5690 950 6030 1036
rect 5690 894 5760 950
rect 5816 894 5902 950
rect 5958 894 6030 950
rect 5690 808 6030 894
rect 5690 752 5760 808
rect 5816 752 5902 808
rect 5958 752 6030 808
rect 5690 666 6030 752
rect 5690 610 5760 666
rect 5816 610 5902 666
rect 5958 610 6030 666
rect 5690 524 6030 610
rect 5690 468 5760 524
rect 5816 468 5902 524
rect 5958 468 6030 524
rect 5690 458 6030 468
rect 6230 12310 6570 12320
rect 6230 12254 6300 12310
rect 6356 12254 6442 12310
rect 6498 12254 6570 12310
rect 6230 12168 6570 12254
rect 6230 12112 6300 12168
rect 6356 12112 6442 12168
rect 6498 12112 6570 12168
rect 6230 12026 6570 12112
rect 6230 11970 6300 12026
rect 6356 11970 6442 12026
rect 6498 11970 6570 12026
rect 6230 11884 6570 11970
rect 6230 11828 6300 11884
rect 6356 11828 6442 11884
rect 6498 11828 6570 11884
rect 6230 11742 6570 11828
rect 6230 11686 6300 11742
rect 6356 11686 6442 11742
rect 6498 11686 6570 11742
rect 6230 11600 6570 11686
rect 6230 11544 6300 11600
rect 6356 11544 6442 11600
rect 6498 11544 6570 11600
rect 6230 11458 6570 11544
rect 6230 11402 6300 11458
rect 6356 11402 6442 11458
rect 6498 11402 6570 11458
rect 6230 11316 6570 11402
rect 6230 11260 6300 11316
rect 6356 11260 6442 11316
rect 6498 11260 6570 11316
rect 6230 11174 6570 11260
rect 6230 11118 6300 11174
rect 6356 11118 6442 11174
rect 6498 11118 6570 11174
rect 6230 11032 6570 11118
rect 6230 10976 6300 11032
rect 6356 10976 6442 11032
rect 6498 10976 6570 11032
rect 6230 10890 6570 10976
rect 6230 10834 6300 10890
rect 6356 10834 6442 10890
rect 6498 10834 6570 10890
rect 6230 10748 6570 10834
rect 6230 10692 6300 10748
rect 6356 10692 6442 10748
rect 6498 10692 6570 10748
rect 6230 10606 6570 10692
rect 6230 10550 6300 10606
rect 6356 10550 6442 10606
rect 6498 10550 6570 10606
rect 6230 10464 6570 10550
rect 6230 10408 6300 10464
rect 6356 10408 6442 10464
rect 6498 10408 6570 10464
rect 6230 10322 6570 10408
rect 6230 10266 6300 10322
rect 6356 10266 6442 10322
rect 6498 10266 6570 10322
rect 6230 10180 6570 10266
rect 6230 10124 6300 10180
rect 6356 10124 6442 10180
rect 6498 10124 6570 10180
rect 6230 10038 6570 10124
rect 6230 9982 6300 10038
rect 6356 9982 6442 10038
rect 6498 9982 6570 10038
rect 6230 9896 6570 9982
rect 6230 9840 6300 9896
rect 6356 9840 6442 9896
rect 6498 9840 6570 9896
rect 6230 9754 6570 9840
rect 6230 9698 6300 9754
rect 6356 9698 6442 9754
rect 6498 9698 6570 9754
rect 6230 9612 6570 9698
rect 6230 9556 6300 9612
rect 6356 9556 6442 9612
rect 6498 9556 6570 9612
rect 6230 9470 6570 9556
rect 6230 9414 6300 9470
rect 6356 9414 6442 9470
rect 6498 9414 6570 9470
rect 6230 9328 6570 9414
rect 6230 9272 6300 9328
rect 6356 9272 6442 9328
rect 6498 9272 6570 9328
rect 6230 9186 6570 9272
rect 6230 9130 6300 9186
rect 6356 9130 6442 9186
rect 6498 9130 6570 9186
rect 6230 9044 6570 9130
rect 6230 8988 6300 9044
rect 6356 8988 6442 9044
rect 6498 8988 6570 9044
rect 6230 8902 6570 8988
rect 6230 8846 6300 8902
rect 6356 8846 6442 8902
rect 6498 8846 6570 8902
rect 6230 8760 6570 8846
rect 6230 8704 6300 8760
rect 6356 8704 6442 8760
rect 6498 8704 6570 8760
rect 6230 8618 6570 8704
rect 6230 8562 6300 8618
rect 6356 8562 6442 8618
rect 6498 8562 6570 8618
rect 6230 8476 6570 8562
rect 6230 8420 6300 8476
rect 6356 8420 6442 8476
rect 6498 8420 6570 8476
rect 6230 8334 6570 8420
rect 6230 8278 6300 8334
rect 6356 8278 6442 8334
rect 6498 8278 6570 8334
rect 6230 8192 6570 8278
rect 6230 8136 6300 8192
rect 6356 8136 6442 8192
rect 6498 8136 6570 8192
rect 6230 8050 6570 8136
rect 6230 7994 6300 8050
rect 6356 7994 6442 8050
rect 6498 7994 6570 8050
rect 6230 7908 6570 7994
rect 6230 7852 6300 7908
rect 6356 7852 6442 7908
rect 6498 7852 6570 7908
rect 6230 7766 6570 7852
rect 6230 7710 6300 7766
rect 6356 7710 6442 7766
rect 6498 7710 6570 7766
rect 6230 7624 6570 7710
rect 6230 7568 6300 7624
rect 6356 7568 6442 7624
rect 6498 7568 6570 7624
rect 6230 7482 6570 7568
rect 6230 7426 6300 7482
rect 6356 7426 6442 7482
rect 6498 7426 6570 7482
rect 6230 7340 6570 7426
rect 6230 7284 6300 7340
rect 6356 7284 6442 7340
rect 6498 7284 6570 7340
rect 6230 7198 6570 7284
rect 6230 7142 6300 7198
rect 6356 7142 6442 7198
rect 6498 7142 6570 7198
rect 6230 7056 6570 7142
rect 6230 7000 6300 7056
rect 6356 7000 6442 7056
rect 6498 7000 6570 7056
rect 6230 6914 6570 7000
rect 6230 6858 6300 6914
rect 6356 6858 6442 6914
rect 6498 6858 6570 6914
rect 6230 6772 6570 6858
rect 6230 6716 6300 6772
rect 6356 6716 6442 6772
rect 6498 6716 6570 6772
rect 6230 6630 6570 6716
rect 6230 6574 6300 6630
rect 6356 6574 6442 6630
rect 6498 6574 6570 6630
rect 6230 6488 6570 6574
rect 6230 6432 6300 6488
rect 6356 6432 6442 6488
rect 6498 6432 6570 6488
rect 6230 6346 6570 6432
rect 6230 6290 6300 6346
rect 6356 6290 6442 6346
rect 6498 6290 6570 6346
rect 6230 6204 6570 6290
rect 6230 6148 6300 6204
rect 6356 6148 6442 6204
rect 6498 6148 6570 6204
rect 6230 6062 6570 6148
rect 6230 6006 6300 6062
rect 6356 6006 6442 6062
rect 6498 6006 6570 6062
rect 6230 5920 6570 6006
rect 6230 5864 6300 5920
rect 6356 5864 6442 5920
rect 6498 5864 6570 5920
rect 6230 5778 6570 5864
rect 6230 5722 6300 5778
rect 6356 5722 6442 5778
rect 6498 5722 6570 5778
rect 6230 5636 6570 5722
rect 6230 5580 6300 5636
rect 6356 5580 6442 5636
rect 6498 5580 6570 5636
rect 6230 5494 6570 5580
rect 6230 5438 6300 5494
rect 6356 5438 6442 5494
rect 6498 5438 6570 5494
rect 6230 5352 6570 5438
rect 6230 5296 6300 5352
rect 6356 5296 6442 5352
rect 6498 5296 6570 5352
rect 6230 5210 6570 5296
rect 6230 5154 6300 5210
rect 6356 5154 6442 5210
rect 6498 5154 6570 5210
rect 6230 5068 6570 5154
rect 6230 5012 6300 5068
rect 6356 5012 6442 5068
rect 6498 5012 6570 5068
rect 6230 4926 6570 5012
rect 6230 4870 6300 4926
rect 6356 4870 6442 4926
rect 6498 4870 6570 4926
rect 6230 4784 6570 4870
rect 6230 4728 6300 4784
rect 6356 4728 6442 4784
rect 6498 4728 6570 4784
rect 6230 4642 6570 4728
rect 6230 4586 6300 4642
rect 6356 4586 6442 4642
rect 6498 4586 6570 4642
rect 6230 4500 6570 4586
rect 6230 4444 6300 4500
rect 6356 4444 6442 4500
rect 6498 4444 6570 4500
rect 6230 4358 6570 4444
rect 6230 4302 6300 4358
rect 6356 4302 6442 4358
rect 6498 4302 6570 4358
rect 6230 4216 6570 4302
rect 6230 4160 6300 4216
rect 6356 4160 6442 4216
rect 6498 4160 6570 4216
rect 6230 4074 6570 4160
rect 6230 4018 6300 4074
rect 6356 4018 6442 4074
rect 6498 4018 6570 4074
rect 6230 3932 6570 4018
rect 6230 3876 6300 3932
rect 6356 3876 6442 3932
rect 6498 3876 6570 3932
rect 6230 3790 6570 3876
rect 6230 3734 6300 3790
rect 6356 3734 6442 3790
rect 6498 3734 6570 3790
rect 6230 3648 6570 3734
rect 6230 3592 6300 3648
rect 6356 3592 6442 3648
rect 6498 3592 6570 3648
rect 6230 3506 6570 3592
rect 6230 3450 6300 3506
rect 6356 3450 6442 3506
rect 6498 3450 6570 3506
rect 6230 3364 6570 3450
rect 6230 3308 6300 3364
rect 6356 3308 6442 3364
rect 6498 3308 6570 3364
rect 6230 3222 6570 3308
rect 6230 3166 6300 3222
rect 6356 3166 6442 3222
rect 6498 3166 6570 3222
rect 6230 3080 6570 3166
rect 6230 3024 6300 3080
rect 6356 3024 6442 3080
rect 6498 3024 6570 3080
rect 6230 2938 6570 3024
rect 6230 2882 6300 2938
rect 6356 2882 6442 2938
rect 6498 2882 6570 2938
rect 6230 2796 6570 2882
rect 6230 2740 6300 2796
rect 6356 2740 6442 2796
rect 6498 2740 6570 2796
rect 6230 2654 6570 2740
rect 6230 2598 6300 2654
rect 6356 2598 6442 2654
rect 6498 2598 6570 2654
rect 6230 2512 6570 2598
rect 6230 2456 6300 2512
rect 6356 2456 6442 2512
rect 6498 2456 6570 2512
rect 6230 2370 6570 2456
rect 6230 2314 6300 2370
rect 6356 2314 6442 2370
rect 6498 2314 6570 2370
rect 6230 2228 6570 2314
rect 6230 2172 6300 2228
rect 6356 2172 6442 2228
rect 6498 2172 6570 2228
rect 6230 2086 6570 2172
rect 6230 2030 6300 2086
rect 6356 2030 6442 2086
rect 6498 2030 6570 2086
rect 6230 1944 6570 2030
rect 6230 1888 6300 1944
rect 6356 1888 6442 1944
rect 6498 1888 6570 1944
rect 6230 1802 6570 1888
rect 6230 1746 6300 1802
rect 6356 1746 6442 1802
rect 6498 1746 6570 1802
rect 6230 1660 6570 1746
rect 6230 1604 6300 1660
rect 6356 1604 6442 1660
rect 6498 1604 6570 1660
rect 6230 1518 6570 1604
rect 6230 1462 6300 1518
rect 6356 1462 6442 1518
rect 6498 1462 6570 1518
rect 6230 1376 6570 1462
rect 6230 1320 6300 1376
rect 6356 1320 6442 1376
rect 6498 1320 6570 1376
rect 6230 1234 6570 1320
rect 6230 1178 6300 1234
rect 6356 1178 6442 1234
rect 6498 1178 6570 1234
rect 6230 1092 6570 1178
rect 6230 1036 6300 1092
rect 6356 1036 6442 1092
rect 6498 1036 6570 1092
rect 6230 950 6570 1036
rect 6230 894 6300 950
rect 6356 894 6442 950
rect 6498 894 6570 950
rect 6230 808 6570 894
rect 6230 752 6300 808
rect 6356 752 6442 808
rect 6498 752 6570 808
rect 6230 666 6570 752
rect 6230 610 6300 666
rect 6356 610 6442 666
rect 6498 610 6570 666
rect 6230 524 6570 610
rect 6230 468 6300 524
rect 6356 468 6442 524
rect 6498 468 6570 524
rect 6230 458 6570 468
rect 6770 12310 7110 12320
rect 6770 12254 6845 12310
rect 6901 12254 6987 12310
rect 7043 12254 7110 12310
rect 6770 12168 7110 12254
rect 6770 12112 6845 12168
rect 6901 12112 6987 12168
rect 7043 12112 7110 12168
rect 6770 12026 7110 12112
rect 6770 11970 6845 12026
rect 6901 11970 6987 12026
rect 7043 11970 7110 12026
rect 6770 11884 7110 11970
rect 6770 11828 6845 11884
rect 6901 11828 6987 11884
rect 7043 11828 7110 11884
rect 6770 11742 7110 11828
rect 6770 11686 6845 11742
rect 6901 11686 6987 11742
rect 7043 11686 7110 11742
rect 6770 11600 7110 11686
rect 6770 11544 6845 11600
rect 6901 11544 6987 11600
rect 7043 11544 7110 11600
rect 6770 11458 7110 11544
rect 6770 11402 6845 11458
rect 6901 11402 6987 11458
rect 7043 11402 7110 11458
rect 6770 11316 7110 11402
rect 6770 11260 6845 11316
rect 6901 11260 6987 11316
rect 7043 11260 7110 11316
rect 6770 11174 7110 11260
rect 6770 11118 6845 11174
rect 6901 11118 6987 11174
rect 7043 11118 7110 11174
rect 6770 11032 7110 11118
rect 6770 10976 6845 11032
rect 6901 10976 6987 11032
rect 7043 10976 7110 11032
rect 6770 10890 7110 10976
rect 6770 10834 6845 10890
rect 6901 10834 6987 10890
rect 7043 10834 7110 10890
rect 6770 10748 7110 10834
rect 6770 10692 6845 10748
rect 6901 10692 6987 10748
rect 7043 10692 7110 10748
rect 6770 10606 7110 10692
rect 6770 10550 6845 10606
rect 6901 10550 6987 10606
rect 7043 10550 7110 10606
rect 6770 10464 7110 10550
rect 6770 10408 6845 10464
rect 6901 10408 6987 10464
rect 7043 10408 7110 10464
rect 6770 10322 7110 10408
rect 6770 10266 6845 10322
rect 6901 10266 6987 10322
rect 7043 10266 7110 10322
rect 6770 10180 7110 10266
rect 6770 10124 6845 10180
rect 6901 10124 6987 10180
rect 7043 10124 7110 10180
rect 6770 10038 7110 10124
rect 6770 9982 6845 10038
rect 6901 9982 6987 10038
rect 7043 9982 7110 10038
rect 6770 9896 7110 9982
rect 6770 9840 6845 9896
rect 6901 9840 6987 9896
rect 7043 9840 7110 9896
rect 6770 9754 7110 9840
rect 6770 9698 6845 9754
rect 6901 9698 6987 9754
rect 7043 9698 7110 9754
rect 6770 9612 7110 9698
rect 6770 9556 6845 9612
rect 6901 9556 6987 9612
rect 7043 9556 7110 9612
rect 6770 9470 7110 9556
rect 6770 9414 6845 9470
rect 6901 9414 6987 9470
rect 7043 9414 7110 9470
rect 6770 9328 7110 9414
rect 6770 9272 6845 9328
rect 6901 9272 6987 9328
rect 7043 9272 7110 9328
rect 6770 9186 7110 9272
rect 6770 9130 6845 9186
rect 6901 9130 6987 9186
rect 7043 9130 7110 9186
rect 6770 9044 7110 9130
rect 6770 8988 6845 9044
rect 6901 8988 6987 9044
rect 7043 8988 7110 9044
rect 6770 8902 7110 8988
rect 6770 8846 6845 8902
rect 6901 8846 6987 8902
rect 7043 8846 7110 8902
rect 6770 8760 7110 8846
rect 6770 8704 6845 8760
rect 6901 8704 6987 8760
rect 7043 8704 7110 8760
rect 6770 8618 7110 8704
rect 6770 8562 6845 8618
rect 6901 8562 6987 8618
rect 7043 8562 7110 8618
rect 6770 8476 7110 8562
rect 6770 8420 6845 8476
rect 6901 8420 6987 8476
rect 7043 8420 7110 8476
rect 6770 8334 7110 8420
rect 6770 8278 6845 8334
rect 6901 8278 6987 8334
rect 7043 8278 7110 8334
rect 6770 8192 7110 8278
rect 6770 8136 6845 8192
rect 6901 8136 6987 8192
rect 7043 8136 7110 8192
rect 6770 8050 7110 8136
rect 6770 7994 6845 8050
rect 6901 7994 6987 8050
rect 7043 7994 7110 8050
rect 6770 7908 7110 7994
rect 6770 7852 6845 7908
rect 6901 7852 6987 7908
rect 7043 7852 7110 7908
rect 6770 7766 7110 7852
rect 6770 7710 6845 7766
rect 6901 7710 6987 7766
rect 7043 7710 7110 7766
rect 6770 7624 7110 7710
rect 6770 7568 6845 7624
rect 6901 7568 6987 7624
rect 7043 7568 7110 7624
rect 6770 7482 7110 7568
rect 6770 7426 6845 7482
rect 6901 7426 6987 7482
rect 7043 7426 7110 7482
rect 6770 7340 7110 7426
rect 6770 7284 6845 7340
rect 6901 7284 6987 7340
rect 7043 7284 7110 7340
rect 6770 7198 7110 7284
rect 6770 7142 6845 7198
rect 6901 7142 6987 7198
rect 7043 7142 7110 7198
rect 6770 7056 7110 7142
rect 6770 7000 6845 7056
rect 6901 7000 6987 7056
rect 7043 7000 7110 7056
rect 6770 6914 7110 7000
rect 6770 6858 6845 6914
rect 6901 6858 6987 6914
rect 7043 6858 7110 6914
rect 6770 6772 7110 6858
rect 6770 6716 6845 6772
rect 6901 6716 6987 6772
rect 7043 6716 7110 6772
rect 6770 6630 7110 6716
rect 6770 6574 6845 6630
rect 6901 6574 6987 6630
rect 7043 6574 7110 6630
rect 6770 6488 7110 6574
rect 6770 6432 6845 6488
rect 6901 6432 6987 6488
rect 7043 6432 7110 6488
rect 6770 6346 7110 6432
rect 6770 6290 6845 6346
rect 6901 6290 6987 6346
rect 7043 6290 7110 6346
rect 6770 6204 7110 6290
rect 6770 6148 6845 6204
rect 6901 6148 6987 6204
rect 7043 6148 7110 6204
rect 6770 6062 7110 6148
rect 6770 6006 6845 6062
rect 6901 6006 6987 6062
rect 7043 6006 7110 6062
rect 6770 5920 7110 6006
rect 6770 5864 6845 5920
rect 6901 5864 6987 5920
rect 7043 5864 7110 5920
rect 6770 5778 7110 5864
rect 6770 5722 6845 5778
rect 6901 5722 6987 5778
rect 7043 5722 7110 5778
rect 6770 5636 7110 5722
rect 6770 5580 6845 5636
rect 6901 5580 6987 5636
rect 7043 5580 7110 5636
rect 6770 5494 7110 5580
rect 6770 5438 6845 5494
rect 6901 5438 6987 5494
rect 7043 5438 7110 5494
rect 6770 5352 7110 5438
rect 6770 5296 6845 5352
rect 6901 5296 6987 5352
rect 7043 5296 7110 5352
rect 6770 5210 7110 5296
rect 6770 5154 6845 5210
rect 6901 5154 6987 5210
rect 7043 5154 7110 5210
rect 6770 5068 7110 5154
rect 6770 5012 6845 5068
rect 6901 5012 6987 5068
rect 7043 5012 7110 5068
rect 6770 4926 7110 5012
rect 6770 4870 6845 4926
rect 6901 4870 6987 4926
rect 7043 4870 7110 4926
rect 6770 4784 7110 4870
rect 6770 4728 6845 4784
rect 6901 4728 6987 4784
rect 7043 4728 7110 4784
rect 6770 4642 7110 4728
rect 6770 4586 6845 4642
rect 6901 4586 6987 4642
rect 7043 4586 7110 4642
rect 6770 4500 7110 4586
rect 6770 4444 6845 4500
rect 6901 4444 6987 4500
rect 7043 4444 7110 4500
rect 6770 4358 7110 4444
rect 6770 4302 6845 4358
rect 6901 4302 6987 4358
rect 7043 4302 7110 4358
rect 6770 4216 7110 4302
rect 6770 4160 6845 4216
rect 6901 4160 6987 4216
rect 7043 4160 7110 4216
rect 6770 4074 7110 4160
rect 6770 4018 6845 4074
rect 6901 4018 6987 4074
rect 7043 4018 7110 4074
rect 6770 3932 7110 4018
rect 6770 3876 6845 3932
rect 6901 3876 6987 3932
rect 7043 3876 7110 3932
rect 6770 3790 7110 3876
rect 6770 3734 6845 3790
rect 6901 3734 6987 3790
rect 7043 3734 7110 3790
rect 6770 3648 7110 3734
rect 6770 3592 6845 3648
rect 6901 3592 6987 3648
rect 7043 3592 7110 3648
rect 6770 3506 7110 3592
rect 6770 3450 6845 3506
rect 6901 3450 6987 3506
rect 7043 3450 7110 3506
rect 6770 3364 7110 3450
rect 6770 3308 6845 3364
rect 6901 3308 6987 3364
rect 7043 3308 7110 3364
rect 6770 3222 7110 3308
rect 6770 3166 6845 3222
rect 6901 3166 6987 3222
rect 7043 3166 7110 3222
rect 6770 3080 7110 3166
rect 6770 3024 6845 3080
rect 6901 3024 6987 3080
rect 7043 3024 7110 3080
rect 6770 2938 7110 3024
rect 6770 2882 6845 2938
rect 6901 2882 6987 2938
rect 7043 2882 7110 2938
rect 6770 2796 7110 2882
rect 6770 2740 6845 2796
rect 6901 2740 6987 2796
rect 7043 2740 7110 2796
rect 6770 2654 7110 2740
rect 6770 2598 6845 2654
rect 6901 2598 6987 2654
rect 7043 2598 7110 2654
rect 6770 2512 7110 2598
rect 6770 2456 6845 2512
rect 6901 2456 6987 2512
rect 7043 2456 7110 2512
rect 6770 2370 7110 2456
rect 6770 2314 6845 2370
rect 6901 2314 6987 2370
rect 7043 2314 7110 2370
rect 6770 2228 7110 2314
rect 6770 2172 6845 2228
rect 6901 2172 6987 2228
rect 7043 2172 7110 2228
rect 6770 2086 7110 2172
rect 6770 2030 6845 2086
rect 6901 2030 6987 2086
rect 7043 2030 7110 2086
rect 6770 1944 7110 2030
rect 6770 1888 6845 1944
rect 6901 1888 6987 1944
rect 7043 1888 7110 1944
rect 6770 1802 7110 1888
rect 6770 1746 6845 1802
rect 6901 1746 6987 1802
rect 7043 1746 7110 1802
rect 6770 1660 7110 1746
rect 6770 1604 6845 1660
rect 6901 1604 6987 1660
rect 7043 1604 7110 1660
rect 6770 1518 7110 1604
rect 6770 1462 6845 1518
rect 6901 1462 6987 1518
rect 7043 1462 7110 1518
rect 6770 1376 7110 1462
rect 6770 1320 6845 1376
rect 6901 1320 6987 1376
rect 7043 1320 7110 1376
rect 6770 1234 7110 1320
rect 6770 1178 6845 1234
rect 6901 1178 6987 1234
rect 7043 1178 7110 1234
rect 6770 1092 7110 1178
rect 6770 1036 6845 1092
rect 6901 1036 6987 1092
rect 7043 1036 7110 1092
rect 6770 950 7110 1036
rect 6770 894 6845 950
rect 6901 894 6987 950
rect 7043 894 7110 950
rect 6770 808 7110 894
rect 6770 752 6845 808
rect 6901 752 6987 808
rect 7043 752 7110 808
rect 6770 666 7110 752
rect 6770 610 6845 666
rect 6901 610 6987 666
rect 7043 610 7110 666
rect 6770 524 7110 610
rect 6770 468 6845 524
rect 6901 468 6987 524
rect 7043 468 7110 524
rect 6770 458 7110 468
rect 7310 12310 7650 12320
rect 7310 12254 7382 12310
rect 7438 12254 7524 12310
rect 7580 12254 7650 12310
rect 7310 12168 7650 12254
rect 7310 12112 7382 12168
rect 7438 12112 7524 12168
rect 7580 12112 7650 12168
rect 7310 12026 7650 12112
rect 7310 11970 7382 12026
rect 7438 11970 7524 12026
rect 7580 11970 7650 12026
rect 7310 11884 7650 11970
rect 7310 11828 7382 11884
rect 7438 11828 7524 11884
rect 7580 11828 7650 11884
rect 7310 11742 7650 11828
rect 7310 11686 7382 11742
rect 7438 11686 7524 11742
rect 7580 11686 7650 11742
rect 7310 11600 7650 11686
rect 7310 11544 7382 11600
rect 7438 11544 7524 11600
rect 7580 11544 7650 11600
rect 7310 11458 7650 11544
rect 7310 11402 7382 11458
rect 7438 11402 7524 11458
rect 7580 11402 7650 11458
rect 7310 11316 7650 11402
rect 7310 11260 7382 11316
rect 7438 11260 7524 11316
rect 7580 11260 7650 11316
rect 7310 11174 7650 11260
rect 7310 11118 7382 11174
rect 7438 11118 7524 11174
rect 7580 11118 7650 11174
rect 7310 11032 7650 11118
rect 7310 10976 7382 11032
rect 7438 10976 7524 11032
rect 7580 10976 7650 11032
rect 7310 10890 7650 10976
rect 7310 10834 7382 10890
rect 7438 10834 7524 10890
rect 7580 10834 7650 10890
rect 7310 10748 7650 10834
rect 7310 10692 7382 10748
rect 7438 10692 7524 10748
rect 7580 10692 7650 10748
rect 7310 10606 7650 10692
rect 7310 10550 7382 10606
rect 7438 10550 7524 10606
rect 7580 10550 7650 10606
rect 7310 10464 7650 10550
rect 7310 10408 7382 10464
rect 7438 10408 7524 10464
rect 7580 10408 7650 10464
rect 7310 10322 7650 10408
rect 7310 10266 7382 10322
rect 7438 10266 7524 10322
rect 7580 10266 7650 10322
rect 7310 10180 7650 10266
rect 7310 10124 7382 10180
rect 7438 10124 7524 10180
rect 7580 10124 7650 10180
rect 7310 10038 7650 10124
rect 7310 9982 7382 10038
rect 7438 9982 7524 10038
rect 7580 9982 7650 10038
rect 7310 9896 7650 9982
rect 7310 9840 7382 9896
rect 7438 9840 7524 9896
rect 7580 9840 7650 9896
rect 7310 9754 7650 9840
rect 7310 9698 7382 9754
rect 7438 9698 7524 9754
rect 7580 9698 7650 9754
rect 7310 9612 7650 9698
rect 7310 9556 7382 9612
rect 7438 9556 7524 9612
rect 7580 9556 7650 9612
rect 7310 9470 7650 9556
rect 7310 9414 7382 9470
rect 7438 9414 7524 9470
rect 7580 9414 7650 9470
rect 7310 9328 7650 9414
rect 7310 9272 7382 9328
rect 7438 9272 7524 9328
rect 7580 9272 7650 9328
rect 7310 9186 7650 9272
rect 7310 9130 7382 9186
rect 7438 9130 7524 9186
rect 7580 9130 7650 9186
rect 7310 9044 7650 9130
rect 7310 8988 7382 9044
rect 7438 8988 7524 9044
rect 7580 8988 7650 9044
rect 7310 8902 7650 8988
rect 7310 8846 7382 8902
rect 7438 8846 7524 8902
rect 7580 8846 7650 8902
rect 7310 8760 7650 8846
rect 7310 8704 7382 8760
rect 7438 8704 7524 8760
rect 7580 8704 7650 8760
rect 7310 8618 7650 8704
rect 7310 8562 7382 8618
rect 7438 8562 7524 8618
rect 7580 8562 7650 8618
rect 7310 8476 7650 8562
rect 7310 8420 7382 8476
rect 7438 8420 7524 8476
rect 7580 8420 7650 8476
rect 7310 8334 7650 8420
rect 7310 8278 7382 8334
rect 7438 8278 7524 8334
rect 7580 8278 7650 8334
rect 7310 8192 7650 8278
rect 7310 8136 7382 8192
rect 7438 8136 7524 8192
rect 7580 8136 7650 8192
rect 7310 8050 7650 8136
rect 7310 7994 7382 8050
rect 7438 7994 7524 8050
rect 7580 7994 7650 8050
rect 7310 7908 7650 7994
rect 7310 7852 7382 7908
rect 7438 7852 7524 7908
rect 7580 7852 7650 7908
rect 7310 7766 7650 7852
rect 7310 7710 7382 7766
rect 7438 7710 7524 7766
rect 7580 7710 7650 7766
rect 7310 7624 7650 7710
rect 7310 7568 7382 7624
rect 7438 7568 7524 7624
rect 7580 7568 7650 7624
rect 7310 7482 7650 7568
rect 7310 7426 7382 7482
rect 7438 7426 7524 7482
rect 7580 7426 7650 7482
rect 7310 7340 7650 7426
rect 7310 7284 7382 7340
rect 7438 7284 7524 7340
rect 7580 7284 7650 7340
rect 7310 7198 7650 7284
rect 7310 7142 7382 7198
rect 7438 7142 7524 7198
rect 7580 7142 7650 7198
rect 7310 7056 7650 7142
rect 7310 7000 7382 7056
rect 7438 7000 7524 7056
rect 7580 7000 7650 7056
rect 7310 6914 7650 7000
rect 7310 6858 7382 6914
rect 7438 6858 7524 6914
rect 7580 6858 7650 6914
rect 7310 6772 7650 6858
rect 7310 6716 7382 6772
rect 7438 6716 7524 6772
rect 7580 6716 7650 6772
rect 7310 6630 7650 6716
rect 7310 6574 7382 6630
rect 7438 6574 7524 6630
rect 7580 6574 7650 6630
rect 7310 6488 7650 6574
rect 7310 6432 7382 6488
rect 7438 6432 7524 6488
rect 7580 6432 7650 6488
rect 7310 6346 7650 6432
rect 7310 6290 7382 6346
rect 7438 6290 7524 6346
rect 7580 6290 7650 6346
rect 7310 6204 7650 6290
rect 7310 6148 7382 6204
rect 7438 6148 7524 6204
rect 7580 6148 7650 6204
rect 7310 6062 7650 6148
rect 7310 6006 7382 6062
rect 7438 6006 7524 6062
rect 7580 6006 7650 6062
rect 7310 5920 7650 6006
rect 7310 5864 7382 5920
rect 7438 5864 7524 5920
rect 7580 5864 7650 5920
rect 7310 5778 7650 5864
rect 7310 5722 7382 5778
rect 7438 5722 7524 5778
rect 7580 5722 7650 5778
rect 7310 5636 7650 5722
rect 7310 5580 7382 5636
rect 7438 5580 7524 5636
rect 7580 5580 7650 5636
rect 7310 5494 7650 5580
rect 7310 5438 7382 5494
rect 7438 5438 7524 5494
rect 7580 5438 7650 5494
rect 7310 5352 7650 5438
rect 7310 5296 7382 5352
rect 7438 5296 7524 5352
rect 7580 5296 7650 5352
rect 7310 5210 7650 5296
rect 7310 5154 7382 5210
rect 7438 5154 7524 5210
rect 7580 5154 7650 5210
rect 7310 5068 7650 5154
rect 7310 5012 7382 5068
rect 7438 5012 7524 5068
rect 7580 5012 7650 5068
rect 7310 4926 7650 5012
rect 7310 4870 7382 4926
rect 7438 4870 7524 4926
rect 7580 4870 7650 4926
rect 7310 4784 7650 4870
rect 7310 4728 7382 4784
rect 7438 4728 7524 4784
rect 7580 4728 7650 4784
rect 7310 4642 7650 4728
rect 7310 4586 7382 4642
rect 7438 4586 7524 4642
rect 7580 4586 7650 4642
rect 7310 4500 7650 4586
rect 7310 4444 7382 4500
rect 7438 4444 7524 4500
rect 7580 4444 7650 4500
rect 7310 4358 7650 4444
rect 7310 4302 7382 4358
rect 7438 4302 7524 4358
rect 7580 4302 7650 4358
rect 7310 4216 7650 4302
rect 7310 4160 7382 4216
rect 7438 4160 7524 4216
rect 7580 4160 7650 4216
rect 7310 4074 7650 4160
rect 7310 4018 7382 4074
rect 7438 4018 7524 4074
rect 7580 4018 7650 4074
rect 7310 3932 7650 4018
rect 7310 3876 7382 3932
rect 7438 3876 7524 3932
rect 7580 3876 7650 3932
rect 7310 3790 7650 3876
rect 7310 3734 7382 3790
rect 7438 3734 7524 3790
rect 7580 3734 7650 3790
rect 7310 3648 7650 3734
rect 7310 3592 7382 3648
rect 7438 3592 7524 3648
rect 7580 3592 7650 3648
rect 7310 3506 7650 3592
rect 7310 3450 7382 3506
rect 7438 3450 7524 3506
rect 7580 3450 7650 3506
rect 7310 3364 7650 3450
rect 7310 3308 7382 3364
rect 7438 3308 7524 3364
rect 7580 3308 7650 3364
rect 7310 3222 7650 3308
rect 7310 3166 7382 3222
rect 7438 3166 7524 3222
rect 7580 3166 7650 3222
rect 7310 3080 7650 3166
rect 7310 3024 7382 3080
rect 7438 3024 7524 3080
rect 7580 3024 7650 3080
rect 7310 2938 7650 3024
rect 7310 2882 7382 2938
rect 7438 2882 7524 2938
rect 7580 2882 7650 2938
rect 7310 2796 7650 2882
rect 7310 2740 7382 2796
rect 7438 2740 7524 2796
rect 7580 2740 7650 2796
rect 7310 2654 7650 2740
rect 7310 2598 7382 2654
rect 7438 2598 7524 2654
rect 7580 2598 7650 2654
rect 7310 2512 7650 2598
rect 7310 2456 7382 2512
rect 7438 2456 7524 2512
rect 7580 2456 7650 2512
rect 7310 2370 7650 2456
rect 7310 2314 7382 2370
rect 7438 2314 7524 2370
rect 7580 2314 7650 2370
rect 7310 2228 7650 2314
rect 7310 2172 7382 2228
rect 7438 2172 7524 2228
rect 7580 2172 7650 2228
rect 7310 2086 7650 2172
rect 7310 2030 7382 2086
rect 7438 2030 7524 2086
rect 7580 2030 7650 2086
rect 7310 1944 7650 2030
rect 7310 1888 7382 1944
rect 7438 1888 7524 1944
rect 7580 1888 7650 1944
rect 7310 1802 7650 1888
rect 7310 1746 7382 1802
rect 7438 1746 7524 1802
rect 7580 1746 7650 1802
rect 7310 1660 7650 1746
rect 7310 1604 7382 1660
rect 7438 1604 7524 1660
rect 7580 1604 7650 1660
rect 7310 1518 7650 1604
rect 7310 1462 7382 1518
rect 7438 1462 7524 1518
rect 7580 1462 7650 1518
rect 7310 1376 7650 1462
rect 7310 1320 7382 1376
rect 7438 1320 7524 1376
rect 7580 1320 7650 1376
rect 7310 1234 7650 1320
rect 7310 1178 7382 1234
rect 7438 1178 7524 1234
rect 7580 1178 7650 1234
rect 7310 1092 7650 1178
rect 7310 1036 7382 1092
rect 7438 1036 7524 1092
rect 7580 1036 7650 1092
rect 7310 950 7650 1036
rect 7310 894 7382 950
rect 7438 894 7524 950
rect 7580 894 7650 950
rect 7310 808 7650 894
rect 7310 752 7382 808
rect 7438 752 7524 808
rect 7580 752 7650 808
rect 7310 666 7650 752
rect 7310 610 7382 666
rect 7438 610 7524 666
rect 7580 610 7650 666
rect 7310 524 7650 610
rect 7310 468 7382 524
rect 7438 468 7524 524
rect 7580 468 7650 524
rect 7310 458 7650 468
rect 7850 12310 8190 12320
rect 7850 12254 7919 12310
rect 7975 12254 8061 12310
rect 8117 12254 8190 12310
rect 7850 12168 8190 12254
rect 7850 12112 7919 12168
rect 7975 12112 8061 12168
rect 8117 12112 8190 12168
rect 7850 12026 8190 12112
rect 7850 11970 7919 12026
rect 7975 11970 8061 12026
rect 8117 11970 8190 12026
rect 7850 11884 8190 11970
rect 7850 11828 7919 11884
rect 7975 11828 8061 11884
rect 8117 11828 8190 11884
rect 7850 11742 8190 11828
rect 7850 11686 7919 11742
rect 7975 11686 8061 11742
rect 8117 11686 8190 11742
rect 7850 11600 8190 11686
rect 7850 11544 7919 11600
rect 7975 11544 8061 11600
rect 8117 11544 8190 11600
rect 7850 11458 8190 11544
rect 7850 11402 7919 11458
rect 7975 11402 8061 11458
rect 8117 11402 8190 11458
rect 7850 11316 8190 11402
rect 7850 11260 7919 11316
rect 7975 11260 8061 11316
rect 8117 11260 8190 11316
rect 7850 11174 8190 11260
rect 7850 11118 7919 11174
rect 7975 11118 8061 11174
rect 8117 11118 8190 11174
rect 7850 11032 8190 11118
rect 7850 10976 7919 11032
rect 7975 10976 8061 11032
rect 8117 10976 8190 11032
rect 7850 10890 8190 10976
rect 7850 10834 7919 10890
rect 7975 10834 8061 10890
rect 8117 10834 8190 10890
rect 7850 10748 8190 10834
rect 7850 10692 7919 10748
rect 7975 10692 8061 10748
rect 8117 10692 8190 10748
rect 7850 10606 8190 10692
rect 7850 10550 7919 10606
rect 7975 10550 8061 10606
rect 8117 10550 8190 10606
rect 7850 10464 8190 10550
rect 7850 10408 7919 10464
rect 7975 10408 8061 10464
rect 8117 10408 8190 10464
rect 7850 10322 8190 10408
rect 7850 10266 7919 10322
rect 7975 10266 8061 10322
rect 8117 10266 8190 10322
rect 7850 10180 8190 10266
rect 7850 10124 7919 10180
rect 7975 10124 8061 10180
rect 8117 10124 8190 10180
rect 7850 10038 8190 10124
rect 7850 9982 7919 10038
rect 7975 9982 8061 10038
rect 8117 9982 8190 10038
rect 7850 9896 8190 9982
rect 7850 9840 7919 9896
rect 7975 9840 8061 9896
rect 8117 9840 8190 9896
rect 7850 9754 8190 9840
rect 7850 9698 7919 9754
rect 7975 9698 8061 9754
rect 8117 9698 8190 9754
rect 7850 9612 8190 9698
rect 7850 9556 7919 9612
rect 7975 9556 8061 9612
rect 8117 9556 8190 9612
rect 7850 9470 8190 9556
rect 7850 9414 7919 9470
rect 7975 9414 8061 9470
rect 8117 9414 8190 9470
rect 7850 9328 8190 9414
rect 7850 9272 7919 9328
rect 7975 9272 8061 9328
rect 8117 9272 8190 9328
rect 7850 9186 8190 9272
rect 7850 9130 7919 9186
rect 7975 9130 8061 9186
rect 8117 9130 8190 9186
rect 7850 9044 8190 9130
rect 7850 8988 7919 9044
rect 7975 8988 8061 9044
rect 8117 8988 8190 9044
rect 7850 8902 8190 8988
rect 7850 8846 7919 8902
rect 7975 8846 8061 8902
rect 8117 8846 8190 8902
rect 7850 8760 8190 8846
rect 7850 8704 7919 8760
rect 7975 8704 8061 8760
rect 8117 8704 8190 8760
rect 7850 8618 8190 8704
rect 7850 8562 7919 8618
rect 7975 8562 8061 8618
rect 8117 8562 8190 8618
rect 7850 8476 8190 8562
rect 7850 8420 7919 8476
rect 7975 8420 8061 8476
rect 8117 8420 8190 8476
rect 7850 8334 8190 8420
rect 7850 8278 7919 8334
rect 7975 8278 8061 8334
rect 8117 8278 8190 8334
rect 7850 8192 8190 8278
rect 7850 8136 7919 8192
rect 7975 8136 8061 8192
rect 8117 8136 8190 8192
rect 7850 8050 8190 8136
rect 7850 7994 7919 8050
rect 7975 7994 8061 8050
rect 8117 7994 8190 8050
rect 7850 7908 8190 7994
rect 7850 7852 7919 7908
rect 7975 7852 8061 7908
rect 8117 7852 8190 7908
rect 7850 7766 8190 7852
rect 7850 7710 7919 7766
rect 7975 7710 8061 7766
rect 8117 7710 8190 7766
rect 7850 7624 8190 7710
rect 7850 7568 7919 7624
rect 7975 7568 8061 7624
rect 8117 7568 8190 7624
rect 7850 7482 8190 7568
rect 7850 7426 7919 7482
rect 7975 7426 8061 7482
rect 8117 7426 8190 7482
rect 7850 7340 8190 7426
rect 7850 7284 7919 7340
rect 7975 7284 8061 7340
rect 8117 7284 8190 7340
rect 7850 7198 8190 7284
rect 7850 7142 7919 7198
rect 7975 7142 8061 7198
rect 8117 7142 8190 7198
rect 7850 7056 8190 7142
rect 7850 7000 7919 7056
rect 7975 7000 8061 7056
rect 8117 7000 8190 7056
rect 7850 6914 8190 7000
rect 7850 6858 7919 6914
rect 7975 6858 8061 6914
rect 8117 6858 8190 6914
rect 7850 6772 8190 6858
rect 7850 6716 7919 6772
rect 7975 6716 8061 6772
rect 8117 6716 8190 6772
rect 7850 6630 8190 6716
rect 7850 6574 7919 6630
rect 7975 6574 8061 6630
rect 8117 6574 8190 6630
rect 7850 6488 8190 6574
rect 7850 6432 7919 6488
rect 7975 6432 8061 6488
rect 8117 6432 8190 6488
rect 7850 6346 8190 6432
rect 7850 6290 7919 6346
rect 7975 6290 8061 6346
rect 8117 6290 8190 6346
rect 7850 6204 8190 6290
rect 7850 6148 7919 6204
rect 7975 6148 8061 6204
rect 8117 6148 8190 6204
rect 7850 6062 8190 6148
rect 7850 6006 7919 6062
rect 7975 6006 8061 6062
rect 8117 6006 8190 6062
rect 7850 5920 8190 6006
rect 7850 5864 7919 5920
rect 7975 5864 8061 5920
rect 8117 5864 8190 5920
rect 7850 5778 8190 5864
rect 7850 5722 7919 5778
rect 7975 5722 8061 5778
rect 8117 5722 8190 5778
rect 7850 5636 8190 5722
rect 7850 5580 7919 5636
rect 7975 5580 8061 5636
rect 8117 5580 8190 5636
rect 7850 5494 8190 5580
rect 7850 5438 7919 5494
rect 7975 5438 8061 5494
rect 8117 5438 8190 5494
rect 7850 5352 8190 5438
rect 7850 5296 7919 5352
rect 7975 5296 8061 5352
rect 8117 5296 8190 5352
rect 7850 5210 8190 5296
rect 7850 5154 7919 5210
rect 7975 5154 8061 5210
rect 8117 5154 8190 5210
rect 7850 5068 8190 5154
rect 7850 5012 7919 5068
rect 7975 5012 8061 5068
rect 8117 5012 8190 5068
rect 7850 4926 8190 5012
rect 7850 4870 7919 4926
rect 7975 4870 8061 4926
rect 8117 4870 8190 4926
rect 7850 4784 8190 4870
rect 7850 4728 7919 4784
rect 7975 4728 8061 4784
rect 8117 4728 8190 4784
rect 7850 4642 8190 4728
rect 7850 4586 7919 4642
rect 7975 4586 8061 4642
rect 8117 4586 8190 4642
rect 7850 4500 8190 4586
rect 7850 4444 7919 4500
rect 7975 4444 8061 4500
rect 8117 4444 8190 4500
rect 7850 4358 8190 4444
rect 7850 4302 7919 4358
rect 7975 4302 8061 4358
rect 8117 4302 8190 4358
rect 7850 4216 8190 4302
rect 7850 4160 7919 4216
rect 7975 4160 8061 4216
rect 8117 4160 8190 4216
rect 7850 4074 8190 4160
rect 7850 4018 7919 4074
rect 7975 4018 8061 4074
rect 8117 4018 8190 4074
rect 7850 3932 8190 4018
rect 7850 3876 7919 3932
rect 7975 3876 8061 3932
rect 8117 3876 8190 3932
rect 7850 3790 8190 3876
rect 7850 3734 7919 3790
rect 7975 3734 8061 3790
rect 8117 3734 8190 3790
rect 7850 3648 8190 3734
rect 7850 3592 7919 3648
rect 7975 3592 8061 3648
rect 8117 3592 8190 3648
rect 7850 3506 8190 3592
rect 7850 3450 7919 3506
rect 7975 3450 8061 3506
rect 8117 3450 8190 3506
rect 7850 3364 8190 3450
rect 7850 3308 7919 3364
rect 7975 3308 8061 3364
rect 8117 3308 8190 3364
rect 7850 3222 8190 3308
rect 7850 3166 7919 3222
rect 7975 3166 8061 3222
rect 8117 3166 8190 3222
rect 7850 3080 8190 3166
rect 7850 3024 7919 3080
rect 7975 3024 8061 3080
rect 8117 3024 8190 3080
rect 7850 2938 8190 3024
rect 7850 2882 7919 2938
rect 7975 2882 8061 2938
rect 8117 2882 8190 2938
rect 7850 2796 8190 2882
rect 7850 2740 7919 2796
rect 7975 2740 8061 2796
rect 8117 2740 8190 2796
rect 7850 2654 8190 2740
rect 7850 2598 7919 2654
rect 7975 2598 8061 2654
rect 8117 2598 8190 2654
rect 7850 2512 8190 2598
rect 7850 2456 7919 2512
rect 7975 2456 8061 2512
rect 8117 2456 8190 2512
rect 7850 2370 8190 2456
rect 7850 2314 7919 2370
rect 7975 2314 8061 2370
rect 8117 2314 8190 2370
rect 7850 2228 8190 2314
rect 7850 2172 7919 2228
rect 7975 2172 8061 2228
rect 8117 2172 8190 2228
rect 7850 2086 8190 2172
rect 7850 2030 7919 2086
rect 7975 2030 8061 2086
rect 8117 2030 8190 2086
rect 7850 1944 8190 2030
rect 7850 1888 7919 1944
rect 7975 1888 8061 1944
rect 8117 1888 8190 1944
rect 7850 1802 8190 1888
rect 7850 1746 7919 1802
rect 7975 1746 8061 1802
rect 8117 1746 8190 1802
rect 7850 1660 8190 1746
rect 7850 1604 7919 1660
rect 7975 1604 8061 1660
rect 8117 1604 8190 1660
rect 7850 1518 8190 1604
rect 7850 1462 7919 1518
rect 7975 1462 8061 1518
rect 8117 1462 8190 1518
rect 7850 1376 8190 1462
rect 7850 1320 7919 1376
rect 7975 1320 8061 1376
rect 8117 1320 8190 1376
rect 7850 1234 8190 1320
rect 7850 1178 7919 1234
rect 7975 1178 8061 1234
rect 8117 1178 8190 1234
rect 7850 1092 8190 1178
rect 7850 1036 7919 1092
rect 7975 1036 8061 1092
rect 8117 1036 8190 1092
rect 7850 950 8190 1036
rect 7850 894 7919 950
rect 7975 894 8061 950
rect 8117 894 8190 950
rect 7850 808 8190 894
rect 7850 752 7919 808
rect 7975 752 8061 808
rect 8117 752 8190 808
rect 7850 666 8190 752
rect 7850 610 7919 666
rect 7975 610 8061 666
rect 8117 610 8190 666
rect 7850 524 8190 610
rect 7850 468 7919 524
rect 7975 468 8061 524
rect 8117 468 8190 524
rect 7850 458 8190 468
rect 8390 12310 8730 12320
rect 8390 12254 8462 12310
rect 8518 12254 8604 12310
rect 8660 12254 8730 12310
rect 8390 12168 8730 12254
rect 8390 12112 8462 12168
rect 8518 12112 8604 12168
rect 8660 12112 8730 12168
rect 8390 12026 8730 12112
rect 8390 11970 8462 12026
rect 8518 11970 8604 12026
rect 8660 11970 8730 12026
rect 8390 11884 8730 11970
rect 8390 11828 8462 11884
rect 8518 11828 8604 11884
rect 8660 11828 8730 11884
rect 8390 11742 8730 11828
rect 8390 11686 8462 11742
rect 8518 11686 8604 11742
rect 8660 11686 8730 11742
rect 8390 11600 8730 11686
rect 8390 11544 8462 11600
rect 8518 11544 8604 11600
rect 8660 11544 8730 11600
rect 8390 11458 8730 11544
rect 8390 11402 8462 11458
rect 8518 11402 8604 11458
rect 8660 11402 8730 11458
rect 8390 11316 8730 11402
rect 8390 11260 8462 11316
rect 8518 11260 8604 11316
rect 8660 11260 8730 11316
rect 8390 11174 8730 11260
rect 8390 11118 8462 11174
rect 8518 11118 8604 11174
rect 8660 11118 8730 11174
rect 8390 11032 8730 11118
rect 8390 10976 8462 11032
rect 8518 10976 8604 11032
rect 8660 10976 8730 11032
rect 8390 10890 8730 10976
rect 8390 10834 8462 10890
rect 8518 10834 8604 10890
rect 8660 10834 8730 10890
rect 8390 10748 8730 10834
rect 8390 10692 8462 10748
rect 8518 10692 8604 10748
rect 8660 10692 8730 10748
rect 8390 10606 8730 10692
rect 8390 10550 8462 10606
rect 8518 10550 8604 10606
rect 8660 10550 8730 10606
rect 8390 10464 8730 10550
rect 8390 10408 8462 10464
rect 8518 10408 8604 10464
rect 8660 10408 8730 10464
rect 8390 10322 8730 10408
rect 8390 10266 8462 10322
rect 8518 10266 8604 10322
rect 8660 10266 8730 10322
rect 8390 10180 8730 10266
rect 8390 10124 8462 10180
rect 8518 10124 8604 10180
rect 8660 10124 8730 10180
rect 8390 10038 8730 10124
rect 8390 9982 8462 10038
rect 8518 9982 8604 10038
rect 8660 9982 8730 10038
rect 8390 9896 8730 9982
rect 8390 9840 8462 9896
rect 8518 9840 8604 9896
rect 8660 9840 8730 9896
rect 8390 9754 8730 9840
rect 8390 9698 8462 9754
rect 8518 9698 8604 9754
rect 8660 9698 8730 9754
rect 8390 9612 8730 9698
rect 8390 9556 8462 9612
rect 8518 9556 8604 9612
rect 8660 9556 8730 9612
rect 8390 9470 8730 9556
rect 8390 9414 8462 9470
rect 8518 9414 8604 9470
rect 8660 9414 8730 9470
rect 8390 9328 8730 9414
rect 8390 9272 8462 9328
rect 8518 9272 8604 9328
rect 8660 9272 8730 9328
rect 8390 9186 8730 9272
rect 8390 9130 8462 9186
rect 8518 9130 8604 9186
rect 8660 9130 8730 9186
rect 8390 9044 8730 9130
rect 8390 8988 8462 9044
rect 8518 8988 8604 9044
rect 8660 8988 8730 9044
rect 8390 8902 8730 8988
rect 8390 8846 8462 8902
rect 8518 8846 8604 8902
rect 8660 8846 8730 8902
rect 8390 8760 8730 8846
rect 8390 8704 8462 8760
rect 8518 8704 8604 8760
rect 8660 8704 8730 8760
rect 8390 8618 8730 8704
rect 8390 8562 8462 8618
rect 8518 8562 8604 8618
rect 8660 8562 8730 8618
rect 8390 8476 8730 8562
rect 8390 8420 8462 8476
rect 8518 8420 8604 8476
rect 8660 8420 8730 8476
rect 8390 8334 8730 8420
rect 8390 8278 8462 8334
rect 8518 8278 8604 8334
rect 8660 8278 8730 8334
rect 8390 8192 8730 8278
rect 8390 8136 8462 8192
rect 8518 8136 8604 8192
rect 8660 8136 8730 8192
rect 8390 8050 8730 8136
rect 8390 7994 8462 8050
rect 8518 7994 8604 8050
rect 8660 7994 8730 8050
rect 8390 7908 8730 7994
rect 8390 7852 8462 7908
rect 8518 7852 8604 7908
rect 8660 7852 8730 7908
rect 8390 7766 8730 7852
rect 8390 7710 8462 7766
rect 8518 7710 8604 7766
rect 8660 7710 8730 7766
rect 8390 7624 8730 7710
rect 8390 7568 8462 7624
rect 8518 7568 8604 7624
rect 8660 7568 8730 7624
rect 8390 7482 8730 7568
rect 8390 7426 8462 7482
rect 8518 7426 8604 7482
rect 8660 7426 8730 7482
rect 8390 7340 8730 7426
rect 8390 7284 8462 7340
rect 8518 7284 8604 7340
rect 8660 7284 8730 7340
rect 8390 7198 8730 7284
rect 8390 7142 8462 7198
rect 8518 7142 8604 7198
rect 8660 7142 8730 7198
rect 8390 7056 8730 7142
rect 8390 7000 8462 7056
rect 8518 7000 8604 7056
rect 8660 7000 8730 7056
rect 8390 6914 8730 7000
rect 8390 6858 8462 6914
rect 8518 6858 8604 6914
rect 8660 6858 8730 6914
rect 8390 6772 8730 6858
rect 8390 6716 8462 6772
rect 8518 6716 8604 6772
rect 8660 6716 8730 6772
rect 8390 6630 8730 6716
rect 8390 6574 8462 6630
rect 8518 6574 8604 6630
rect 8660 6574 8730 6630
rect 8390 6488 8730 6574
rect 8390 6432 8462 6488
rect 8518 6432 8604 6488
rect 8660 6432 8730 6488
rect 8390 6346 8730 6432
rect 8390 6290 8462 6346
rect 8518 6290 8604 6346
rect 8660 6290 8730 6346
rect 8390 6204 8730 6290
rect 8390 6148 8462 6204
rect 8518 6148 8604 6204
rect 8660 6148 8730 6204
rect 8390 6062 8730 6148
rect 8390 6006 8462 6062
rect 8518 6006 8604 6062
rect 8660 6006 8730 6062
rect 8390 5920 8730 6006
rect 8390 5864 8462 5920
rect 8518 5864 8604 5920
rect 8660 5864 8730 5920
rect 8390 5778 8730 5864
rect 8390 5722 8462 5778
rect 8518 5722 8604 5778
rect 8660 5722 8730 5778
rect 8390 5636 8730 5722
rect 8390 5580 8462 5636
rect 8518 5580 8604 5636
rect 8660 5580 8730 5636
rect 8390 5494 8730 5580
rect 8390 5438 8462 5494
rect 8518 5438 8604 5494
rect 8660 5438 8730 5494
rect 8390 5352 8730 5438
rect 8390 5296 8462 5352
rect 8518 5296 8604 5352
rect 8660 5296 8730 5352
rect 8390 5210 8730 5296
rect 8390 5154 8462 5210
rect 8518 5154 8604 5210
rect 8660 5154 8730 5210
rect 8390 5068 8730 5154
rect 8390 5012 8462 5068
rect 8518 5012 8604 5068
rect 8660 5012 8730 5068
rect 8390 4926 8730 5012
rect 8390 4870 8462 4926
rect 8518 4870 8604 4926
rect 8660 4870 8730 4926
rect 8390 4784 8730 4870
rect 8390 4728 8462 4784
rect 8518 4728 8604 4784
rect 8660 4728 8730 4784
rect 8390 4642 8730 4728
rect 8390 4586 8462 4642
rect 8518 4586 8604 4642
rect 8660 4586 8730 4642
rect 8390 4500 8730 4586
rect 8390 4444 8462 4500
rect 8518 4444 8604 4500
rect 8660 4444 8730 4500
rect 8390 4358 8730 4444
rect 8390 4302 8462 4358
rect 8518 4302 8604 4358
rect 8660 4302 8730 4358
rect 8390 4216 8730 4302
rect 8390 4160 8462 4216
rect 8518 4160 8604 4216
rect 8660 4160 8730 4216
rect 8390 4074 8730 4160
rect 8390 4018 8462 4074
rect 8518 4018 8604 4074
rect 8660 4018 8730 4074
rect 8390 3932 8730 4018
rect 8390 3876 8462 3932
rect 8518 3876 8604 3932
rect 8660 3876 8730 3932
rect 8390 3790 8730 3876
rect 8390 3734 8462 3790
rect 8518 3734 8604 3790
rect 8660 3734 8730 3790
rect 8390 3648 8730 3734
rect 8390 3592 8462 3648
rect 8518 3592 8604 3648
rect 8660 3592 8730 3648
rect 8390 3506 8730 3592
rect 8390 3450 8462 3506
rect 8518 3450 8604 3506
rect 8660 3450 8730 3506
rect 8390 3364 8730 3450
rect 8390 3308 8462 3364
rect 8518 3308 8604 3364
rect 8660 3308 8730 3364
rect 8390 3222 8730 3308
rect 8390 3166 8462 3222
rect 8518 3166 8604 3222
rect 8660 3166 8730 3222
rect 8390 3080 8730 3166
rect 8390 3024 8462 3080
rect 8518 3024 8604 3080
rect 8660 3024 8730 3080
rect 8390 2938 8730 3024
rect 8390 2882 8462 2938
rect 8518 2882 8604 2938
rect 8660 2882 8730 2938
rect 8390 2796 8730 2882
rect 8390 2740 8462 2796
rect 8518 2740 8604 2796
rect 8660 2740 8730 2796
rect 8390 2654 8730 2740
rect 8390 2598 8462 2654
rect 8518 2598 8604 2654
rect 8660 2598 8730 2654
rect 8390 2512 8730 2598
rect 8390 2456 8462 2512
rect 8518 2456 8604 2512
rect 8660 2456 8730 2512
rect 8390 2370 8730 2456
rect 8390 2314 8462 2370
rect 8518 2314 8604 2370
rect 8660 2314 8730 2370
rect 8390 2228 8730 2314
rect 8390 2172 8462 2228
rect 8518 2172 8604 2228
rect 8660 2172 8730 2228
rect 8390 2086 8730 2172
rect 8390 2030 8462 2086
rect 8518 2030 8604 2086
rect 8660 2030 8730 2086
rect 8390 1944 8730 2030
rect 8390 1888 8462 1944
rect 8518 1888 8604 1944
rect 8660 1888 8730 1944
rect 8390 1802 8730 1888
rect 8390 1746 8462 1802
rect 8518 1746 8604 1802
rect 8660 1746 8730 1802
rect 8390 1660 8730 1746
rect 8390 1604 8462 1660
rect 8518 1604 8604 1660
rect 8660 1604 8730 1660
rect 8390 1518 8730 1604
rect 8390 1462 8462 1518
rect 8518 1462 8604 1518
rect 8660 1462 8730 1518
rect 8390 1376 8730 1462
rect 8390 1320 8462 1376
rect 8518 1320 8604 1376
rect 8660 1320 8730 1376
rect 8390 1234 8730 1320
rect 8390 1178 8462 1234
rect 8518 1178 8604 1234
rect 8660 1178 8730 1234
rect 8390 1092 8730 1178
rect 8390 1036 8462 1092
rect 8518 1036 8604 1092
rect 8660 1036 8730 1092
rect 8390 950 8730 1036
rect 8390 894 8462 950
rect 8518 894 8604 950
rect 8660 894 8730 950
rect 8390 808 8730 894
rect 8390 752 8462 808
rect 8518 752 8604 808
rect 8660 752 8730 808
rect 8390 666 8730 752
rect 8390 610 8462 666
rect 8518 610 8604 666
rect 8660 610 8730 666
rect 8390 524 8730 610
rect 8390 468 8462 524
rect 8518 468 8604 524
rect 8660 468 8730 524
rect 8390 458 8730 468
rect 8930 12310 9270 12320
rect 8930 12254 9004 12310
rect 9060 12254 9146 12310
rect 9202 12254 9270 12310
rect 8930 12168 9270 12254
rect 8930 12112 9004 12168
rect 9060 12112 9146 12168
rect 9202 12112 9270 12168
rect 8930 12026 9270 12112
rect 8930 11970 9004 12026
rect 9060 11970 9146 12026
rect 9202 11970 9270 12026
rect 8930 11884 9270 11970
rect 8930 11828 9004 11884
rect 9060 11828 9146 11884
rect 9202 11828 9270 11884
rect 8930 11742 9270 11828
rect 8930 11686 9004 11742
rect 9060 11686 9146 11742
rect 9202 11686 9270 11742
rect 8930 11600 9270 11686
rect 8930 11544 9004 11600
rect 9060 11544 9146 11600
rect 9202 11544 9270 11600
rect 8930 11458 9270 11544
rect 8930 11402 9004 11458
rect 9060 11402 9146 11458
rect 9202 11402 9270 11458
rect 8930 11316 9270 11402
rect 8930 11260 9004 11316
rect 9060 11260 9146 11316
rect 9202 11260 9270 11316
rect 8930 11174 9270 11260
rect 8930 11118 9004 11174
rect 9060 11118 9146 11174
rect 9202 11118 9270 11174
rect 8930 11032 9270 11118
rect 8930 10976 9004 11032
rect 9060 10976 9146 11032
rect 9202 10976 9270 11032
rect 8930 10890 9270 10976
rect 8930 10834 9004 10890
rect 9060 10834 9146 10890
rect 9202 10834 9270 10890
rect 8930 10748 9270 10834
rect 8930 10692 9004 10748
rect 9060 10692 9146 10748
rect 9202 10692 9270 10748
rect 8930 10606 9270 10692
rect 8930 10550 9004 10606
rect 9060 10550 9146 10606
rect 9202 10550 9270 10606
rect 8930 10464 9270 10550
rect 8930 10408 9004 10464
rect 9060 10408 9146 10464
rect 9202 10408 9270 10464
rect 8930 10322 9270 10408
rect 8930 10266 9004 10322
rect 9060 10266 9146 10322
rect 9202 10266 9270 10322
rect 8930 10180 9270 10266
rect 8930 10124 9004 10180
rect 9060 10124 9146 10180
rect 9202 10124 9270 10180
rect 8930 10038 9270 10124
rect 8930 9982 9004 10038
rect 9060 9982 9146 10038
rect 9202 9982 9270 10038
rect 8930 9896 9270 9982
rect 8930 9840 9004 9896
rect 9060 9840 9146 9896
rect 9202 9840 9270 9896
rect 8930 9754 9270 9840
rect 8930 9698 9004 9754
rect 9060 9698 9146 9754
rect 9202 9698 9270 9754
rect 8930 9612 9270 9698
rect 8930 9556 9004 9612
rect 9060 9556 9146 9612
rect 9202 9556 9270 9612
rect 8930 9470 9270 9556
rect 8930 9414 9004 9470
rect 9060 9414 9146 9470
rect 9202 9414 9270 9470
rect 8930 9328 9270 9414
rect 8930 9272 9004 9328
rect 9060 9272 9146 9328
rect 9202 9272 9270 9328
rect 8930 9186 9270 9272
rect 8930 9130 9004 9186
rect 9060 9130 9146 9186
rect 9202 9130 9270 9186
rect 8930 9044 9270 9130
rect 8930 8988 9004 9044
rect 9060 8988 9146 9044
rect 9202 8988 9270 9044
rect 8930 8902 9270 8988
rect 8930 8846 9004 8902
rect 9060 8846 9146 8902
rect 9202 8846 9270 8902
rect 8930 8760 9270 8846
rect 8930 8704 9004 8760
rect 9060 8704 9146 8760
rect 9202 8704 9270 8760
rect 8930 8618 9270 8704
rect 8930 8562 9004 8618
rect 9060 8562 9146 8618
rect 9202 8562 9270 8618
rect 8930 8476 9270 8562
rect 8930 8420 9004 8476
rect 9060 8420 9146 8476
rect 9202 8420 9270 8476
rect 8930 8334 9270 8420
rect 8930 8278 9004 8334
rect 9060 8278 9146 8334
rect 9202 8278 9270 8334
rect 8930 8192 9270 8278
rect 8930 8136 9004 8192
rect 9060 8136 9146 8192
rect 9202 8136 9270 8192
rect 8930 8050 9270 8136
rect 8930 7994 9004 8050
rect 9060 7994 9146 8050
rect 9202 7994 9270 8050
rect 8930 7908 9270 7994
rect 8930 7852 9004 7908
rect 9060 7852 9146 7908
rect 9202 7852 9270 7908
rect 8930 7766 9270 7852
rect 8930 7710 9004 7766
rect 9060 7710 9146 7766
rect 9202 7710 9270 7766
rect 8930 7624 9270 7710
rect 8930 7568 9004 7624
rect 9060 7568 9146 7624
rect 9202 7568 9270 7624
rect 8930 7482 9270 7568
rect 8930 7426 9004 7482
rect 9060 7426 9146 7482
rect 9202 7426 9270 7482
rect 8930 7340 9270 7426
rect 8930 7284 9004 7340
rect 9060 7284 9146 7340
rect 9202 7284 9270 7340
rect 8930 7198 9270 7284
rect 8930 7142 9004 7198
rect 9060 7142 9146 7198
rect 9202 7142 9270 7198
rect 8930 7056 9270 7142
rect 8930 7000 9004 7056
rect 9060 7000 9146 7056
rect 9202 7000 9270 7056
rect 8930 6914 9270 7000
rect 8930 6858 9004 6914
rect 9060 6858 9146 6914
rect 9202 6858 9270 6914
rect 8930 6772 9270 6858
rect 8930 6716 9004 6772
rect 9060 6716 9146 6772
rect 9202 6716 9270 6772
rect 8930 6630 9270 6716
rect 8930 6574 9004 6630
rect 9060 6574 9146 6630
rect 9202 6574 9270 6630
rect 8930 6488 9270 6574
rect 8930 6432 9004 6488
rect 9060 6432 9146 6488
rect 9202 6432 9270 6488
rect 8930 6346 9270 6432
rect 8930 6290 9004 6346
rect 9060 6290 9146 6346
rect 9202 6290 9270 6346
rect 8930 6204 9270 6290
rect 8930 6148 9004 6204
rect 9060 6148 9146 6204
rect 9202 6148 9270 6204
rect 8930 6062 9270 6148
rect 8930 6006 9004 6062
rect 9060 6006 9146 6062
rect 9202 6006 9270 6062
rect 8930 5920 9270 6006
rect 8930 5864 9004 5920
rect 9060 5864 9146 5920
rect 9202 5864 9270 5920
rect 8930 5778 9270 5864
rect 8930 5722 9004 5778
rect 9060 5722 9146 5778
rect 9202 5722 9270 5778
rect 8930 5636 9270 5722
rect 8930 5580 9004 5636
rect 9060 5580 9146 5636
rect 9202 5580 9270 5636
rect 8930 5494 9270 5580
rect 8930 5438 9004 5494
rect 9060 5438 9146 5494
rect 9202 5438 9270 5494
rect 8930 5352 9270 5438
rect 8930 5296 9004 5352
rect 9060 5296 9146 5352
rect 9202 5296 9270 5352
rect 8930 5210 9270 5296
rect 8930 5154 9004 5210
rect 9060 5154 9146 5210
rect 9202 5154 9270 5210
rect 8930 5068 9270 5154
rect 8930 5012 9004 5068
rect 9060 5012 9146 5068
rect 9202 5012 9270 5068
rect 8930 4926 9270 5012
rect 8930 4870 9004 4926
rect 9060 4870 9146 4926
rect 9202 4870 9270 4926
rect 8930 4784 9270 4870
rect 8930 4728 9004 4784
rect 9060 4728 9146 4784
rect 9202 4728 9270 4784
rect 8930 4642 9270 4728
rect 8930 4586 9004 4642
rect 9060 4586 9146 4642
rect 9202 4586 9270 4642
rect 8930 4500 9270 4586
rect 8930 4444 9004 4500
rect 9060 4444 9146 4500
rect 9202 4444 9270 4500
rect 8930 4358 9270 4444
rect 8930 4302 9004 4358
rect 9060 4302 9146 4358
rect 9202 4302 9270 4358
rect 8930 4216 9270 4302
rect 8930 4160 9004 4216
rect 9060 4160 9146 4216
rect 9202 4160 9270 4216
rect 8930 4074 9270 4160
rect 8930 4018 9004 4074
rect 9060 4018 9146 4074
rect 9202 4018 9270 4074
rect 8930 3932 9270 4018
rect 8930 3876 9004 3932
rect 9060 3876 9146 3932
rect 9202 3876 9270 3932
rect 8930 3790 9270 3876
rect 8930 3734 9004 3790
rect 9060 3734 9146 3790
rect 9202 3734 9270 3790
rect 8930 3648 9270 3734
rect 8930 3592 9004 3648
rect 9060 3592 9146 3648
rect 9202 3592 9270 3648
rect 8930 3506 9270 3592
rect 8930 3450 9004 3506
rect 9060 3450 9146 3506
rect 9202 3450 9270 3506
rect 8930 3364 9270 3450
rect 8930 3308 9004 3364
rect 9060 3308 9146 3364
rect 9202 3308 9270 3364
rect 8930 3222 9270 3308
rect 8930 3166 9004 3222
rect 9060 3166 9146 3222
rect 9202 3166 9270 3222
rect 8930 3080 9270 3166
rect 8930 3024 9004 3080
rect 9060 3024 9146 3080
rect 9202 3024 9270 3080
rect 8930 2938 9270 3024
rect 8930 2882 9004 2938
rect 9060 2882 9146 2938
rect 9202 2882 9270 2938
rect 8930 2796 9270 2882
rect 8930 2740 9004 2796
rect 9060 2740 9146 2796
rect 9202 2740 9270 2796
rect 8930 2654 9270 2740
rect 8930 2598 9004 2654
rect 9060 2598 9146 2654
rect 9202 2598 9270 2654
rect 8930 2512 9270 2598
rect 8930 2456 9004 2512
rect 9060 2456 9146 2512
rect 9202 2456 9270 2512
rect 8930 2370 9270 2456
rect 8930 2314 9004 2370
rect 9060 2314 9146 2370
rect 9202 2314 9270 2370
rect 8930 2228 9270 2314
rect 8930 2172 9004 2228
rect 9060 2172 9146 2228
rect 9202 2172 9270 2228
rect 8930 2086 9270 2172
rect 8930 2030 9004 2086
rect 9060 2030 9146 2086
rect 9202 2030 9270 2086
rect 8930 1944 9270 2030
rect 8930 1888 9004 1944
rect 9060 1888 9146 1944
rect 9202 1888 9270 1944
rect 8930 1802 9270 1888
rect 8930 1746 9004 1802
rect 9060 1746 9146 1802
rect 9202 1746 9270 1802
rect 8930 1660 9270 1746
rect 8930 1604 9004 1660
rect 9060 1604 9146 1660
rect 9202 1604 9270 1660
rect 8930 1518 9270 1604
rect 8930 1462 9004 1518
rect 9060 1462 9146 1518
rect 9202 1462 9270 1518
rect 8930 1376 9270 1462
rect 8930 1320 9004 1376
rect 9060 1320 9146 1376
rect 9202 1320 9270 1376
rect 8930 1234 9270 1320
rect 8930 1178 9004 1234
rect 9060 1178 9146 1234
rect 9202 1178 9270 1234
rect 8930 1092 9270 1178
rect 8930 1036 9004 1092
rect 9060 1036 9146 1092
rect 9202 1036 9270 1092
rect 8930 950 9270 1036
rect 8930 894 9004 950
rect 9060 894 9146 950
rect 9202 894 9270 950
rect 8930 808 9270 894
rect 8930 752 9004 808
rect 9060 752 9146 808
rect 9202 752 9270 808
rect 8930 666 9270 752
rect 8930 610 9004 666
rect 9060 610 9146 666
rect 9202 610 9270 666
rect 8930 524 9270 610
rect 8930 468 9004 524
rect 9060 468 9146 524
rect 9202 468 9270 524
rect 8930 458 9270 468
rect 9470 12310 9810 12320
rect 9470 12254 9547 12310
rect 9603 12254 9689 12310
rect 9745 12254 9810 12310
rect 9470 12168 9810 12254
rect 9470 12112 9547 12168
rect 9603 12112 9689 12168
rect 9745 12112 9810 12168
rect 9470 12026 9810 12112
rect 9470 11970 9547 12026
rect 9603 11970 9689 12026
rect 9745 11970 9810 12026
rect 9470 11884 9810 11970
rect 9470 11828 9547 11884
rect 9603 11828 9689 11884
rect 9745 11828 9810 11884
rect 9470 11742 9810 11828
rect 9470 11686 9547 11742
rect 9603 11686 9689 11742
rect 9745 11686 9810 11742
rect 9470 11600 9810 11686
rect 9470 11544 9547 11600
rect 9603 11544 9689 11600
rect 9745 11544 9810 11600
rect 9470 11458 9810 11544
rect 9470 11402 9547 11458
rect 9603 11402 9689 11458
rect 9745 11402 9810 11458
rect 9470 11316 9810 11402
rect 9470 11260 9547 11316
rect 9603 11260 9689 11316
rect 9745 11260 9810 11316
rect 9470 11174 9810 11260
rect 9470 11118 9547 11174
rect 9603 11118 9689 11174
rect 9745 11118 9810 11174
rect 9470 11032 9810 11118
rect 9470 10976 9547 11032
rect 9603 10976 9689 11032
rect 9745 10976 9810 11032
rect 9470 10890 9810 10976
rect 9470 10834 9547 10890
rect 9603 10834 9689 10890
rect 9745 10834 9810 10890
rect 9470 10748 9810 10834
rect 9470 10692 9547 10748
rect 9603 10692 9689 10748
rect 9745 10692 9810 10748
rect 9470 10606 9810 10692
rect 9470 10550 9547 10606
rect 9603 10550 9689 10606
rect 9745 10550 9810 10606
rect 9470 10464 9810 10550
rect 9470 10408 9547 10464
rect 9603 10408 9689 10464
rect 9745 10408 9810 10464
rect 9470 10322 9810 10408
rect 9470 10266 9547 10322
rect 9603 10266 9689 10322
rect 9745 10266 9810 10322
rect 9470 10180 9810 10266
rect 9470 10124 9547 10180
rect 9603 10124 9689 10180
rect 9745 10124 9810 10180
rect 9470 10038 9810 10124
rect 9470 9982 9547 10038
rect 9603 9982 9689 10038
rect 9745 9982 9810 10038
rect 9470 9896 9810 9982
rect 9470 9840 9547 9896
rect 9603 9840 9689 9896
rect 9745 9840 9810 9896
rect 9470 9754 9810 9840
rect 9470 9698 9547 9754
rect 9603 9698 9689 9754
rect 9745 9698 9810 9754
rect 9470 9612 9810 9698
rect 9470 9556 9547 9612
rect 9603 9556 9689 9612
rect 9745 9556 9810 9612
rect 9470 9470 9810 9556
rect 9470 9414 9547 9470
rect 9603 9414 9689 9470
rect 9745 9414 9810 9470
rect 9470 9328 9810 9414
rect 9470 9272 9547 9328
rect 9603 9272 9689 9328
rect 9745 9272 9810 9328
rect 9470 9186 9810 9272
rect 9470 9130 9547 9186
rect 9603 9130 9689 9186
rect 9745 9130 9810 9186
rect 9470 9044 9810 9130
rect 9470 8988 9547 9044
rect 9603 8988 9689 9044
rect 9745 8988 9810 9044
rect 9470 8902 9810 8988
rect 9470 8846 9547 8902
rect 9603 8846 9689 8902
rect 9745 8846 9810 8902
rect 9470 8760 9810 8846
rect 9470 8704 9547 8760
rect 9603 8704 9689 8760
rect 9745 8704 9810 8760
rect 9470 8618 9810 8704
rect 9470 8562 9547 8618
rect 9603 8562 9689 8618
rect 9745 8562 9810 8618
rect 9470 8476 9810 8562
rect 9470 8420 9547 8476
rect 9603 8420 9689 8476
rect 9745 8420 9810 8476
rect 9470 8334 9810 8420
rect 9470 8278 9547 8334
rect 9603 8278 9689 8334
rect 9745 8278 9810 8334
rect 9470 8192 9810 8278
rect 9470 8136 9547 8192
rect 9603 8136 9689 8192
rect 9745 8136 9810 8192
rect 9470 8050 9810 8136
rect 9470 7994 9547 8050
rect 9603 7994 9689 8050
rect 9745 7994 9810 8050
rect 9470 7908 9810 7994
rect 9470 7852 9547 7908
rect 9603 7852 9689 7908
rect 9745 7852 9810 7908
rect 9470 7766 9810 7852
rect 9470 7710 9547 7766
rect 9603 7710 9689 7766
rect 9745 7710 9810 7766
rect 9470 7624 9810 7710
rect 9470 7568 9547 7624
rect 9603 7568 9689 7624
rect 9745 7568 9810 7624
rect 9470 7482 9810 7568
rect 9470 7426 9547 7482
rect 9603 7426 9689 7482
rect 9745 7426 9810 7482
rect 9470 7340 9810 7426
rect 9470 7284 9547 7340
rect 9603 7284 9689 7340
rect 9745 7284 9810 7340
rect 9470 7198 9810 7284
rect 9470 7142 9547 7198
rect 9603 7142 9689 7198
rect 9745 7142 9810 7198
rect 9470 7056 9810 7142
rect 9470 7000 9547 7056
rect 9603 7000 9689 7056
rect 9745 7000 9810 7056
rect 9470 6914 9810 7000
rect 9470 6858 9547 6914
rect 9603 6858 9689 6914
rect 9745 6858 9810 6914
rect 9470 6772 9810 6858
rect 9470 6716 9547 6772
rect 9603 6716 9689 6772
rect 9745 6716 9810 6772
rect 9470 6630 9810 6716
rect 9470 6574 9547 6630
rect 9603 6574 9689 6630
rect 9745 6574 9810 6630
rect 9470 6488 9810 6574
rect 9470 6432 9547 6488
rect 9603 6432 9689 6488
rect 9745 6432 9810 6488
rect 9470 6346 9810 6432
rect 9470 6290 9547 6346
rect 9603 6290 9689 6346
rect 9745 6290 9810 6346
rect 9470 6204 9810 6290
rect 9470 6148 9547 6204
rect 9603 6148 9689 6204
rect 9745 6148 9810 6204
rect 9470 6062 9810 6148
rect 9470 6006 9547 6062
rect 9603 6006 9689 6062
rect 9745 6006 9810 6062
rect 9470 5920 9810 6006
rect 9470 5864 9547 5920
rect 9603 5864 9689 5920
rect 9745 5864 9810 5920
rect 9470 5778 9810 5864
rect 9470 5722 9547 5778
rect 9603 5722 9689 5778
rect 9745 5722 9810 5778
rect 9470 5636 9810 5722
rect 9470 5580 9547 5636
rect 9603 5580 9689 5636
rect 9745 5580 9810 5636
rect 9470 5494 9810 5580
rect 9470 5438 9547 5494
rect 9603 5438 9689 5494
rect 9745 5438 9810 5494
rect 9470 5352 9810 5438
rect 9470 5296 9547 5352
rect 9603 5296 9689 5352
rect 9745 5296 9810 5352
rect 9470 5210 9810 5296
rect 9470 5154 9547 5210
rect 9603 5154 9689 5210
rect 9745 5154 9810 5210
rect 9470 5068 9810 5154
rect 9470 5012 9547 5068
rect 9603 5012 9689 5068
rect 9745 5012 9810 5068
rect 9470 4926 9810 5012
rect 9470 4870 9547 4926
rect 9603 4870 9689 4926
rect 9745 4870 9810 4926
rect 9470 4784 9810 4870
rect 9470 4728 9547 4784
rect 9603 4728 9689 4784
rect 9745 4728 9810 4784
rect 9470 4642 9810 4728
rect 9470 4586 9547 4642
rect 9603 4586 9689 4642
rect 9745 4586 9810 4642
rect 9470 4500 9810 4586
rect 9470 4444 9547 4500
rect 9603 4444 9689 4500
rect 9745 4444 9810 4500
rect 9470 4358 9810 4444
rect 9470 4302 9547 4358
rect 9603 4302 9689 4358
rect 9745 4302 9810 4358
rect 9470 4216 9810 4302
rect 9470 4160 9547 4216
rect 9603 4160 9689 4216
rect 9745 4160 9810 4216
rect 9470 4074 9810 4160
rect 9470 4018 9547 4074
rect 9603 4018 9689 4074
rect 9745 4018 9810 4074
rect 9470 3932 9810 4018
rect 9470 3876 9547 3932
rect 9603 3876 9689 3932
rect 9745 3876 9810 3932
rect 9470 3790 9810 3876
rect 9470 3734 9547 3790
rect 9603 3734 9689 3790
rect 9745 3734 9810 3790
rect 9470 3648 9810 3734
rect 9470 3592 9547 3648
rect 9603 3592 9689 3648
rect 9745 3592 9810 3648
rect 9470 3506 9810 3592
rect 9470 3450 9547 3506
rect 9603 3450 9689 3506
rect 9745 3450 9810 3506
rect 9470 3364 9810 3450
rect 9470 3308 9547 3364
rect 9603 3308 9689 3364
rect 9745 3308 9810 3364
rect 9470 3222 9810 3308
rect 9470 3166 9547 3222
rect 9603 3166 9689 3222
rect 9745 3166 9810 3222
rect 9470 3080 9810 3166
rect 9470 3024 9547 3080
rect 9603 3024 9689 3080
rect 9745 3024 9810 3080
rect 9470 2938 9810 3024
rect 9470 2882 9547 2938
rect 9603 2882 9689 2938
rect 9745 2882 9810 2938
rect 9470 2796 9810 2882
rect 9470 2740 9547 2796
rect 9603 2740 9689 2796
rect 9745 2740 9810 2796
rect 9470 2654 9810 2740
rect 9470 2598 9547 2654
rect 9603 2598 9689 2654
rect 9745 2598 9810 2654
rect 9470 2512 9810 2598
rect 9470 2456 9547 2512
rect 9603 2456 9689 2512
rect 9745 2456 9810 2512
rect 9470 2370 9810 2456
rect 9470 2314 9547 2370
rect 9603 2314 9689 2370
rect 9745 2314 9810 2370
rect 9470 2228 9810 2314
rect 9470 2172 9547 2228
rect 9603 2172 9689 2228
rect 9745 2172 9810 2228
rect 9470 2086 9810 2172
rect 9470 2030 9547 2086
rect 9603 2030 9689 2086
rect 9745 2030 9810 2086
rect 9470 1944 9810 2030
rect 9470 1888 9547 1944
rect 9603 1888 9689 1944
rect 9745 1888 9810 1944
rect 9470 1802 9810 1888
rect 9470 1746 9547 1802
rect 9603 1746 9689 1802
rect 9745 1746 9810 1802
rect 9470 1660 9810 1746
rect 9470 1604 9547 1660
rect 9603 1604 9689 1660
rect 9745 1604 9810 1660
rect 9470 1518 9810 1604
rect 9470 1462 9547 1518
rect 9603 1462 9689 1518
rect 9745 1462 9810 1518
rect 9470 1376 9810 1462
rect 9470 1320 9547 1376
rect 9603 1320 9689 1376
rect 9745 1320 9810 1376
rect 9470 1234 9810 1320
rect 9470 1178 9547 1234
rect 9603 1178 9689 1234
rect 9745 1178 9810 1234
rect 9470 1092 9810 1178
rect 9470 1036 9547 1092
rect 9603 1036 9689 1092
rect 9745 1036 9810 1092
rect 9470 950 9810 1036
rect 9470 894 9547 950
rect 9603 894 9689 950
rect 9745 894 9810 950
rect 9470 808 9810 894
rect 9470 752 9547 808
rect 9603 752 9689 808
rect 9745 752 9810 808
rect 9470 666 9810 752
rect 9470 610 9547 666
rect 9603 610 9689 666
rect 9745 610 9810 666
rect 9470 524 9810 610
rect 9470 468 9547 524
rect 9603 468 9689 524
rect 9745 468 9810 524
rect 9470 458 9810 468
rect 10010 12310 10350 12320
rect 10010 12254 10081 12310
rect 10137 12254 10223 12310
rect 10279 12254 10350 12310
rect 10010 12168 10350 12254
rect 10010 12112 10081 12168
rect 10137 12112 10223 12168
rect 10279 12112 10350 12168
rect 10010 12026 10350 12112
rect 10010 11970 10081 12026
rect 10137 11970 10223 12026
rect 10279 11970 10350 12026
rect 10010 11884 10350 11970
rect 10010 11828 10081 11884
rect 10137 11828 10223 11884
rect 10279 11828 10350 11884
rect 10010 11742 10350 11828
rect 10010 11686 10081 11742
rect 10137 11686 10223 11742
rect 10279 11686 10350 11742
rect 10010 11600 10350 11686
rect 10010 11544 10081 11600
rect 10137 11544 10223 11600
rect 10279 11544 10350 11600
rect 10010 11458 10350 11544
rect 10010 11402 10081 11458
rect 10137 11402 10223 11458
rect 10279 11402 10350 11458
rect 10010 11316 10350 11402
rect 10010 11260 10081 11316
rect 10137 11260 10223 11316
rect 10279 11260 10350 11316
rect 10010 11174 10350 11260
rect 10010 11118 10081 11174
rect 10137 11118 10223 11174
rect 10279 11118 10350 11174
rect 10010 11032 10350 11118
rect 10010 10976 10081 11032
rect 10137 10976 10223 11032
rect 10279 10976 10350 11032
rect 10010 10890 10350 10976
rect 10010 10834 10081 10890
rect 10137 10834 10223 10890
rect 10279 10834 10350 10890
rect 10010 10748 10350 10834
rect 10010 10692 10081 10748
rect 10137 10692 10223 10748
rect 10279 10692 10350 10748
rect 10010 10606 10350 10692
rect 10010 10550 10081 10606
rect 10137 10550 10223 10606
rect 10279 10550 10350 10606
rect 10010 10464 10350 10550
rect 10010 10408 10081 10464
rect 10137 10408 10223 10464
rect 10279 10408 10350 10464
rect 10010 10322 10350 10408
rect 10010 10266 10081 10322
rect 10137 10266 10223 10322
rect 10279 10266 10350 10322
rect 10010 10180 10350 10266
rect 10010 10124 10081 10180
rect 10137 10124 10223 10180
rect 10279 10124 10350 10180
rect 10010 10038 10350 10124
rect 10010 9982 10081 10038
rect 10137 9982 10223 10038
rect 10279 9982 10350 10038
rect 10010 9896 10350 9982
rect 10010 9840 10081 9896
rect 10137 9840 10223 9896
rect 10279 9840 10350 9896
rect 10010 9754 10350 9840
rect 10010 9698 10081 9754
rect 10137 9698 10223 9754
rect 10279 9698 10350 9754
rect 10010 9612 10350 9698
rect 10010 9556 10081 9612
rect 10137 9556 10223 9612
rect 10279 9556 10350 9612
rect 10010 9470 10350 9556
rect 10010 9414 10081 9470
rect 10137 9414 10223 9470
rect 10279 9414 10350 9470
rect 10010 9328 10350 9414
rect 10010 9272 10081 9328
rect 10137 9272 10223 9328
rect 10279 9272 10350 9328
rect 10010 9186 10350 9272
rect 10010 9130 10081 9186
rect 10137 9130 10223 9186
rect 10279 9130 10350 9186
rect 10010 9044 10350 9130
rect 10010 8988 10081 9044
rect 10137 8988 10223 9044
rect 10279 8988 10350 9044
rect 10010 8902 10350 8988
rect 10010 8846 10081 8902
rect 10137 8846 10223 8902
rect 10279 8846 10350 8902
rect 10010 8760 10350 8846
rect 10010 8704 10081 8760
rect 10137 8704 10223 8760
rect 10279 8704 10350 8760
rect 10010 8618 10350 8704
rect 10010 8562 10081 8618
rect 10137 8562 10223 8618
rect 10279 8562 10350 8618
rect 10010 8476 10350 8562
rect 10010 8420 10081 8476
rect 10137 8420 10223 8476
rect 10279 8420 10350 8476
rect 10010 8334 10350 8420
rect 10010 8278 10081 8334
rect 10137 8278 10223 8334
rect 10279 8278 10350 8334
rect 10010 8192 10350 8278
rect 10010 8136 10081 8192
rect 10137 8136 10223 8192
rect 10279 8136 10350 8192
rect 10010 8050 10350 8136
rect 10010 7994 10081 8050
rect 10137 7994 10223 8050
rect 10279 7994 10350 8050
rect 10010 7908 10350 7994
rect 10010 7852 10081 7908
rect 10137 7852 10223 7908
rect 10279 7852 10350 7908
rect 10010 7766 10350 7852
rect 10010 7710 10081 7766
rect 10137 7710 10223 7766
rect 10279 7710 10350 7766
rect 10010 7624 10350 7710
rect 10010 7568 10081 7624
rect 10137 7568 10223 7624
rect 10279 7568 10350 7624
rect 10010 7482 10350 7568
rect 10010 7426 10081 7482
rect 10137 7426 10223 7482
rect 10279 7426 10350 7482
rect 10010 7340 10350 7426
rect 10010 7284 10081 7340
rect 10137 7284 10223 7340
rect 10279 7284 10350 7340
rect 10010 7198 10350 7284
rect 10010 7142 10081 7198
rect 10137 7142 10223 7198
rect 10279 7142 10350 7198
rect 10010 7056 10350 7142
rect 10010 7000 10081 7056
rect 10137 7000 10223 7056
rect 10279 7000 10350 7056
rect 10010 6914 10350 7000
rect 10010 6858 10081 6914
rect 10137 6858 10223 6914
rect 10279 6858 10350 6914
rect 10010 6772 10350 6858
rect 10010 6716 10081 6772
rect 10137 6716 10223 6772
rect 10279 6716 10350 6772
rect 10010 6630 10350 6716
rect 10010 6574 10081 6630
rect 10137 6574 10223 6630
rect 10279 6574 10350 6630
rect 10010 6488 10350 6574
rect 10010 6432 10081 6488
rect 10137 6432 10223 6488
rect 10279 6432 10350 6488
rect 10010 6346 10350 6432
rect 10010 6290 10081 6346
rect 10137 6290 10223 6346
rect 10279 6290 10350 6346
rect 10010 6204 10350 6290
rect 10010 6148 10081 6204
rect 10137 6148 10223 6204
rect 10279 6148 10350 6204
rect 10010 6062 10350 6148
rect 10010 6006 10081 6062
rect 10137 6006 10223 6062
rect 10279 6006 10350 6062
rect 10010 5920 10350 6006
rect 10010 5864 10081 5920
rect 10137 5864 10223 5920
rect 10279 5864 10350 5920
rect 10010 5778 10350 5864
rect 10010 5722 10081 5778
rect 10137 5722 10223 5778
rect 10279 5722 10350 5778
rect 10010 5636 10350 5722
rect 10010 5580 10081 5636
rect 10137 5580 10223 5636
rect 10279 5580 10350 5636
rect 10010 5494 10350 5580
rect 10010 5438 10081 5494
rect 10137 5438 10223 5494
rect 10279 5438 10350 5494
rect 10010 5352 10350 5438
rect 10010 5296 10081 5352
rect 10137 5296 10223 5352
rect 10279 5296 10350 5352
rect 10010 5210 10350 5296
rect 10010 5154 10081 5210
rect 10137 5154 10223 5210
rect 10279 5154 10350 5210
rect 10010 5068 10350 5154
rect 10010 5012 10081 5068
rect 10137 5012 10223 5068
rect 10279 5012 10350 5068
rect 10010 4926 10350 5012
rect 10010 4870 10081 4926
rect 10137 4870 10223 4926
rect 10279 4870 10350 4926
rect 10010 4784 10350 4870
rect 10010 4728 10081 4784
rect 10137 4728 10223 4784
rect 10279 4728 10350 4784
rect 10010 4642 10350 4728
rect 10010 4586 10081 4642
rect 10137 4586 10223 4642
rect 10279 4586 10350 4642
rect 10010 4500 10350 4586
rect 10010 4444 10081 4500
rect 10137 4444 10223 4500
rect 10279 4444 10350 4500
rect 10010 4358 10350 4444
rect 10010 4302 10081 4358
rect 10137 4302 10223 4358
rect 10279 4302 10350 4358
rect 10010 4216 10350 4302
rect 10010 4160 10081 4216
rect 10137 4160 10223 4216
rect 10279 4160 10350 4216
rect 10010 4074 10350 4160
rect 10010 4018 10081 4074
rect 10137 4018 10223 4074
rect 10279 4018 10350 4074
rect 10010 3932 10350 4018
rect 10010 3876 10081 3932
rect 10137 3876 10223 3932
rect 10279 3876 10350 3932
rect 10010 3790 10350 3876
rect 10010 3734 10081 3790
rect 10137 3734 10223 3790
rect 10279 3734 10350 3790
rect 10010 3648 10350 3734
rect 10010 3592 10081 3648
rect 10137 3592 10223 3648
rect 10279 3592 10350 3648
rect 10010 3506 10350 3592
rect 10010 3450 10081 3506
rect 10137 3450 10223 3506
rect 10279 3450 10350 3506
rect 10010 3364 10350 3450
rect 10010 3308 10081 3364
rect 10137 3308 10223 3364
rect 10279 3308 10350 3364
rect 10010 3222 10350 3308
rect 10010 3166 10081 3222
rect 10137 3166 10223 3222
rect 10279 3166 10350 3222
rect 10010 3080 10350 3166
rect 10010 3024 10081 3080
rect 10137 3024 10223 3080
rect 10279 3024 10350 3080
rect 10010 2938 10350 3024
rect 10010 2882 10081 2938
rect 10137 2882 10223 2938
rect 10279 2882 10350 2938
rect 10010 2796 10350 2882
rect 10010 2740 10081 2796
rect 10137 2740 10223 2796
rect 10279 2740 10350 2796
rect 10010 2654 10350 2740
rect 10010 2598 10081 2654
rect 10137 2598 10223 2654
rect 10279 2598 10350 2654
rect 10010 2512 10350 2598
rect 10010 2456 10081 2512
rect 10137 2456 10223 2512
rect 10279 2456 10350 2512
rect 10010 2370 10350 2456
rect 10010 2314 10081 2370
rect 10137 2314 10223 2370
rect 10279 2314 10350 2370
rect 10010 2228 10350 2314
rect 10010 2172 10081 2228
rect 10137 2172 10223 2228
rect 10279 2172 10350 2228
rect 10010 2086 10350 2172
rect 10010 2030 10081 2086
rect 10137 2030 10223 2086
rect 10279 2030 10350 2086
rect 10010 1944 10350 2030
rect 10010 1888 10081 1944
rect 10137 1888 10223 1944
rect 10279 1888 10350 1944
rect 10010 1802 10350 1888
rect 10010 1746 10081 1802
rect 10137 1746 10223 1802
rect 10279 1746 10350 1802
rect 10010 1660 10350 1746
rect 10010 1604 10081 1660
rect 10137 1604 10223 1660
rect 10279 1604 10350 1660
rect 10010 1518 10350 1604
rect 10010 1462 10081 1518
rect 10137 1462 10223 1518
rect 10279 1462 10350 1518
rect 10010 1376 10350 1462
rect 10010 1320 10081 1376
rect 10137 1320 10223 1376
rect 10279 1320 10350 1376
rect 10010 1234 10350 1320
rect 10010 1178 10081 1234
rect 10137 1178 10223 1234
rect 10279 1178 10350 1234
rect 10010 1092 10350 1178
rect 10010 1036 10081 1092
rect 10137 1036 10223 1092
rect 10279 1036 10350 1092
rect 10010 950 10350 1036
rect 10010 894 10081 950
rect 10137 894 10223 950
rect 10279 894 10350 950
rect 10010 808 10350 894
rect 10010 752 10081 808
rect 10137 752 10223 808
rect 10279 752 10350 808
rect 10010 666 10350 752
rect 10010 610 10081 666
rect 10137 610 10223 666
rect 10279 610 10350 666
rect 10010 524 10350 610
rect 10010 468 10081 524
rect 10137 468 10223 524
rect 10279 468 10350 524
rect 10010 458 10350 468
rect 10550 12310 10890 12320
rect 10550 12254 10622 12310
rect 10678 12254 10764 12310
rect 10820 12254 10890 12310
rect 10550 12168 10890 12254
rect 10550 12112 10622 12168
rect 10678 12112 10764 12168
rect 10820 12112 10890 12168
rect 10550 12026 10890 12112
rect 10550 11970 10622 12026
rect 10678 11970 10764 12026
rect 10820 11970 10890 12026
rect 10550 11884 10890 11970
rect 10550 11828 10622 11884
rect 10678 11828 10764 11884
rect 10820 11828 10890 11884
rect 10550 11742 10890 11828
rect 10550 11686 10622 11742
rect 10678 11686 10764 11742
rect 10820 11686 10890 11742
rect 10550 11600 10890 11686
rect 10550 11544 10622 11600
rect 10678 11544 10764 11600
rect 10820 11544 10890 11600
rect 10550 11458 10890 11544
rect 10550 11402 10622 11458
rect 10678 11402 10764 11458
rect 10820 11402 10890 11458
rect 10550 11316 10890 11402
rect 10550 11260 10622 11316
rect 10678 11260 10764 11316
rect 10820 11260 10890 11316
rect 10550 11174 10890 11260
rect 10550 11118 10622 11174
rect 10678 11118 10764 11174
rect 10820 11118 10890 11174
rect 10550 11032 10890 11118
rect 10550 10976 10622 11032
rect 10678 10976 10764 11032
rect 10820 10976 10890 11032
rect 10550 10890 10890 10976
rect 10550 10834 10622 10890
rect 10678 10834 10764 10890
rect 10820 10834 10890 10890
rect 10550 10748 10890 10834
rect 10550 10692 10622 10748
rect 10678 10692 10764 10748
rect 10820 10692 10890 10748
rect 10550 10606 10890 10692
rect 10550 10550 10622 10606
rect 10678 10550 10764 10606
rect 10820 10550 10890 10606
rect 10550 10464 10890 10550
rect 10550 10408 10622 10464
rect 10678 10408 10764 10464
rect 10820 10408 10890 10464
rect 10550 10322 10890 10408
rect 10550 10266 10622 10322
rect 10678 10266 10764 10322
rect 10820 10266 10890 10322
rect 10550 10180 10890 10266
rect 10550 10124 10622 10180
rect 10678 10124 10764 10180
rect 10820 10124 10890 10180
rect 10550 10038 10890 10124
rect 10550 9982 10622 10038
rect 10678 9982 10764 10038
rect 10820 9982 10890 10038
rect 10550 9896 10890 9982
rect 10550 9840 10622 9896
rect 10678 9840 10764 9896
rect 10820 9840 10890 9896
rect 10550 9754 10890 9840
rect 10550 9698 10622 9754
rect 10678 9698 10764 9754
rect 10820 9698 10890 9754
rect 10550 9612 10890 9698
rect 10550 9556 10622 9612
rect 10678 9556 10764 9612
rect 10820 9556 10890 9612
rect 10550 9470 10890 9556
rect 10550 9414 10622 9470
rect 10678 9414 10764 9470
rect 10820 9414 10890 9470
rect 10550 9328 10890 9414
rect 10550 9272 10622 9328
rect 10678 9272 10764 9328
rect 10820 9272 10890 9328
rect 10550 9186 10890 9272
rect 10550 9130 10622 9186
rect 10678 9130 10764 9186
rect 10820 9130 10890 9186
rect 10550 9044 10890 9130
rect 10550 8988 10622 9044
rect 10678 8988 10764 9044
rect 10820 8988 10890 9044
rect 10550 8902 10890 8988
rect 10550 8846 10622 8902
rect 10678 8846 10764 8902
rect 10820 8846 10890 8902
rect 10550 8760 10890 8846
rect 10550 8704 10622 8760
rect 10678 8704 10764 8760
rect 10820 8704 10890 8760
rect 10550 8618 10890 8704
rect 10550 8562 10622 8618
rect 10678 8562 10764 8618
rect 10820 8562 10890 8618
rect 10550 8476 10890 8562
rect 10550 8420 10622 8476
rect 10678 8420 10764 8476
rect 10820 8420 10890 8476
rect 10550 8334 10890 8420
rect 10550 8278 10622 8334
rect 10678 8278 10764 8334
rect 10820 8278 10890 8334
rect 10550 8192 10890 8278
rect 10550 8136 10622 8192
rect 10678 8136 10764 8192
rect 10820 8136 10890 8192
rect 10550 8050 10890 8136
rect 10550 7994 10622 8050
rect 10678 7994 10764 8050
rect 10820 7994 10890 8050
rect 10550 7908 10890 7994
rect 10550 7852 10622 7908
rect 10678 7852 10764 7908
rect 10820 7852 10890 7908
rect 10550 7766 10890 7852
rect 10550 7710 10622 7766
rect 10678 7710 10764 7766
rect 10820 7710 10890 7766
rect 10550 7624 10890 7710
rect 10550 7568 10622 7624
rect 10678 7568 10764 7624
rect 10820 7568 10890 7624
rect 10550 7482 10890 7568
rect 10550 7426 10622 7482
rect 10678 7426 10764 7482
rect 10820 7426 10890 7482
rect 10550 7340 10890 7426
rect 10550 7284 10622 7340
rect 10678 7284 10764 7340
rect 10820 7284 10890 7340
rect 10550 7198 10890 7284
rect 10550 7142 10622 7198
rect 10678 7142 10764 7198
rect 10820 7142 10890 7198
rect 10550 7056 10890 7142
rect 10550 7000 10622 7056
rect 10678 7000 10764 7056
rect 10820 7000 10890 7056
rect 10550 6914 10890 7000
rect 10550 6858 10622 6914
rect 10678 6858 10764 6914
rect 10820 6858 10890 6914
rect 10550 6772 10890 6858
rect 10550 6716 10622 6772
rect 10678 6716 10764 6772
rect 10820 6716 10890 6772
rect 10550 6630 10890 6716
rect 10550 6574 10622 6630
rect 10678 6574 10764 6630
rect 10820 6574 10890 6630
rect 10550 6488 10890 6574
rect 10550 6432 10622 6488
rect 10678 6432 10764 6488
rect 10820 6432 10890 6488
rect 10550 6346 10890 6432
rect 10550 6290 10622 6346
rect 10678 6290 10764 6346
rect 10820 6290 10890 6346
rect 10550 6204 10890 6290
rect 10550 6148 10622 6204
rect 10678 6148 10764 6204
rect 10820 6148 10890 6204
rect 10550 6062 10890 6148
rect 10550 6006 10622 6062
rect 10678 6006 10764 6062
rect 10820 6006 10890 6062
rect 10550 5920 10890 6006
rect 10550 5864 10622 5920
rect 10678 5864 10764 5920
rect 10820 5864 10890 5920
rect 10550 5778 10890 5864
rect 10550 5722 10622 5778
rect 10678 5722 10764 5778
rect 10820 5722 10890 5778
rect 10550 5636 10890 5722
rect 10550 5580 10622 5636
rect 10678 5580 10764 5636
rect 10820 5580 10890 5636
rect 10550 5494 10890 5580
rect 10550 5438 10622 5494
rect 10678 5438 10764 5494
rect 10820 5438 10890 5494
rect 10550 5352 10890 5438
rect 10550 5296 10622 5352
rect 10678 5296 10764 5352
rect 10820 5296 10890 5352
rect 10550 5210 10890 5296
rect 10550 5154 10622 5210
rect 10678 5154 10764 5210
rect 10820 5154 10890 5210
rect 10550 5068 10890 5154
rect 10550 5012 10622 5068
rect 10678 5012 10764 5068
rect 10820 5012 10890 5068
rect 10550 4926 10890 5012
rect 10550 4870 10622 4926
rect 10678 4870 10764 4926
rect 10820 4870 10890 4926
rect 10550 4784 10890 4870
rect 10550 4728 10622 4784
rect 10678 4728 10764 4784
rect 10820 4728 10890 4784
rect 10550 4642 10890 4728
rect 10550 4586 10622 4642
rect 10678 4586 10764 4642
rect 10820 4586 10890 4642
rect 10550 4500 10890 4586
rect 10550 4444 10622 4500
rect 10678 4444 10764 4500
rect 10820 4444 10890 4500
rect 10550 4358 10890 4444
rect 10550 4302 10622 4358
rect 10678 4302 10764 4358
rect 10820 4302 10890 4358
rect 10550 4216 10890 4302
rect 10550 4160 10622 4216
rect 10678 4160 10764 4216
rect 10820 4160 10890 4216
rect 10550 4074 10890 4160
rect 10550 4018 10622 4074
rect 10678 4018 10764 4074
rect 10820 4018 10890 4074
rect 10550 3932 10890 4018
rect 10550 3876 10622 3932
rect 10678 3876 10764 3932
rect 10820 3876 10890 3932
rect 10550 3790 10890 3876
rect 10550 3734 10622 3790
rect 10678 3734 10764 3790
rect 10820 3734 10890 3790
rect 10550 3648 10890 3734
rect 10550 3592 10622 3648
rect 10678 3592 10764 3648
rect 10820 3592 10890 3648
rect 10550 3506 10890 3592
rect 10550 3450 10622 3506
rect 10678 3450 10764 3506
rect 10820 3450 10890 3506
rect 10550 3364 10890 3450
rect 10550 3308 10622 3364
rect 10678 3308 10764 3364
rect 10820 3308 10890 3364
rect 10550 3222 10890 3308
rect 10550 3166 10622 3222
rect 10678 3166 10764 3222
rect 10820 3166 10890 3222
rect 10550 3080 10890 3166
rect 10550 3024 10622 3080
rect 10678 3024 10764 3080
rect 10820 3024 10890 3080
rect 10550 2938 10890 3024
rect 10550 2882 10622 2938
rect 10678 2882 10764 2938
rect 10820 2882 10890 2938
rect 10550 2796 10890 2882
rect 10550 2740 10622 2796
rect 10678 2740 10764 2796
rect 10820 2740 10890 2796
rect 10550 2654 10890 2740
rect 10550 2598 10622 2654
rect 10678 2598 10764 2654
rect 10820 2598 10890 2654
rect 10550 2512 10890 2598
rect 10550 2456 10622 2512
rect 10678 2456 10764 2512
rect 10820 2456 10890 2512
rect 10550 2370 10890 2456
rect 10550 2314 10622 2370
rect 10678 2314 10764 2370
rect 10820 2314 10890 2370
rect 10550 2228 10890 2314
rect 10550 2172 10622 2228
rect 10678 2172 10764 2228
rect 10820 2172 10890 2228
rect 10550 2086 10890 2172
rect 10550 2030 10622 2086
rect 10678 2030 10764 2086
rect 10820 2030 10890 2086
rect 10550 1944 10890 2030
rect 10550 1888 10622 1944
rect 10678 1888 10764 1944
rect 10820 1888 10890 1944
rect 10550 1802 10890 1888
rect 10550 1746 10622 1802
rect 10678 1746 10764 1802
rect 10820 1746 10890 1802
rect 10550 1660 10890 1746
rect 10550 1604 10622 1660
rect 10678 1604 10764 1660
rect 10820 1604 10890 1660
rect 10550 1518 10890 1604
rect 10550 1462 10622 1518
rect 10678 1462 10764 1518
rect 10820 1462 10890 1518
rect 10550 1376 10890 1462
rect 10550 1320 10622 1376
rect 10678 1320 10764 1376
rect 10820 1320 10890 1376
rect 10550 1234 10890 1320
rect 10550 1178 10622 1234
rect 10678 1178 10764 1234
rect 10820 1178 10890 1234
rect 10550 1092 10890 1178
rect 10550 1036 10622 1092
rect 10678 1036 10764 1092
rect 10820 1036 10890 1092
rect 10550 950 10890 1036
rect 10550 894 10622 950
rect 10678 894 10764 950
rect 10820 894 10890 950
rect 10550 808 10890 894
rect 10550 752 10622 808
rect 10678 752 10764 808
rect 10820 752 10890 808
rect 10550 666 10890 752
rect 10550 610 10622 666
rect 10678 610 10764 666
rect 10820 610 10890 666
rect 10550 524 10890 610
rect 10550 468 10622 524
rect 10678 468 10764 524
rect 10820 468 10890 524
rect 10550 458 10890 468
rect 11090 12310 11430 12320
rect 11090 12254 11162 12310
rect 11218 12254 11304 12310
rect 11360 12254 11430 12310
rect 11090 12168 11430 12254
rect 11090 12112 11162 12168
rect 11218 12112 11304 12168
rect 11360 12112 11430 12168
rect 11090 12026 11430 12112
rect 11090 11970 11162 12026
rect 11218 11970 11304 12026
rect 11360 11970 11430 12026
rect 11090 11884 11430 11970
rect 11090 11828 11162 11884
rect 11218 11828 11304 11884
rect 11360 11828 11430 11884
rect 11090 11742 11430 11828
rect 11090 11686 11162 11742
rect 11218 11686 11304 11742
rect 11360 11686 11430 11742
rect 11090 11600 11430 11686
rect 11090 11544 11162 11600
rect 11218 11544 11304 11600
rect 11360 11544 11430 11600
rect 11090 11458 11430 11544
rect 11090 11402 11162 11458
rect 11218 11402 11304 11458
rect 11360 11402 11430 11458
rect 11090 11316 11430 11402
rect 11090 11260 11162 11316
rect 11218 11260 11304 11316
rect 11360 11260 11430 11316
rect 11090 11174 11430 11260
rect 11090 11118 11162 11174
rect 11218 11118 11304 11174
rect 11360 11118 11430 11174
rect 11090 11032 11430 11118
rect 11090 10976 11162 11032
rect 11218 10976 11304 11032
rect 11360 10976 11430 11032
rect 11090 10890 11430 10976
rect 11090 10834 11162 10890
rect 11218 10834 11304 10890
rect 11360 10834 11430 10890
rect 11090 10748 11430 10834
rect 11090 10692 11162 10748
rect 11218 10692 11304 10748
rect 11360 10692 11430 10748
rect 11090 10606 11430 10692
rect 11090 10550 11162 10606
rect 11218 10550 11304 10606
rect 11360 10550 11430 10606
rect 11090 10464 11430 10550
rect 11090 10408 11162 10464
rect 11218 10408 11304 10464
rect 11360 10408 11430 10464
rect 11090 10322 11430 10408
rect 11090 10266 11162 10322
rect 11218 10266 11304 10322
rect 11360 10266 11430 10322
rect 11090 10180 11430 10266
rect 11090 10124 11162 10180
rect 11218 10124 11304 10180
rect 11360 10124 11430 10180
rect 11090 10038 11430 10124
rect 11090 9982 11162 10038
rect 11218 9982 11304 10038
rect 11360 9982 11430 10038
rect 11090 9896 11430 9982
rect 11090 9840 11162 9896
rect 11218 9840 11304 9896
rect 11360 9840 11430 9896
rect 11090 9754 11430 9840
rect 11090 9698 11162 9754
rect 11218 9698 11304 9754
rect 11360 9698 11430 9754
rect 11090 9612 11430 9698
rect 11090 9556 11162 9612
rect 11218 9556 11304 9612
rect 11360 9556 11430 9612
rect 11090 9470 11430 9556
rect 11090 9414 11162 9470
rect 11218 9414 11304 9470
rect 11360 9414 11430 9470
rect 11090 9328 11430 9414
rect 11090 9272 11162 9328
rect 11218 9272 11304 9328
rect 11360 9272 11430 9328
rect 11090 9186 11430 9272
rect 11090 9130 11162 9186
rect 11218 9130 11304 9186
rect 11360 9130 11430 9186
rect 11090 9044 11430 9130
rect 11090 8988 11162 9044
rect 11218 8988 11304 9044
rect 11360 8988 11430 9044
rect 11090 8902 11430 8988
rect 11090 8846 11162 8902
rect 11218 8846 11304 8902
rect 11360 8846 11430 8902
rect 11090 8760 11430 8846
rect 11090 8704 11162 8760
rect 11218 8704 11304 8760
rect 11360 8704 11430 8760
rect 11090 8618 11430 8704
rect 11090 8562 11162 8618
rect 11218 8562 11304 8618
rect 11360 8562 11430 8618
rect 11090 8476 11430 8562
rect 11090 8420 11162 8476
rect 11218 8420 11304 8476
rect 11360 8420 11430 8476
rect 11090 8334 11430 8420
rect 11090 8278 11162 8334
rect 11218 8278 11304 8334
rect 11360 8278 11430 8334
rect 11090 8192 11430 8278
rect 11090 8136 11162 8192
rect 11218 8136 11304 8192
rect 11360 8136 11430 8192
rect 11090 8050 11430 8136
rect 11090 7994 11162 8050
rect 11218 7994 11304 8050
rect 11360 7994 11430 8050
rect 11090 7908 11430 7994
rect 11090 7852 11162 7908
rect 11218 7852 11304 7908
rect 11360 7852 11430 7908
rect 11090 7766 11430 7852
rect 11090 7710 11162 7766
rect 11218 7710 11304 7766
rect 11360 7710 11430 7766
rect 11090 7624 11430 7710
rect 11090 7568 11162 7624
rect 11218 7568 11304 7624
rect 11360 7568 11430 7624
rect 11090 7482 11430 7568
rect 11090 7426 11162 7482
rect 11218 7426 11304 7482
rect 11360 7426 11430 7482
rect 11090 7340 11430 7426
rect 11090 7284 11162 7340
rect 11218 7284 11304 7340
rect 11360 7284 11430 7340
rect 11090 7198 11430 7284
rect 11090 7142 11162 7198
rect 11218 7142 11304 7198
rect 11360 7142 11430 7198
rect 11090 7056 11430 7142
rect 11090 7000 11162 7056
rect 11218 7000 11304 7056
rect 11360 7000 11430 7056
rect 11090 6914 11430 7000
rect 11090 6858 11162 6914
rect 11218 6858 11304 6914
rect 11360 6858 11430 6914
rect 11090 6772 11430 6858
rect 11090 6716 11162 6772
rect 11218 6716 11304 6772
rect 11360 6716 11430 6772
rect 11090 6630 11430 6716
rect 11090 6574 11162 6630
rect 11218 6574 11304 6630
rect 11360 6574 11430 6630
rect 11090 6488 11430 6574
rect 11090 6432 11162 6488
rect 11218 6432 11304 6488
rect 11360 6432 11430 6488
rect 11090 6346 11430 6432
rect 11090 6290 11162 6346
rect 11218 6290 11304 6346
rect 11360 6290 11430 6346
rect 11090 6204 11430 6290
rect 11090 6148 11162 6204
rect 11218 6148 11304 6204
rect 11360 6148 11430 6204
rect 11090 6062 11430 6148
rect 11090 6006 11162 6062
rect 11218 6006 11304 6062
rect 11360 6006 11430 6062
rect 11090 5920 11430 6006
rect 11090 5864 11162 5920
rect 11218 5864 11304 5920
rect 11360 5864 11430 5920
rect 11090 5778 11430 5864
rect 11090 5722 11162 5778
rect 11218 5722 11304 5778
rect 11360 5722 11430 5778
rect 11090 5636 11430 5722
rect 11090 5580 11162 5636
rect 11218 5580 11304 5636
rect 11360 5580 11430 5636
rect 11090 5494 11430 5580
rect 11090 5438 11162 5494
rect 11218 5438 11304 5494
rect 11360 5438 11430 5494
rect 11090 5352 11430 5438
rect 11090 5296 11162 5352
rect 11218 5296 11304 5352
rect 11360 5296 11430 5352
rect 11090 5210 11430 5296
rect 11090 5154 11162 5210
rect 11218 5154 11304 5210
rect 11360 5154 11430 5210
rect 11090 5068 11430 5154
rect 11090 5012 11162 5068
rect 11218 5012 11304 5068
rect 11360 5012 11430 5068
rect 11090 4926 11430 5012
rect 11090 4870 11162 4926
rect 11218 4870 11304 4926
rect 11360 4870 11430 4926
rect 11090 4784 11430 4870
rect 11090 4728 11162 4784
rect 11218 4728 11304 4784
rect 11360 4728 11430 4784
rect 11090 4642 11430 4728
rect 11090 4586 11162 4642
rect 11218 4586 11304 4642
rect 11360 4586 11430 4642
rect 11090 4500 11430 4586
rect 11090 4444 11162 4500
rect 11218 4444 11304 4500
rect 11360 4444 11430 4500
rect 11090 4358 11430 4444
rect 11090 4302 11162 4358
rect 11218 4302 11304 4358
rect 11360 4302 11430 4358
rect 11090 4216 11430 4302
rect 11090 4160 11162 4216
rect 11218 4160 11304 4216
rect 11360 4160 11430 4216
rect 11090 4074 11430 4160
rect 11090 4018 11162 4074
rect 11218 4018 11304 4074
rect 11360 4018 11430 4074
rect 11090 3932 11430 4018
rect 11090 3876 11162 3932
rect 11218 3876 11304 3932
rect 11360 3876 11430 3932
rect 11090 3790 11430 3876
rect 11090 3734 11162 3790
rect 11218 3734 11304 3790
rect 11360 3734 11430 3790
rect 11090 3648 11430 3734
rect 11090 3592 11162 3648
rect 11218 3592 11304 3648
rect 11360 3592 11430 3648
rect 11090 3506 11430 3592
rect 11090 3450 11162 3506
rect 11218 3450 11304 3506
rect 11360 3450 11430 3506
rect 11090 3364 11430 3450
rect 11090 3308 11162 3364
rect 11218 3308 11304 3364
rect 11360 3308 11430 3364
rect 11090 3222 11430 3308
rect 11090 3166 11162 3222
rect 11218 3166 11304 3222
rect 11360 3166 11430 3222
rect 11090 3080 11430 3166
rect 11090 3024 11162 3080
rect 11218 3024 11304 3080
rect 11360 3024 11430 3080
rect 11090 2938 11430 3024
rect 11090 2882 11162 2938
rect 11218 2882 11304 2938
rect 11360 2882 11430 2938
rect 11090 2796 11430 2882
rect 11090 2740 11162 2796
rect 11218 2740 11304 2796
rect 11360 2740 11430 2796
rect 11090 2654 11430 2740
rect 11090 2598 11162 2654
rect 11218 2598 11304 2654
rect 11360 2598 11430 2654
rect 11090 2512 11430 2598
rect 11090 2456 11162 2512
rect 11218 2456 11304 2512
rect 11360 2456 11430 2512
rect 11090 2370 11430 2456
rect 11090 2314 11162 2370
rect 11218 2314 11304 2370
rect 11360 2314 11430 2370
rect 11090 2228 11430 2314
rect 11090 2172 11162 2228
rect 11218 2172 11304 2228
rect 11360 2172 11430 2228
rect 11090 2086 11430 2172
rect 11090 2030 11162 2086
rect 11218 2030 11304 2086
rect 11360 2030 11430 2086
rect 11090 1944 11430 2030
rect 11090 1888 11162 1944
rect 11218 1888 11304 1944
rect 11360 1888 11430 1944
rect 11090 1802 11430 1888
rect 11090 1746 11162 1802
rect 11218 1746 11304 1802
rect 11360 1746 11430 1802
rect 11090 1660 11430 1746
rect 11090 1604 11162 1660
rect 11218 1604 11304 1660
rect 11360 1604 11430 1660
rect 11090 1518 11430 1604
rect 11090 1462 11162 1518
rect 11218 1462 11304 1518
rect 11360 1462 11430 1518
rect 11090 1376 11430 1462
rect 11090 1320 11162 1376
rect 11218 1320 11304 1376
rect 11360 1320 11430 1376
rect 11090 1234 11430 1320
rect 11090 1178 11162 1234
rect 11218 1178 11304 1234
rect 11360 1178 11430 1234
rect 11090 1092 11430 1178
rect 11090 1036 11162 1092
rect 11218 1036 11304 1092
rect 11360 1036 11430 1092
rect 11090 950 11430 1036
rect 11090 894 11162 950
rect 11218 894 11304 950
rect 11360 894 11430 950
rect 11090 808 11430 894
rect 11090 752 11162 808
rect 11218 752 11304 808
rect 11360 752 11430 808
rect 11090 666 11430 752
rect 11090 610 11162 666
rect 11218 610 11304 666
rect 11360 610 11430 666
rect 11090 524 11430 610
rect 11090 468 11162 524
rect 11218 468 11304 524
rect 11360 468 11430 524
rect 11090 458 11430 468
rect 11630 12310 11970 12320
rect 11630 12254 11702 12310
rect 11758 12254 11844 12310
rect 11900 12254 11970 12310
rect 11630 12168 11970 12254
rect 11630 12112 11702 12168
rect 11758 12112 11844 12168
rect 11900 12112 11970 12168
rect 11630 12026 11970 12112
rect 11630 11970 11702 12026
rect 11758 11970 11844 12026
rect 11900 11970 11970 12026
rect 11630 11884 11970 11970
rect 11630 11828 11702 11884
rect 11758 11828 11844 11884
rect 11900 11828 11970 11884
rect 11630 11742 11970 11828
rect 11630 11686 11702 11742
rect 11758 11686 11844 11742
rect 11900 11686 11970 11742
rect 11630 11600 11970 11686
rect 11630 11544 11702 11600
rect 11758 11544 11844 11600
rect 11900 11544 11970 11600
rect 11630 11458 11970 11544
rect 11630 11402 11702 11458
rect 11758 11402 11844 11458
rect 11900 11402 11970 11458
rect 11630 11316 11970 11402
rect 11630 11260 11702 11316
rect 11758 11260 11844 11316
rect 11900 11260 11970 11316
rect 11630 11174 11970 11260
rect 11630 11118 11702 11174
rect 11758 11118 11844 11174
rect 11900 11118 11970 11174
rect 11630 11032 11970 11118
rect 11630 10976 11702 11032
rect 11758 10976 11844 11032
rect 11900 10976 11970 11032
rect 11630 10890 11970 10976
rect 11630 10834 11702 10890
rect 11758 10834 11844 10890
rect 11900 10834 11970 10890
rect 11630 10748 11970 10834
rect 11630 10692 11702 10748
rect 11758 10692 11844 10748
rect 11900 10692 11970 10748
rect 11630 10606 11970 10692
rect 11630 10550 11702 10606
rect 11758 10550 11844 10606
rect 11900 10550 11970 10606
rect 11630 10464 11970 10550
rect 11630 10408 11702 10464
rect 11758 10408 11844 10464
rect 11900 10408 11970 10464
rect 11630 10322 11970 10408
rect 11630 10266 11702 10322
rect 11758 10266 11844 10322
rect 11900 10266 11970 10322
rect 11630 10180 11970 10266
rect 11630 10124 11702 10180
rect 11758 10124 11844 10180
rect 11900 10124 11970 10180
rect 11630 10038 11970 10124
rect 11630 9982 11702 10038
rect 11758 9982 11844 10038
rect 11900 9982 11970 10038
rect 11630 9896 11970 9982
rect 11630 9840 11702 9896
rect 11758 9840 11844 9896
rect 11900 9840 11970 9896
rect 11630 9754 11970 9840
rect 11630 9698 11702 9754
rect 11758 9698 11844 9754
rect 11900 9698 11970 9754
rect 11630 9612 11970 9698
rect 11630 9556 11702 9612
rect 11758 9556 11844 9612
rect 11900 9556 11970 9612
rect 11630 9470 11970 9556
rect 11630 9414 11702 9470
rect 11758 9414 11844 9470
rect 11900 9414 11970 9470
rect 11630 9328 11970 9414
rect 11630 9272 11702 9328
rect 11758 9272 11844 9328
rect 11900 9272 11970 9328
rect 11630 9186 11970 9272
rect 11630 9130 11702 9186
rect 11758 9130 11844 9186
rect 11900 9130 11970 9186
rect 11630 9044 11970 9130
rect 11630 8988 11702 9044
rect 11758 8988 11844 9044
rect 11900 8988 11970 9044
rect 11630 8902 11970 8988
rect 11630 8846 11702 8902
rect 11758 8846 11844 8902
rect 11900 8846 11970 8902
rect 11630 8760 11970 8846
rect 11630 8704 11702 8760
rect 11758 8704 11844 8760
rect 11900 8704 11970 8760
rect 11630 8618 11970 8704
rect 11630 8562 11702 8618
rect 11758 8562 11844 8618
rect 11900 8562 11970 8618
rect 11630 8476 11970 8562
rect 11630 8420 11702 8476
rect 11758 8420 11844 8476
rect 11900 8420 11970 8476
rect 11630 8334 11970 8420
rect 11630 8278 11702 8334
rect 11758 8278 11844 8334
rect 11900 8278 11970 8334
rect 11630 8192 11970 8278
rect 11630 8136 11702 8192
rect 11758 8136 11844 8192
rect 11900 8136 11970 8192
rect 11630 8050 11970 8136
rect 11630 7994 11702 8050
rect 11758 7994 11844 8050
rect 11900 7994 11970 8050
rect 11630 7908 11970 7994
rect 11630 7852 11702 7908
rect 11758 7852 11844 7908
rect 11900 7852 11970 7908
rect 11630 7766 11970 7852
rect 11630 7710 11702 7766
rect 11758 7710 11844 7766
rect 11900 7710 11970 7766
rect 11630 7624 11970 7710
rect 11630 7568 11702 7624
rect 11758 7568 11844 7624
rect 11900 7568 11970 7624
rect 11630 7482 11970 7568
rect 11630 7426 11702 7482
rect 11758 7426 11844 7482
rect 11900 7426 11970 7482
rect 11630 7340 11970 7426
rect 11630 7284 11702 7340
rect 11758 7284 11844 7340
rect 11900 7284 11970 7340
rect 11630 7198 11970 7284
rect 11630 7142 11702 7198
rect 11758 7142 11844 7198
rect 11900 7142 11970 7198
rect 11630 7056 11970 7142
rect 11630 7000 11702 7056
rect 11758 7000 11844 7056
rect 11900 7000 11970 7056
rect 11630 6914 11970 7000
rect 11630 6858 11702 6914
rect 11758 6858 11844 6914
rect 11900 6858 11970 6914
rect 11630 6772 11970 6858
rect 11630 6716 11702 6772
rect 11758 6716 11844 6772
rect 11900 6716 11970 6772
rect 11630 6630 11970 6716
rect 11630 6574 11702 6630
rect 11758 6574 11844 6630
rect 11900 6574 11970 6630
rect 11630 6488 11970 6574
rect 11630 6432 11702 6488
rect 11758 6432 11844 6488
rect 11900 6432 11970 6488
rect 11630 6346 11970 6432
rect 11630 6290 11702 6346
rect 11758 6290 11844 6346
rect 11900 6290 11970 6346
rect 11630 6204 11970 6290
rect 11630 6148 11702 6204
rect 11758 6148 11844 6204
rect 11900 6148 11970 6204
rect 11630 6062 11970 6148
rect 11630 6006 11702 6062
rect 11758 6006 11844 6062
rect 11900 6006 11970 6062
rect 11630 5920 11970 6006
rect 11630 5864 11702 5920
rect 11758 5864 11844 5920
rect 11900 5864 11970 5920
rect 11630 5778 11970 5864
rect 11630 5722 11702 5778
rect 11758 5722 11844 5778
rect 11900 5722 11970 5778
rect 11630 5636 11970 5722
rect 11630 5580 11702 5636
rect 11758 5580 11844 5636
rect 11900 5580 11970 5636
rect 11630 5494 11970 5580
rect 11630 5438 11702 5494
rect 11758 5438 11844 5494
rect 11900 5438 11970 5494
rect 11630 5352 11970 5438
rect 11630 5296 11702 5352
rect 11758 5296 11844 5352
rect 11900 5296 11970 5352
rect 11630 5210 11970 5296
rect 11630 5154 11702 5210
rect 11758 5154 11844 5210
rect 11900 5154 11970 5210
rect 11630 5068 11970 5154
rect 11630 5012 11702 5068
rect 11758 5012 11844 5068
rect 11900 5012 11970 5068
rect 11630 4926 11970 5012
rect 11630 4870 11702 4926
rect 11758 4870 11844 4926
rect 11900 4870 11970 4926
rect 11630 4784 11970 4870
rect 11630 4728 11702 4784
rect 11758 4728 11844 4784
rect 11900 4728 11970 4784
rect 11630 4642 11970 4728
rect 11630 4586 11702 4642
rect 11758 4586 11844 4642
rect 11900 4586 11970 4642
rect 11630 4500 11970 4586
rect 11630 4444 11702 4500
rect 11758 4444 11844 4500
rect 11900 4444 11970 4500
rect 11630 4358 11970 4444
rect 11630 4302 11702 4358
rect 11758 4302 11844 4358
rect 11900 4302 11970 4358
rect 11630 4216 11970 4302
rect 11630 4160 11702 4216
rect 11758 4160 11844 4216
rect 11900 4160 11970 4216
rect 11630 4074 11970 4160
rect 11630 4018 11702 4074
rect 11758 4018 11844 4074
rect 11900 4018 11970 4074
rect 11630 3932 11970 4018
rect 11630 3876 11702 3932
rect 11758 3876 11844 3932
rect 11900 3876 11970 3932
rect 11630 3790 11970 3876
rect 11630 3734 11702 3790
rect 11758 3734 11844 3790
rect 11900 3734 11970 3790
rect 11630 3648 11970 3734
rect 11630 3592 11702 3648
rect 11758 3592 11844 3648
rect 11900 3592 11970 3648
rect 11630 3506 11970 3592
rect 11630 3450 11702 3506
rect 11758 3450 11844 3506
rect 11900 3450 11970 3506
rect 11630 3364 11970 3450
rect 11630 3308 11702 3364
rect 11758 3308 11844 3364
rect 11900 3308 11970 3364
rect 11630 3222 11970 3308
rect 11630 3166 11702 3222
rect 11758 3166 11844 3222
rect 11900 3166 11970 3222
rect 11630 3080 11970 3166
rect 11630 3024 11702 3080
rect 11758 3024 11844 3080
rect 11900 3024 11970 3080
rect 11630 2938 11970 3024
rect 11630 2882 11702 2938
rect 11758 2882 11844 2938
rect 11900 2882 11970 2938
rect 11630 2796 11970 2882
rect 11630 2740 11702 2796
rect 11758 2740 11844 2796
rect 11900 2740 11970 2796
rect 11630 2654 11970 2740
rect 11630 2598 11702 2654
rect 11758 2598 11844 2654
rect 11900 2598 11970 2654
rect 11630 2512 11970 2598
rect 11630 2456 11702 2512
rect 11758 2456 11844 2512
rect 11900 2456 11970 2512
rect 11630 2370 11970 2456
rect 11630 2314 11702 2370
rect 11758 2314 11844 2370
rect 11900 2314 11970 2370
rect 11630 2228 11970 2314
rect 11630 2172 11702 2228
rect 11758 2172 11844 2228
rect 11900 2172 11970 2228
rect 11630 2086 11970 2172
rect 11630 2030 11702 2086
rect 11758 2030 11844 2086
rect 11900 2030 11970 2086
rect 11630 1944 11970 2030
rect 11630 1888 11702 1944
rect 11758 1888 11844 1944
rect 11900 1888 11970 1944
rect 11630 1802 11970 1888
rect 11630 1746 11702 1802
rect 11758 1746 11844 1802
rect 11900 1746 11970 1802
rect 11630 1660 11970 1746
rect 11630 1604 11702 1660
rect 11758 1604 11844 1660
rect 11900 1604 11970 1660
rect 11630 1518 11970 1604
rect 11630 1462 11702 1518
rect 11758 1462 11844 1518
rect 11900 1462 11970 1518
rect 11630 1376 11970 1462
rect 11630 1320 11702 1376
rect 11758 1320 11844 1376
rect 11900 1320 11970 1376
rect 11630 1234 11970 1320
rect 11630 1178 11702 1234
rect 11758 1178 11844 1234
rect 11900 1178 11970 1234
rect 11630 1092 11970 1178
rect 11630 1036 11702 1092
rect 11758 1036 11844 1092
rect 11900 1036 11970 1092
rect 11630 950 11970 1036
rect 11630 894 11702 950
rect 11758 894 11844 950
rect 11900 894 11970 950
rect 11630 808 11970 894
rect 11630 752 11702 808
rect 11758 752 11844 808
rect 11900 752 11970 808
rect 11630 666 11970 752
rect 11630 610 11702 666
rect 11758 610 11844 666
rect 11900 610 11970 666
rect 11630 524 11970 610
rect 11630 468 11702 524
rect 11758 468 11844 524
rect 11900 468 11970 524
rect 11630 458 11970 468
rect 12400 12302 12526 12320
rect 12582 12302 12650 12358
rect 12706 12302 12774 12358
rect 12830 12302 12898 12358
rect 12954 12302 13022 12358
rect 13078 12302 13200 12358
rect 12400 12234 13200 12302
rect 12400 12178 12526 12234
rect 12582 12178 12650 12234
rect 12706 12178 12774 12234
rect 12830 12178 12898 12234
rect 12954 12178 13022 12234
rect 13078 12178 13200 12234
rect 12400 12110 13200 12178
rect 12400 12054 12526 12110
rect 12582 12054 12650 12110
rect 12706 12054 12774 12110
rect 12830 12054 12898 12110
rect 12954 12054 13022 12110
rect 13078 12054 13200 12110
rect 12400 11986 13200 12054
rect 12400 11930 12526 11986
rect 12582 11930 12650 11986
rect 12706 11930 12774 11986
rect 12830 11930 12898 11986
rect 12954 11930 13022 11986
rect 13078 11930 13200 11986
rect 12400 11862 13200 11930
rect 12400 11806 12526 11862
rect 12582 11806 12650 11862
rect 12706 11806 12774 11862
rect 12830 11806 12898 11862
rect 12954 11806 13022 11862
rect 13078 11806 13200 11862
rect 12400 11738 13200 11806
rect 12400 11682 12526 11738
rect 12582 11682 12650 11738
rect 12706 11682 12774 11738
rect 12830 11682 12898 11738
rect 12954 11682 13022 11738
rect 13078 11682 13200 11738
rect 12400 11614 13200 11682
rect 12400 11558 12526 11614
rect 12582 11558 12650 11614
rect 12706 11558 12774 11614
rect 12830 11558 12898 11614
rect 12954 11558 13022 11614
rect 13078 11558 13200 11614
rect 12400 11490 13200 11558
rect 12400 11434 12526 11490
rect 12582 11434 12650 11490
rect 12706 11434 12774 11490
rect 12830 11434 12898 11490
rect 12954 11434 13022 11490
rect 13078 11434 13200 11490
rect 12400 11366 13200 11434
rect 12400 11310 12526 11366
rect 12582 11310 12650 11366
rect 12706 11310 12774 11366
rect 12830 11310 12898 11366
rect 12954 11310 13022 11366
rect 13078 11310 13200 11366
rect 12400 11242 13200 11310
rect 12400 11186 12526 11242
rect 12582 11186 12650 11242
rect 12706 11186 12774 11242
rect 12830 11186 12898 11242
rect 12954 11186 13022 11242
rect 13078 11186 13200 11242
rect 12400 11118 13200 11186
rect 12400 11062 12526 11118
rect 12582 11062 12650 11118
rect 12706 11062 12774 11118
rect 12830 11062 12898 11118
rect 12954 11062 13022 11118
rect 13078 11062 13200 11118
rect 12400 10994 13200 11062
rect 12400 10938 12526 10994
rect 12582 10938 12650 10994
rect 12706 10938 12774 10994
rect 12830 10938 12898 10994
rect 12954 10938 13022 10994
rect 13078 10938 13200 10994
rect 12400 10870 13200 10938
rect 12400 10814 12526 10870
rect 12582 10814 12650 10870
rect 12706 10814 12774 10870
rect 12830 10814 12898 10870
rect 12954 10814 13022 10870
rect 13078 10814 13200 10870
rect 12400 10746 13200 10814
rect 12400 10690 12526 10746
rect 12582 10690 12650 10746
rect 12706 10690 12774 10746
rect 12830 10690 12898 10746
rect 12954 10690 13022 10746
rect 13078 10690 13200 10746
rect 12400 10622 13200 10690
rect 12400 10566 12526 10622
rect 12582 10566 12650 10622
rect 12706 10566 12774 10622
rect 12830 10566 12898 10622
rect 12954 10566 13022 10622
rect 13078 10566 13200 10622
rect 12400 10498 13200 10566
rect 12400 10442 12526 10498
rect 12582 10442 12650 10498
rect 12706 10442 12774 10498
rect 12830 10442 12898 10498
rect 12954 10442 13022 10498
rect 13078 10442 13200 10498
rect 12400 10374 13200 10442
rect 12400 10318 12526 10374
rect 12582 10318 12650 10374
rect 12706 10318 12774 10374
rect 12830 10318 12898 10374
rect 12954 10318 13022 10374
rect 13078 10318 13200 10374
rect 12400 10250 13200 10318
rect 12400 10194 12526 10250
rect 12582 10194 12650 10250
rect 12706 10194 12774 10250
rect 12830 10194 12898 10250
rect 12954 10194 13022 10250
rect 13078 10194 13200 10250
rect 12400 10126 13200 10194
rect 12400 10070 12526 10126
rect 12582 10070 12650 10126
rect 12706 10070 12774 10126
rect 12830 10070 12898 10126
rect 12954 10070 13022 10126
rect 13078 10070 13200 10126
rect 12400 10002 13200 10070
rect 12400 9946 12526 10002
rect 12582 9946 12650 10002
rect 12706 9946 12774 10002
rect 12830 9946 12898 10002
rect 12954 9946 13022 10002
rect 13078 9946 13200 10002
rect 12400 9878 13200 9946
rect 12400 9822 12526 9878
rect 12582 9822 12650 9878
rect 12706 9822 12774 9878
rect 12830 9822 12898 9878
rect 12954 9822 13022 9878
rect 13078 9822 13200 9878
rect 12400 9754 13200 9822
rect 12400 9698 12526 9754
rect 12582 9698 12650 9754
rect 12706 9698 12774 9754
rect 12830 9698 12898 9754
rect 12954 9698 13022 9754
rect 13078 9698 13200 9754
rect 12400 9630 13200 9698
rect 12400 9574 12526 9630
rect 12582 9574 12650 9630
rect 12706 9574 12774 9630
rect 12830 9574 12898 9630
rect 12954 9574 13022 9630
rect 13078 9574 13200 9630
rect 12400 9506 13200 9574
rect 12400 9450 12526 9506
rect 12582 9450 12650 9506
rect 12706 9450 12774 9506
rect 12830 9450 12898 9506
rect 12954 9450 13022 9506
rect 13078 9450 13200 9506
rect 12400 9382 13200 9450
rect 12400 9326 12526 9382
rect 12582 9326 12650 9382
rect 12706 9326 12774 9382
rect 12830 9326 12898 9382
rect 12954 9326 13022 9382
rect 13078 9326 13200 9382
rect 12400 9258 13200 9326
rect 12400 9202 12526 9258
rect 12582 9202 12650 9258
rect 12706 9202 12774 9258
rect 12830 9202 12898 9258
rect 12954 9202 13022 9258
rect 13078 9202 13200 9258
rect 12400 9134 13200 9202
rect 12400 9078 12526 9134
rect 12582 9078 12650 9134
rect 12706 9078 12774 9134
rect 12830 9078 12898 9134
rect 12954 9078 13022 9134
rect 13078 9078 13200 9134
rect 12400 9010 13200 9078
rect 12400 8954 12526 9010
rect 12582 8954 12650 9010
rect 12706 8954 12774 9010
rect 12830 8954 12898 9010
rect 12954 8954 13022 9010
rect 13078 8954 13200 9010
rect 12400 8886 13200 8954
rect 12400 8830 12526 8886
rect 12582 8830 12650 8886
rect 12706 8830 12774 8886
rect 12830 8830 12898 8886
rect 12954 8830 13022 8886
rect 13078 8830 13200 8886
rect 12400 8762 13200 8830
rect 12400 8706 12526 8762
rect 12582 8706 12650 8762
rect 12706 8706 12774 8762
rect 12830 8706 12898 8762
rect 12954 8706 13022 8762
rect 13078 8706 13200 8762
rect 12400 8638 13200 8706
rect 12400 8582 12526 8638
rect 12582 8582 12650 8638
rect 12706 8582 12774 8638
rect 12830 8582 12898 8638
rect 12954 8582 13022 8638
rect 13078 8582 13200 8638
rect 12400 8514 13200 8582
rect 12400 8458 12526 8514
rect 12582 8458 12650 8514
rect 12706 8458 12774 8514
rect 12830 8458 12898 8514
rect 12954 8458 13022 8514
rect 13078 8458 13200 8514
rect 12400 8390 13200 8458
rect 12400 8334 12526 8390
rect 12582 8334 12650 8390
rect 12706 8334 12774 8390
rect 12830 8334 12898 8390
rect 12954 8334 13022 8390
rect 13078 8334 13200 8390
rect 12400 8266 13200 8334
rect 12400 8210 12526 8266
rect 12582 8210 12650 8266
rect 12706 8210 12774 8266
rect 12830 8210 12898 8266
rect 12954 8210 13022 8266
rect 13078 8210 13200 8266
rect 12400 8142 13200 8210
rect 12400 8086 12526 8142
rect 12582 8086 12650 8142
rect 12706 8086 12774 8142
rect 12830 8086 12898 8142
rect 12954 8086 13022 8142
rect 13078 8086 13200 8142
rect 12400 8018 13200 8086
rect 12400 7962 12526 8018
rect 12582 7962 12650 8018
rect 12706 7962 12774 8018
rect 12830 7962 12898 8018
rect 12954 7962 13022 8018
rect 13078 7962 13200 8018
rect 12400 7894 13200 7962
rect 12400 7838 12526 7894
rect 12582 7838 12650 7894
rect 12706 7838 12774 7894
rect 12830 7838 12898 7894
rect 12954 7838 13022 7894
rect 13078 7838 13200 7894
rect 12400 7770 13200 7838
rect 12400 7714 12526 7770
rect 12582 7714 12650 7770
rect 12706 7714 12774 7770
rect 12830 7714 12898 7770
rect 12954 7714 13022 7770
rect 13078 7714 13200 7770
rect 12400 7646 13200 7714
rect 12400 7590 12526 7646
rect 12582 7590 12650 7646
rect 12706 7590 12774 7646
rect 12830 7590 12898 7646
rect 12954 7590 13022 7646
rect 13078 7590 13200 7646
rect 12400 7522 13200 7590
rect 12400 7466 12526 7522
rect 12582 7466 12650 7522
rect 12706 7466 12774 7522
rect 12830 7466 12898 7522
rect 12954 7466 13022 7522
rect 13078 7466 13200 7522
rect 12400 7398 13200 7466
rect 12400 7342 12526 7398
rect 12582 7342 12650 7398
rect 12706 7342 12774 7398
rect 12830 7342 12898 7398
rect 12954 7342 13022 7398
rect 13078 7342 13200 7398
rect 12400 7274 13200 7342
rect 12400 7218 12526 7274
rect 12582 7218 12650 7274
rect 12706 7218 12774 7274
rect 12830 7218 12898 7274
rect 12954 7218 13022 7274
rect 13078 7218 13200 7274
rect 12400 7150 13200 7218
rect 12400 7094 12526 7150
rect 12582 7094 12650 7150
rect 12706 7094 12774 7150
rect 12830 7094 12898 7150
rect 12954 7094 13022 7150
rect 13078 7094 13200 7150
rect 12400 7026 13200 7094
rect 12400 6970 12526 7026
rect 12582 6970 12650 7026
rect 12706 6970 12774 7026
rect 12830 6970 12898 7026
rect 12954 6970 13022 7026
rect 13078 6970 13200 7026
rect 12400 6902 13200 6970
rect 12400 6846 12526 6902
rect 12582 6846 12650 6902
rect 12706 6846 12774 6902
rect 12830 6846 12898 6902
rect 12954 6846 13022 6902
rect 13078 6846 13200 6902
rect 12400 6778 13200 6846
rect 12400 6722 12526 6778
rect 12582 6722 12650 6778
rect 12706 6722 12774 6778
rect 12830 6722 12898 6778
rect 12954 6722 13022 6778
rect 13078 6722 13200 6778
rect 12400 6654 13200 6722
rect 12400 6598 12526 6654
rect 12582 6598 12650 6654
rect 12706 6598 12774 6654
rect 12830 6598 12898 6654
rect 12954 6598 13022 6654
rect 13078 6598 13200 6654
rect 12400 6530 13200 6598
rect 12400 6474 12526 6530
rect 12582 6474 12650 6530
rect 12706 6474 12774 6530
rect 12830 6474 12898 6530
rect 12954 6474 13022 6530
rect 13078 6474 13200 6530
rect 12400 6406 13200 6474
rect 12400 6350 12526 6406
rect 12582 6350 12650 6406
rect 12706 6350 12774 6406
rect 12830 6350 12898 6406
rect 12954 6350 13022 6406
rect 13078 6350 13200 6406
rect 12400 6282 13200 6350
rect 12400 6226 12526 6282
rect 12582 6226 12650 6282
rect 12706 6226 12774 6282
rect 12830 6226 12898 6282
rect 12954 6226 13022 6282
rect 13078 6226 13200 6282
rect 12400 6158 13200 6226
rect 12400 6102 12526 6158
rect 12582 6102 12650 6158
rect 12706 6102 12774 6158
rect 12830 6102 12898 6158
rect 12954 6102 13022 6158
rect 13078 6102 13200 6158
rect 12400 6034 13200 6102
rect 12400 5978 12526 6034
rect 12582 5978 12650 6034
rect 12706 5978 12774 6034
rect 12830 5978 12898 6034
rect 12954 5978 13022 6034
rect 13078 5978 13200 6034
rect 12400 5910 13200 5978
rect 12400 5854 12526 5910
rect 12582 5854 12650 5910
rect 12706 5854 12774 5910
rect 12830 5854 12898 5910
rect 12954 5854 13022 5910
rect 13078 5854 13200 5910
rect 12400 5786 13200 5854
rect 12400 5730 12526 5786
rect 12582 5730 12650 5786
rect 12706 5730 12774 5786
rect 12830 5730 12898 5786
rect 12954 5730 13022 5786
rect 13078 5730 13200 5786
rect 12400 5662 13200 5730
rect 12400 5606 12526 5662
rect 12582 5606 12650 5662
rect 12706 5606 12774 5662
rect 12830 5606 12898 5662
rect 12954 5606 13022 5662
rect 13078 5606 13200 5662
rect 12400 5538 13200 5606
rect 12400 5482 12526 5538
rect 12582 5482 12650 5538
rect 12706 5482 12774 5538
rect 12830 5482 12898 5538
rect 12954 5482 13022 5538
rect 13078 5482 13200 5538
rect 12400 5414 13200 5482
rect 12400 5358 12526 5414
rect 12582 5358 12650 5414
rect 12706 5358 12774 5414
rect 12830 5358 12898 5414
rect 12954 5358 13022 5414
rect 13078 5358 13200 5414
rect 12400 5290 13200 5358
rect 12400 5234 12526 5290
rect 12582 5234 12650 5290
rect 12706 5234 12774 5290
rect 12830 5234 12898 5290
rect 12954 5234 13022 5290
rect 13078 5234 13200 5290
rect 12400 5166 13200 5234
rect 12400 5110 12526 5166
rect 12582 5110 12650 5166
rect 12706 5110 12774 5166
rect 12830 5110 12898 5166
rect 12954 5110 13022 5166
rect 13078 5110 13200 5166
rect 12400 5042 13200 5110
rect 12400 4986 12526 5042
rect 12582 4986 12650 5042
rect 12706 4986 12774 5042
rect 12830 4986 12898 5042
rect 12954 4986 13022 5042
rect 13078 4986 13200 5042
rect 12400 4918 13200 4986
rect 12400 4862 12526 4918
rect 12582 4862 12650 4918
rect 12706 4862 12774 4918
rect 12830 4862 12898 4918
rect 12954 4862 13022 4918
rect 13078 4862 13200 4918
rect 12400 4794 13200 4862
rect 12400 4738 12526 4794
rect 12582 4738 12650 4794
rect 12706 4738 12774 4794
rect 12830 4738 12898 4794
rect 12954 4738 13022 4794
rect 13078 4738 13200 4794
rect 12400 4670 13200 4738
rect 12400 4614 12526 4670
rect 12582 4614 12650 4670
rect 12706 4614 12774 4670
rect 12830 4614 12898 4670
rect 12954 4614 13022 4670
rect 13078 4614 13200 4670
rect 12400 4546 13200 4614
rect 12400 4490 12526 4546
rect 12582 4490 12650 4546
rect 12706 4490 12774 4546
rect 12830 4490 12898 4546
rect 12954 4490 13022 4546
rect 13078 4490 13200 4546
rect 12400 4422 13200 4490
rect 12400 4366 12526 4422
rect 12582 4366 12650 4422
rect 12706 4366 12774 4422
rect 12830 4366 12898 4422
rect 12954 4366 13022 4422
rect 13078 4366 13200 4422
rect 12400 4298 13200 4366
rect 12400 4242 12526 4298
rect 12582 4242 12650 4298
rect 12706 4242 12774 4298
rect 12830 4242 12898 4298
rect 12954 4242 13022 4298
rect 13078 4242 13200 4298
rect 12400 4174 13200 4242
rect 12400 4118 12526 4174
rect 12582 4118 12650 4174
rect 12706 4118 12774 4174
rect 12830 4118 12898 4174
rect 12954 4118 13022 4174
rect 13078 4118 13200 4174
rect 12400 4050 13200 4118
rect 12400 3994 12526 4050
rect 12582 3994 12650 4050
rect 12706 3994 12774 4050
rect 12830 3994 12898 4050
rect 12954 3994 13022 4050
rect 13078 3994 13200 4050
rect 12400 3926 13200 3994
rect 12400 3870 12526 3926
rect 12582 3870 12650 3926
rect 12706 3870 12774 3926
rect 12830 3870 12898 3926
rect 12954 3870 13022 3926
rect 13078 3870 13200 3926
rect 12400 3802 13200 3870
rect 12400 3746 12526 3802
rect 12582 3746 12650 3802
rect 12706 3746 12774 3802
rect 12830 3746 12898 3802
rect 12954 3746 13022 3802
rect 13078 3746 13200 3802
rect 12400 3678 13200 3746
rect 12400 3622 12526 3678
rect 12582 3622 12650 3678
rect 12706 3622 12774 3678
rect 12830 3622 12898 3678
rect 12954 3622 13022 3678
rect 13078 3622 13200 3678
rect 12400 3554 13200 3622
rect 12400 3498 12526 3554
rect 12582 3498 12650 3554
rect 12706 3498 12774 3554
rect 12830 3498 12898 3554
rect 12954 3498 13022 3554
rect 13078 3498 13200 3554
rect 12400 3430 13200 3498
rect 12400 3374 12526 3430
rect 12582 3374 12650 3430
rect 12706 3374 12774 3430
rect 12830 3374 12898 3430
rect 12954 3374 13022 3430
rect 13078 3374 13200 3430
rect 12400 3306 13200 3374
rect 12400 3250 12526 3306
rect 12582 3250 12650 3306
rect 12706 3250 12774 3306
rect 12830 3250 12898 3306
rect 12954 3250 13022 3306
rect 13078 3250 13200 3306
rect 12400 3182 13200 3250
rect 12400 3126 12526 3182
rect 12582 3126 12650 3182
rect 12706 3126 12774 3182
rect 12830 3126 12898 3182
rect 12954 3126 13022 3182
rect 13078 3126 13200 3182
rect 12400 3058 13200 3126
rect 12400 3002 12526 3058
rect 12582 3002 12650 3058
rect 12706 3002 12774 3058
rect 12830 3002 12898 3058
rect 12954 3002 13022 3058
rect 13078 3002 13200 3058
rect 12400 2934 13200 3002
rect 12400 2878 12526 2934
rect 12582 2878 12650 2934
rect 12706 2878 12774 2934
rect 12830 2878 12898 2934
rect 12954 2878 13022 2934
rect 13078 2878 13200 2934
rect 12400 2810 13200 2878
rect 12400 2754 12526 2810
rect 12582 2754 12650 2810
rect 12706 2754 12774 2810
rect 12830 2754 12898 2810
rect 12954 2754 13022 2810
rect 13078 2754 13200 2810
rect 12400 2686 13200 2754
rect 12400 2630 12526 2686
rect 12582 2630 12650 2686
rect 12706 2630 12774 2686
rect 12830 2630 12898 2686
rect 12954 2630 13022 2686
rect 13078 2630 13200 2686
rect 12400 2562 13200 2630
rect 12400 2506 12526 2562
rect 12582 2506 12650 2562
rect 12706 2506 12774 2562
rect 12830 2506 12898 2562
rect 12954 2506 13022 2562
rect 13078 2506 13200 2562
rect 12400 2438 13200 2506
rect 12400 2382 12526 2438
rect 12582 2382 12650 2438
rect 12706 2382 12774 2438
rect 12830 2382 12898 2438
rect 12954 2382 13022 2438
rect 13078 2382 13200 2438
rect 12400 2314 13200 2382
rect 12400 2258 12526 2314
rect 12582 2258 12650 2314
rect 12706 2258 12774 2314
rect 12830 2258 12898 2314
rect 12954 2258 13022 2314
rect 13078 2258 13200 2314
rect 12400 2190 13200 2258
rect 12400 2134 12526 2190
rect 12582 2134 12650 2190
rect 12706 2134 12774 2190
rect 12830 2134 12898 2190
rect 12954 2134 13022 2190
rect 13078 2134 13200 2190
rect 12400 2066 13200 2134
rect 12400 2010 12526 2066
rect 12582 2010 12650 2066
rect 12706 2010 12774 2066
rect 12830 2010 12898 2066
rect 12954 2010 13022 2066
rect 13078 2010 13200 2066
rect 12400 1942 13200 2010
rect 12400 1886 12526 1942
rect 12582 1886 12650 1942
rect 12706 1886 12774 1942
rect 12830 1886 12898 1942
rect 12954 1886 13022 1942
rect 13078 1886 13200 1942
rect 12400 1818 13200 1886
rect 12400 1762 12526 1818
rect 12582 1762 12650 1818
rect 12706 1762 12774 1818
rect 12830 1762 12898 1818
rect 12954 1762 13022 1818
rect 13078 1762 13200 1818
rect 12400 1694 13200 1762
rect 12400 1638 12526 1694
rect 12582 1638 12650 1694
rect 12706 1638 12774 1694
rect 12830 1638 12898 1694
rect 12954 1638 13022 1694
rect 13078 1638 13200 1694
rect 12400 1570 13200 1638
rect 12400 1514 12526 1570
rect 12582 1514 12650 1570
rect 12706 1514 12774 1570
rect 12830 1514 12898 1570
rect 12954 1514 13022 1570
rect 13078 1514 13200 1570
rect 12400 1446 13200 1514
rect 12400 1390 12526 1446
rect 12582 1390 12650 1446
rect 12706 1390 12774 1446
rect 12830 1390 12898 1446
rect 12954 1390 13022 1446
rect 13078 1390 13200 1446
rect 12400 1322 13200 1390
rect 12400 1266 12526 1322
rect 12582 1266 12650 1322
rect 12706 1266 12774 1322
rect 12830 1266 12898 1322
rect 12954 1266 13022 1322
rect 13078 1266 13200 1322
rect 12400 1198 13200 1266
rect 12400 1142 12526 1198
rect 12582 1142 12650 1198
rect 12706 1142 12774 1198
rect 12830 1142 12898 1198
rect 12954 1142 13022 1198
rect 13078 1142 13200 1198
rect 12400 1074 13200 1142
rect 12400 1018 12526 1074
rect 12582 1018 12650 1074
rect 12706 1018 12774 1074
rect 12830 1018 12898 1074
rect 12954 1018 13022 1074
rect 13078 1018 13200 1074
rect 12400 950 13200 1018
rect 12400 894 12526 950
rect 12582 894 12650 950
rect 12706 894 12774 950
rect 12830 894 12898 950
rect 12954 894 13022 950
rect 13078 894 13200 950
rect 12400 826 13200 894
rect 12400 770 12526 826
rect 12582 770 12650 826
rect 12706 770 12774 826
rect 12830 770 12898 826
rect 12954 770 13022 826
rect 13078 770 13200 826
rect 12400 702 13200 770
rect 12400 646 12526 702
rect 12582 646 12650 702
rect 12706 646 12774 702
rect 12830 646 12898 702
rect 12954 646 13022 702
rect 13078 646 13200 702
rect 12400 578 13200 646
rect 12400 522 12526 578
rect 12582 522 12650 578
rect 12706 522 12774 578
rect 12830 522 12898 578
rect 12954 522 13022 578
rect 13078 522 13200 578
rect 12400 458 13200 522
rect -400 454 13200 458
rect -400 398 -286 454
rect -230 398 -162 454
rect -106 398 -38 454
rect 18 398 86 454
rect 142 398 210 454
rect 266 398 12526 454
rect 12582 398 12650 454
rect 12706 398 12774 454
rect 12830 398 12898 454
rect 12954 398 13022 454
rect 13078 398 13200 454
rect -400 330 13200 398
rect -400 274 -286 330
rect -230 274 -162 330
rect -106 274 -38 330
rect 18 274 86 330
rect 142 274 210 330
rect 266 302 12526 330
rect 266 274 415 302
rect -400 246 415 274
rect 471 246 557 302
rect 613 246 699 302
rect 755 246 841 302
rect 897 246 983 302
rect 1039 246 1125 302
rect 1181 246 1267 302
rect 1323 246 1409 302
rect 1465 246 1551 302
rect 1607 246 1693 302
rect 1749 246 1835 302
rect 1891 246 1977 302
rect 2033 246 2119 302
rect 2175 246 2261 302
rect 2317 246 2403 302
rect 2459 246 2545 302
rect 2601 246 2687 302
rect 2743 246 2829 302
rect 2885 246 2971 302
rect 3027 246 3113 302
rect 3169 246 3255 302
rect 3311 246 3397 302
rect 3453 246 3539 302
rect 3595 246 3681 302
rect 3737 246 3823 302
rect 3879 246 3965 302
rect 4021 246 4107 302
rect 4163 246 4249 302
rect 4305 246 4391 302
rect 4447 246 4533 302
rect 4589 246 4675 302
rect 4731 246 4817 302
rect 4873 246 4959 302
rect 5015 246 5101 302
rect 5157 246 5243 302
rect 5299 246 5385 302
rect 5441 246 5527 302
rect 5583 246 5669 302
rect 5725 246 5811 302
rect 5867 246 5953 302
rect 6009 246 6095 302
rect 6151 246 6237 302
rect 6293 246 6379 302
rect 6435 246 6521 302
rect 6577 246 6663 302
rect 6719 246 6805 302
rect 6861 246 6947 302
rect 7003 246 7089 302
rect 7145 246 7231 302
rect 7287 246 7373 302
rect 7429 246 7515 302
rect 7571 246 7657 302
rect 7713 246 7799 302
rect 7855 246 7941 302
rect 7997 246 8083 302
rect 8139 246 8225 302
rect 8281 246 8367 302
rect 8423 246 8509 302
rect 8565 246 8651 302
rect 8707 246 8793 302
rect 8849 246 8935 302
rect 8991 246 9077 302
rect 9133 246 9219 302
rect 9275 246 9361 302
rect 9417 246 9503 302
rect 9559 246 9645 302
rect 9701 246 9787 302
rect 9843 246 9929 302
rect 9985 246 10071 302
rect 10127 246 10213 302
rect 10269 246 10355 302
rect 10411 246 10497 302
rect 10553 246 10639 302
rect 10695 246 10781 302
rect 10837 246 10923 302
rect 10979 246 11065 302
rect 11121 246 11207 302
rect 11263 246 11349 302
rect 11405 246 11491 302
rect 11547 246 11633 302
rect 11689 246 11775 302
rect 11831 246 11917 302
rect 11973 246 12059 302
rect 12115 246 12201 302
rect 12257 246 12343 302
rect 12399 274 12526 302
rect 12582 274 12650 330
rect 12706 274 12774 330
rect 12830 274 12898 330
rect 12954 274 13022 330
rect 13078 274 13200 330
rect 12399 246 13200 274
rect -400 206 13200 246
rect -400 150 -286 206
rect -230 150 -162 206
rect -106 150 -38 206
rect 18 150 86 206
rect 142 150 210 206
rect 266 160 12526 206
rect 266 150 415 160
rect -400 104 415 150
rect 471 104 557 160
rect 613 104 699 160
rect 755 104 841 160
rect 897 104 983 160
rect 1039 104 1125 160
rect 1181 104 1267 160
rect 1323 104 1409 160
rect 1465 104 1551 160
rect 1607 104 1693 160
rect 1749 104 1835 160
rect 1891 104 1977 160
rect 2033 104 2119 160
rect 2175 104 2261 160
rect 2317 104 2403 160
rect 2459 104 2545 160
rect 2601 104 2687 160
rect 2743 104 2829 160
rect 2885 104 2971 160
rect 3027 104 3113 160
rect 3169 104 3255 160
rect 3311 104 3397 160
rect 3453 104 3539 160
rect 3595 104 3681 160
rect 3737 104 3823 160
rect 3879 104 3965 160
rect 4021 104 4107 160
rect 4163 104 4249 160
rect 4305 104 4391 160
rect 4447 104 4533 160
rect 4589 104 4675 160
rect 4731 104 4817 160
rect 4873 104 4959 160
rect 5015 104 5101 160
rect 5157 104 5243 160
rect 5299 104 5385 160
rect 5441 104 5527 160
rect 5583 104 5669 160
rect 5725 104 5811 160
rect 5867 104 5953 160
rect 6009 104 6095 160
rect 6151 104 6237 160
rect 6293 104 6379 160
rect 6435 104 6521 160
rect 6577 104 6663 160
rect 6719 104 6805 160
rect 6861 104 6947 160
rect 7003 104 7089 160
rect 7145 104 7231 160
rect 7287 104 7373 160
rect 7429 104 7515 160
rect 7571 104 7657 160
rect 7713 104 7799 160
rect 7855 104 7941 160
rect 7997 104 8083 160
rect 8139 104 8225 160
rect 8281 104 8367 160
rect 8423 104 8509 160
rect 8565 104 8651 160
rect 8707 104 8793 160
rect 8849 104 8935 160
rect 8991 104 9077 160
rect 9133 104 9219 160
rect 9275 104 9361 160
rect 9417 104 9503 160
rect 9559 104 9645 160
rect 9701 104 9787 160
rect 9843 104 9929 160
rect 9985 104 10071 160
rect 10127 104 10213 160
rect 10269 104 10355 160
rect 10411 104 10497 160
rect 10553 104 10639 160
rect 10695 104 10781 160
rect 10837 104 10923 160
rect 10979 104 11065 160
rect 11121 104 11207 160
rect 11263 104 11349 160
rect 11405 104 11491 160
rect 11547 104 11633 160
rect 11689 104 11775 160
rect 11831 104 11917 160
rect 11973 104 12059 160
rect 12115 104 12201 160
rect 12257 104 12343 160
rect 12399 150 12526 160
rect 12582 150 12650 206
rect 12706 150 12774 206
rect 12830 150 12898 206
rect 12954 150 13022 206
rect 13078 150 13200 206
rect 12399 104 13200 150
rect -400 0 13200 104
<< via3 >>
rect -254 12893 -198 12949
rect -130 12893 -74 12949
rect -6 12893 50 12949
rect 118 12893 174 12949
rect 242 12893 298 12949
rect 366 12893 422 12949
rect 490 12893 546 12949
rect 614 12893 670 12949
rect 738 12893 794 12949
rect 862 12893 918 12949
rect 986 12893 1042 12949
rect 1110 12893 1166 12949
rect 1234 12893 1290 12949
rect 1358 12893 1414 12949
rect 1482 12893 1538 12949
rect 1606 12893 1662 12949
rect 1730 12893 1786 12949
rect 1854 12893 1910 12949
rect 1978 12893 2034 12949
rect 2102 12893 2158 12949
rect 2226 12893 2282 12949
rect 2350 12893 2406 12949
rect 2474 12893 2530 12949
rect 2598 12893 2654 12949
rect 2722 12893 2778 12949
rect 2846 12893 2902 12949
rect 2970 12893 3026 12949
rect 3094 12893 3150 12949
rect 3218 12893 3274 12949
rect 3342 12893 3398 12949
rect 3466 12893 3522 12949
rect 3590 12893 3646 12949
rect 3714 12893 3770 12949
rect 3838 12893 3894 12949
rect 3962 12893 4018 12949
rect 4086 12893 4142 12949
rect 4210 12893 4266 12949
rect 4334 12893 4390 12949
rect 4458 12893 4514 12949
rect 4582 12893 4638 12949
rect 4706 12893 4762 12949
rect 4830 12893 4886 12949
rect 4954 12893 5010 12949
rect 5078 12893 5134 12949
rect 5202 12893 5258 12949
rect 5326 12893 5382 12949
rect 5450 12893 5506 12949
rect 5574 12893 5630 12949
rect 5698 12893 5754 12949
rect 5822 12893 5878 12949
rect 5946 12893 6002 12949
rect 6070 12893 6126 12949
rect 6194 12893 6250 12949
rect 6318 12893 6374 12949
rect 6442 12893 6498 12949
rect 6566 12893 6622 12949
rect 6690 12893 6746 12949
rect 6814 12893 6870 12949
rect 6938 12893 6994 12949
rect 7062 12893 7118 12949
rect 7186 12893 7242 12949
rect 7310 12893 7366 12949
rect 7434 12893 7490 12949
rect 7558 12893 7614 12949
rect 7682 12893 7738 12949
rect 7806 12893 7862 12949
rect 7930 12893 7986 12949
rect 8054 12893 8110 12949
rect 8178 12893 8234 12949
rect 8302 12893 8358 12949
rect 8426 12893 8482 12949
rect 8550 12893 8606 12949
rect 8674 12893 8730 12949
rect 8798 12893 8854 12949
rect 8922 12893 8978 12949
rect 9046 12893 9102 12949
rect 9170 12893 9226 12949
rect 9294 12893 9350 12949
rect 9418 12893 9474 12949
rect 9542 12893 9598 12949
rect 9666 12893 9722 12949
rect 9790 12893 9846 12949
rect 9914 12893 9970 12949
rect 10038 12893 10094 12949
rect 10162 12893 10218 12949
rect 10286 12893 10342 12949
rect 10410 12893 10466 12949
rect 10534 12893 10590 12949
rect 10658 12893 10714 12949
rect 10782 12893 10838 12949
rect 10906 12893 10962 12949
rect 11030 12893 11086 12949
rect 11154 12893 11210 12949
rect 11278 12893 11334 12949
rect 11402 12893 11458 12949
rect 11526 12893 11582 12949
rect 11650 12893 11706 12949
rect 11774 12893 11830 12949
rect 11898 12893 11954 12949
rect 12022 12893 12078 12949
rect 12146 12893 12202 12949
rect 12270 12893 12326 12949
rect 12394 12893 12450 12949
rect 12518 12893 12574 12949
rect 12642 12893 12698 12949
rect 12766 12893 12822 12949
rect 12890 12893 12946 12949
rect 13014 12893 13070 12949
rect -254 12769 -198 12825
rect -130 12769 -74 12825
rect -6 12769 50 12825
rect 118 12769 174 12825
rect 242 12769 298 12825
rect 366 12769 422 12825
rect 490 12769 546 12825
rect 614 12769 670 12825
rect 738 12769 794 12825
rect 862 12769 918 12825
rect 986 12769 1042 12825
rect 1110 12769 1166 12825
rect 1234 12769 1290 12825
rect 1358 12769 1414 12825
rect 1482 12769 1538 12825
rect 1606 12769 1662 12825
rect 1730 12769 1786 12825
rect 1854 12769 1910 12825
rect 1978 12769 2034 12825
rect 2102 12769 2158 12825
rect 2226 12769 2282 12825
rect 2350 12769 2406 12825
rect 2474 12769 2530 12825
rect 2598 12769 2654 12825
rect 2722 12769 2778 12825
rect 2846 12769 2902 12825
rect 2970 12769 3026 12825
rect 3094 12769 3150 12825
rect 3218 12769 3274 12825
rect 3342 12769 3398 12825
rect 3466 12769 3522 12825
rect 3590 12769 3646 12825
rect 3714 12769 3770 12825
rect 3838 12769 3894 12825
rect 3962 12769 4018 12825
rect 4086 12769 4142 12825
rect 4210 12769 4266 12825
rect 4334 12769 4390 12825
rect 4458 12769 4514 12825
rect 4582 12769 4638 12825
rect 4706 12769 4762 12825
rect 4830 12769 4886 12825
rect 4954 12769 5010 12825
rect 5078 12769 5134 12825
rect 5202 12769 5258 12825
rect 5326 12769 5382 12825
rect 5450 12769 5506 12825
rect 5574 12769 5630 12825
rect 5698 12769 5754 12825
rect 5822 12769 5878 12825
rect 5946 12769 6002 12825
rect 6070 12769 6126 12825
rect 6194 12769 6250 12825
rect 6318 12769 6374 12825
rect 6442 12769 6498 12825
rect 6566 12769 6622 12825
rect 6690 12769 6746 12825
rect 6814 12769 6870 12825
rect 6938 12769 6994 12825
rect 7062 12769 7118 12825
rect 7186 12769 7242 12825
rect 7310 12769 7366 12825
rect 7434 12769 7490 12825
rect 7558 12769 7614 12825
rect 7682 12769 7738 12825
rect 7806 12769 7862 12825
rect 7930 12769 7986 12825
rect 8054 12769 8110 12825
rect 8178 12769 8234 12825
rect 8302 12769 8358 12825
rect 8426 12769 8482 12825
rect 8550 12769 8606 12825
rect 8674 12769 8730 12825
rect 8798 12769 8854 12825
rect 8922 12769 8978 12825
rect 9046 12769 9102 12825
rect 9170 12769 9226 12825
rect 9294 12769 9350 12825
rect 9418 12769 9474 12825
rect 9542 12769 9598 12825
rect 9666 12769 9722 12825
rect 9790 12769 9846 12825
rect 9914 12769 9970 12825
rect 10038 12769 10094 12825
rect 10162 12769 10218 12825
rect 10286 12769 10342 12825
rect 10410 12769 10466 12825
rect 10534 12769 10590 12825
rect 10658 12769 10714 12825
rect 10782 12769 10838 12825
rect 10906 12769 10962 12825
rect 11030 12769 11086 12825
rect 11154 12769 11210 12825
rect 11278 12769 11334 12825
rect 11402 12769 11458 12825
rect 11526 12769 11582 12825
rect 11650 12769 11706 12825
rect 11774 12769 11830 12825
rect 11898 12769 11954 12825
rect 12022 12769 12078 12825
rect 12146 12769 12202 12825
rect 12270 12769 12326 12825
rect 12394 12769 12450 12825
rect 12518 12769 12574 12825
rect 12642 12769 12698 12825
rect 12766 12769 12822 12825
rect 12890 12769 12946 12825
rect 13014 12769 13070 12825
rect -254 12645 -198 12701
rect -130 12645 -74 12701
rect -6 12645 50 12701
rect 118 12645 174 12701
rect 242 12645 298 12701
rect 366 12645 422 12701
rect 490 12645 546 12701
rect 614 12645 670 12701
rect 738 12645 794 12701
rect 862 12645 918 12701
rect 986 12645 1042 12701
rect 1110 12645 1166 12701
rect 1234 12645 1290 12701
rect 1358 12645 1414 12701
rect 1482 12645 1538 12701
rect 1606 12645 1662 12701
rect 1730 12645 1786 12701
rect 1854 12645 1910 12701
rect 1978 12645 2034 12701
rect 2102 12645 2158 12701
rect 2226 12645 2282 12701
rect 2350 12645 2406 12701
rect 2474 12645 2530 12701
rect 2598 12645 2654 12701
rect 2722 12645 2778 12701
rect 2846 12645 2902 12701
rect 2970 12645 3026 12701
rect 3094 12645 3150 12701
rect 3218 12645 3274 12701
rect 3342 12645 3398 12701
rect 3466 12645 3522 12701
rect 3590 12645 3646 12701
rect 3714 12645 3770 12701
rect 3838 12645 3894 12701
rect 3962 12645 4018 12701
rect 4086 12645 4142 12701
rect 4210 12645 4266 12701
rect 4334 12645 4390 12701
rect 4458 12645 4514 12701
rect 4582 12645 4638 12701
rect 4706 12645 4762 12701
rect 4830 12645 4886 12701
rect 4954 12645 5010 12701
rect 5078 12645 5134 12701
rect 5202 12645 5258 12701
rect 5326 12645 5382 12701
rect 5450 12645 5506 12701
rect 5574 12645 5630 12701
rect 5698 12645 5754 12701
rect 5822 12645 5878 12701
rect 5946 12645 6002 12701
rect 6070 12645 6126 12701
rect 6194 12645 6250 12701
rect 6318 12645 6374 12701
rect 6442 12645 6498 12701
rect 6566 12645 6622 12701
rect 6690 12645 6746 12701
rect 6814 12645 6870 12701
rect 6938 12645 6994 12701
rect 7062 12645 7118 12701
rect 7186 12645 7242 12701
rect 7310 12645 7366 12701
rect 7434 12645 7490 12701
rect 7558 12645 7614 12701
rect 7682 12645 7738 12701
rect 7806 12645 7862 12701
rect 7930 12645 7986 12701
rect 8054 12645 8110 12701
rect 8178 12645 8234 12701
rect 8302 12645 8358 12701
rect 8426 12645 8482 12701
rect 8550 12645 8606 12701
rect 8674 12645 8730 12701
rect 8798 12645 8854 12701
rect 8922 12645 8978 12701
rect 9046 12645 9102 12701
rect 9170 12645 9226 12701
rect 9294 12645 9350 12701
rect 9418 12645 9474 12701
rect 9542 12645 9598 12701
rect 9666 12645 9722 12701
rect 9790 12645 9846 12701
rect 9914 12645 9970 12701
rect 10038 12645 10094 12701
rect 10162 12645 10218 12701
rect 10286 12645 10342 12701
rect 10410 12645 10466 12701
rect 10534 12645 10590 12701
rect 10658 12645 10714 12701
rect 10782 12645 10838 12701
rect 10906 12645 10962 12701
rect 11030 12645 11086 12701
rect 11154 12645 11210 12701
rect 11278 12645 11334 12701
rect 11402 12645 11458 12701
rect 11526 12645 11582 12701
rect 11650 12645 11706 12701
rect 11774 12645 11830 12701
rect 11898 12645 11954 12701
rect 12022 12645 12078 12701
rect 12146 12645 12202 12701
rect 12270 12645 12326 12701
rect 12394 12645 12450 12701
rect 12518 12645 12574 12701
rect 12642 12645 12698 12701
rect 12766 12645 12822 12701
rect 12890 12645 12946 12701
rect 13014 12645 13070 12701
rect -254 12521 -198 12577
rect -130 12521 -74 12577
rect -6 12521 50 12577
rect 118 12521 174 12577
rect 242 12521 298 12577
rect 366 12521 422 12577
rect 490 12521 546 12577
rect 614 12521 670 12577
rect 738 12521 794 12577
rect 862 12521 918 12577
rect 986 12521 1042 12577
rect 1110 12521 1166 12577
rect 1234 12521 1290 12577
rect 1358 12521 1414 12577
rect 1482 12521 1538 12577
rect 1606 12521 1662 12577
rect 1730 12521 1786 12577
rect 1854 12521 1910 12577
rect 1978 12521 2034 12577
rect 2102 12521 2158 12577
rect 2226 12521 2282 12577
rect 2350 12521 2406 12577
rect 2474 12521 2530 12577
rect 2598 12521 2654 12577
rect 2722 12521 2778 12577
rect 2846 12521 2902 12577
rect 2970 12521 3026 12577
rect 3094 12521 3150 12577
rect 3218 12521 3274 12577
rect 3342 12521 3398 12577
rect 3466 12521 3522 12577
rect 3590 12521 3646 12577
rect 3714 12521 3770 12577
rect 3838 12521 3894 12577
rect 3962 12521 4018 12577
rect 4086 12521 4142 12577
rect 4210 12521 4266 12577
rect 4334 12521 4390 12577
rect 4458 12521 4514 12577
rect 4582 12521 4638 12577
rect 4706 12521 4762 12577
rect 4830 12521 4886 12577
rect 4954 12521 5010 12577
rect 5078 12521 5134 12577
rect 5202 12521 5258 12577
rect 5326 12521 5382 12577
rect 5450 12521 5506 12577
rect 5574 12521 5630 12577
rect 5698 12521 5754 12577
rect 5822 12521 5878 12577
rect 5946 12521 6002 12577
rect 6070 12521 6126 12577
rect 6194 12521 6250 12577
rect 6318 12521 6374 12577
rect 6442 12521 6498 12577
rect 6566 12521 6622 12577
rect 6690 12521 6746 12577
rect 6814 12521 6870 12577
rect 6938 12521 6994 12577
rect 7062 12521 7118 12577
rect 7186 12521 7242 12577
rect 7310 12521 7366 12577
rect 7434 12521 7490 12577
rect 7558 12521 7614 12577
rect 7682 12521 7738 12577
rect 7806 12521 7862 12577
rect 7930 12521 7986 12577
rect 8054 12521 8110 12577
rect 8178 12521 8234 12577
rect 8302 12521 8358 12577
rect 8426 12521 8482 12577
rect 8550 12521 8606 12577
rect 8674 12521 8730 12577
rect 8798 12521 8854 12577
rect 8922 12521 8978 12577
rect 9046 12521 9102 12577
rect 9170 12521 9226 12577
rect 9294 12521 9350 12577
rect 9418 12521 9474 12577
rect 9542 12521 9598 12577
rect 9666 12521 9722 12577
rect 9790 12521 9846 12577
rect 9914 12521 9970 12577
rect 10038 12521 10094 12577
rect 10162 12521 10218 12577
rect 10286 12521 10342 12577
rect 10410 12521 10466 12577
rect 10534 12521 10590 12577
rect 10658 12521 10714 12577
rect 10782 12521 10838 12577
rect 10906 12521 10962 12577
rect 11030 12521 11086 12577
rect 11154 12521 11210 12577
rect 11278 12521 11334 12577
rect 11402 12521 11458 12577
rect 11526 12521 11582 12577
rect 11650 12521 11706 12577
rect 11774 12521 11830 12577
rect 11898 12521 11954 12577
rect 12022 12521 12078 12577
rect 12146 12521 12202 12577
rect 12270 12521 12326 12577
rect 12394 12521 12450 12577
rect 12518 12521 12574 12577
rect 12642 12521 12698 12577
rect 12766 12521 12822 12577
rect 12890 12521 12946 12577
rect 13014 12521 13070 12577
rect -286 12302 -230 12358
rect -162 12302 -106 12358
rect -38 12302 18 12358
rect 86 12302 142 12358
rect 210 12302 266 12358
rect -286 12178 -230 12234
rect -162 12178 -106 12234
rect -38 12178 18 12234
rect 86 12178 142 12234
rect 210 12178 266 12234
rect -286 12054 -230 12110
rect -162 12054 -106 12110
rect -38 12054 18 12110
rect 86 12054 142 12110
rect 210 12054 266 12110
rect -286 11930 -230 11986
rect -162 11930 -106 11986
rect -38 11930 18 11986
rect 86 11930 142 11986
rect 210 11930 266 11986
rect -286 11806 -230 11862
rect -162 11806 -106 11862
rect -38 11806 18 11862
rect 86 11806 142 11862
rect 210 11806 266 11862
rect -286 11682 -230 11738
rect -162 11682 -106 11738
rect -38 11682 18 11738
rect 86 11682 142 11738
rect 210 11682 266 11738
rect -286 11558 -230 11614
rect -162 11558 -106 11614
rect -38 11558 18 11614
rect 86 11558 142 11614
rect 210 11558 266 11614
rect -286 11434 -230 11490
rect -162 11434 -106 11490
rect -38 11434 18 11490
rect 86 11434 142 11490
rect 210 11434 266 11490
rect -286 11310 -230 11366
rect -162 11310 -106 11366
rect -38 11310 18 11366
rect 86 11310 142 11366
rect 210 11310 266 11366
rect -286 11186 -230 11242
rect -162 11186 -106 11242
rect -38 11186 18 11242
rect 86 11186 142 11242
rect 210 11186 266 11242
rect -286 11062 -230 11118
rect -162 11062 -106 11118
rect -38 11062 18 11118
rect 86 11062 142 11118
rect 210 11062 266 11118
rect -286 10938 -230 10994
rect -162 10938 -106 10994
rect -38 10938 18 10994
rect 86 10938 142 10994
rect 210 10938 266 10994
rect -286 10814 -230 10870
rect -162 10814 -106 10870
rect -38 10814 18 10870
rect 86 10814 142 10870
rect 210 10814 266 10870
rect -286 10690 -230 10746
rect -162 10690 -106 10746
rect -38 10690 18 10746
rect 86 10690 142 10746
rect 210 10690 266 10746
rect -286 10566 -230 10622
rect -162 10566 -106 10622
rect -38 10566 18 10622
rect 86 10566 142 10622
rect 210 10566 266 10622
rect -286 10442 -230 10498
rect -162 10442 -106 10498
rect -38 10442 18 10498
rect 86 10442 142 10498
rect 210 10442 266 10498
rect -286 10318 -230 10374
rect -162 10318 -106 10374
rect -38 10318 18 10374
rect 86 10318 142 10374
rect 210 10318 266 10374
rect -286 10194 -230 10250
rect -162 10194 -106 10250
rect -38 10194 18 10250
rect 86 10194 142 10250
rect 210 10194 266 10250
rect -286 10070 -230 10126
rect -162 10070 -106 10126
rect -38 10070 18 10126
rect 86 10070 142 10126
rect 210 10070 266 10126
rect -286 9946 -230 10002
rect -162 9946 -106 10002
rect -38 9946 18 10002
rect 86 9946 142 10002
rect 210 9946 266 10002
rect -286 9822 -230 9878
rect -162 9822 -106 9878
rect -38 9822 18 9878
rect 86 9822 142 9878
rect 210 9822 266 9878
rect -286 9698 -230 9754
rect -162 9698 -106 9754
rect -38 9698 18 9754
rect 86 9698 142 9754
rect 210 9698 266 9754
rect -286 9574 -230 9630
rect -162 9574 -106 9630
rect -38 9574 18 9630
rect 86 9574 142 9630
rect 210 9574 266 9630
rect -286 9450 -230 9506
rect -162 9450 -106 9506
rect -38 9450 18 9506
rect 86 9450 142 9506
rect 210 9450 266 9506
rect -286 9326 -230 9382
rect -162 9326 -106 9382
rect -38 9326 18 9382
rect 86 9326 142 9382
rect 210 9326 266 9382
rect -286 9202 -230 9258
rect -162 9202 -106 9258
rect -38 9202 18 9258
rect 86 9202 142 9258
rect 210 9202 266 9258
rect -286 9078 -230 9134
rect -162 9078 -106 9134
rect -38 9078 18 9134
rect 86 9078 142 9134
rect 210 9078 266 9134
rect -286 8954 -230 9010
rect -162 8954 -106 9010
rect -38 8954 18 9010
rect 86 8954 142 9010
rect 210 8954 266 9010
rect -286 8830 -230 8886
rect -162 8830 -106 8886
rect -38 8830 18 8886
rect 86 8830 142 8886
rect 210 8830 266 8886
rect -286 8706 -230 8762
rect -162 8706 -106 8762
rect -38 8706 18 8762
rect 86 8706 142 8762
rect 210 8706 266 8762
rect -286 8582 -230 8638
rect -162 8582 -106 8638
rect -38 8582 18 8638
rect 86 8582 142 8638
rect 210 8582 266 8638
rect -286 8458 -230 8514
rect -162 8458 -106 8514
rect -38 8458 18 8514
rect 86 8458 142 8514
rect 210 8458 266 8514
rect -286 8334 -230 8390
rect -162 8334 -106 8390
rect -38 8334 18 8390
rect 86 8334 142 8390
rect 210 8334 266 8390
rect -286 8210 -230 8266
rect -162 8210 -106 8266
rect -38 8210 18 8266
rect 86 8210 142 8266
rect 210 8210 266 8266
rect -286 8086 -230 8142
rect -162 8086 -106 8142
rect -38 8086 18 8142
rect 86 8086 142 8142
rect 210 8086 266 8142
rect -286 7962 -230 8018
rect -162 7962 -106 8018
rect -38 7962 18 8018
rect 86 7962 142 8018
rect 210 7962 266 8018
rect -286 7838 -230 7894
rect -162 7838 -106 7894
rect -38 7838 18 7894
rect 86 7838 142 7894
rect 210 7838 266 7894
rect -286 7714 -230 7770
rect -162 7714 -106 7770
rect -38 7714 18 7770
rect 86 7714 142 7770
rect 210 7714 266 7770
rect -286 7590 -230 7646
rect -162 7590 -106 7646
rect -38 7590 18 7646
rect 86 7590 142 7646
rect 210 7590 266 7646
rect -286 7466 -230 7522
rect -162 7466 -106 7522
rect -38 7466 18 7522
rect 86 7466 142 7522
rect 210 7466 266 7522
rect -286 7342 -230 7398
rect -162 7342 -106 7398
rect -38 7342 18 7398
rect 86 7342 142 7398
rect 210 7342 266 7398
rect -286 7218 -230 7274
rect -162 7218 -106 7274
rect -38 7218 18 7274
rect 86 7218 142 7274
rect 210 7218 266 7274
rect -286 7094 -230 7150
rect -162 7094 -106 7150
rect -38 7094 18 7150
rect 86 7094 142 7150
rect 210 7094 266 7150
rect -286 6970 -230 7026
rect -162 6970 -106 7026
rect -38 6970 18 7026
rect 86 6970 142 7026
rect 210 6970 266 7026
rect -286 6846 -230 6902
rect -162 6846 -106 6902
rect -38 6846 18 6902
rect 86 6846 142 6902
rect 210 6846 266 6902
rect -286 6722 -230 6778
rect -162 6722 -106 6778
rect -38 6722 18 6778
rect 86 6722 142 6778
rect 210 6722 266 6778
rect -286 6598 -230 6654
rect -162 6598 -106 6654
rect -38 6598 18 6654
rect 86 6598 142 6654
rect 210 6598 266 6654
rect -286 6474 -230 6530
rect -162 6474 -106 6530
rect -38 6474 18 6530
rect 86 6474 142 6530
rect 210 6474 266 6530
rect -286 6350 -230 6406
rect -162 6350 -106 6406
rect -38 6350 18 6406
rect 86 6350 142 6406
rect 210 6350 266 6406
rect -286 6226 -230 6282
rect -162 6226 -106 6282
rect -38 6226 18 6282
rect 86 6226 142 6282
rect 210 6226 266 6282
rect -286 6102 -230 6158
rect -162 6102 -106 6158
rect -38 6102 18 6158
rect 86 6102 142 6158
rect 210 6102 266 6158
rect -286 5978 -230 6034
rect -162 5978 -106 6034
rect -38 5978 18 6034
rect 86 5978 142 6034
rect 210 5978 266 6034
rect -286 5854 -230 5910
rect -162 5854 -106 5910
rect -38 5854 18 5910
rect 86 5854 142 5910
rect 210 5854 266 5910
rect -286 5730 -230 5786
rect -162 5730 -106 5786
rect -38 5730 18 5786
rect 86 5730 142 5786
rect 210 5730 266 5786
rect -286 5606 -230 5662
rect -162 5606 -106 5662
rect -38 5606 18 5662
rect 86 5606 142 5662
rect 210 5606 266 5662
rect -286 5482 -230 5538
rect -162 5482 -106 5538
rect -38 5482 18 5538
rect 86 5482 142 5538
rect 210 5482 266 5538
rect -286 5358 -230 5414
rect -162 5358 -106 5414
rect -38 5358 18 5414
rect 86 5358 142 5414
rect 210 5358 266 5414
rect -286 5234 -230 5290
rect -162 5234 -106 5290
rect -38 5234 18 5290
rect 86 5234 142 5290
rect 210 5234 266 5290
rect -286 5110 -230 5166
rect -162 5110 -106 5166
rect -38 5110 18 5166
rect 86 5110 142 5166
rect 210 5110 266 5166
rect -286 4986 -230 5042
rect -162 4986 -106 5042
rect -38 4986 18 5042
rect 86 4986 142 5042
rect 210 4986 266 5042
rect -286 4862 -230 4918
rect -162 4862 -106 4918
rect -38 4862 18 4918
rect 86 4862 142 4918
rect 210 4862 266 4918
rect -286 4738 -230 4794
rect -162 4738 -106 4794
rect -38 4738 18 4794
rect 86 4738 142 4794
rect 210 4738 266 4794
rect -286 4614 -230 4670
rect -162 4614 -106 4670
rect -38 4614 18 4670
rect 86 4614 142 4670
rect 210 4614 266 4670
rect -286 4490 -230 4546
rect -162 4490 -106 4546
rect -38 4490 18 4546
rect 86 4490 142 4546
rect 210 4490 266 4546
rect -286 4366 -230 4422
rect -162 4366 -106 4422
rect -38 4366 18 4422
rect 86 4366 142 4422
rect 210 4366 266 4422
rect -286 4242 -230 4298
rect -162 4242 -106 4298
rect -38 4242 18 4298
rect 86 4242 142 4298
rect 210 4242 266 4298
rect -286 4118 -230 4174
rect -162 4118 -106 4174
rect -38 4118 18 4174
rect 86 4118 142 4174
rect 210 4118 266 4174
rect -286 3994 -230 4050
rect -162 3994 -106 4050
rect -38 3994 18 4050
rect 86 3994 142 4050
rect 210 3994 266 4050
rect -286 3870 -230 3926
rect -162 3870 -106 3926
rect -38 3870 18 3926
rect 86 3870 142 3926
rect 210 3870 266 3926
rect -286 3746 -230 3802
rect -162 3746 -106 3802
rect -38 3746 18 3802
rect 86 3746 142 3802
rect 210 3746 266 3802
rect -286 3622 -230 3678
rect -162 3622 -106 3678
rect -38 3622 18 3678
rect 86 3622 142 3678
rect 210 3622 266 3678
rect -286 3498 -230 3554
rect -162 3498 -106 3554
rect -38 3498 18 3554
rect 86 3498 142 3554
rect 210 3498 266 3554
rect -286 3374 -230 3430
rect -162 3374 -106 3430
rect -38 3374 18 3430
rect 86 3374 142 3430
rect 210 3374 266 3430
rect -286 3250 -230 3306
rect -162 3250 -106 3306
rect -38 3250 18 3306
rect 86 3250 142 3306
rect 210 3250 266 3306
rect -286 3126 -230 3182
rect -162 3126 -106 3182
rect -38 3126 18 3182
rect 86 3126 142 3182
rect 210 3126 266 3182
rect -286 3002 -230 3058
rect -162 3002 -106 3058
rect -38 3002 18 3058
rect 86 3002 142 3058
rect 210 3002 266 3058
rect -286 2878 -230 2934
rect -162 2878 -106 2934
rect -38 2878 18 2934
rect 86 2878 142 2934
rect 210 2878 266 2934
rect -286 2754 -230 2810
rect -162 2754 -106 2810
rect -38 2754 18 2810
rect 86 2754 142 2810
rect 210 2754 266 2810
rect -286 2630 -230 2686
rect -162 2630 -106 2686
rect -38 2630 18 2686
rect 86 2630 142 2686
rect 210 2630 266 2686
rect -286 2506 -230 2562
rect -162 2506 -106 2562
rect -38 2506 18 2562
rect 86 2506 142 2562
rect 210 2506 266 2562
rect -286 2382 -230 2438
rect -162 2382 -106 2438
rect -38 2382 18 2438
rect 86 2382 142 2438
rect 210 2382 266 2438
rect -286 2258 -230 2314
rect -162 2258 -106 2314
rect -38 2258 18 2314
rect 86 2258 142 2314
rect 210 2258 266 2314
rect -286 2134 -230 2190
rect -162 2134 -106 2190
rect -38 2134 18 2190
rect 86 2134 142 2190
rect 210 2134 266 2190
rect -286 2010 -230 2066
rect -162 2010 -106 2066
rect -38 2010 18 2066
rect 86 2010 142 2066
rect 210 2010 266 2066
rect -286 1886 -230 1942
rect -162 1886 -106 1942
rect -38 1886 18 1942
rect 86 1886 142 1942
rect 210 1886 266 1942
rect -286 1762 -230 1818
rect -162 1762 -106 1818
rect -38 1762 18 1818
rect 86 1762 142 1818
rect 210 1762 266 1818
rect -286 1638 -230 1694
rect -162 1638 -106 1694
rect -38 1638 18 1694
rect 86 1638 142 1694
rect 210 1638 266 1694
rect -286 1514 -230 1570
rect -162 1514 -106 1570
rect -38 1514 18 1570
rect 86 1514 142 1570
rect 210 1514 266 1570
rect -286 1390 -230 1446
rect -162 1390 -106 1446
rect -38 1390 18 1446
rect 86 1390 142 1446
rect 210 1390 266 1446
rect -286 1266 -230 1322
rect -162 1266 -106 1322
rect -38 1266 18 1322
rect 86 1266 142 1322
rect 210 1266 266 1322
rect -286 1142 -230 1198
rect -162 1142 -106 1198
rect -38 1142 18 1198
rect 86 1142 142 1198
rect 210 1142 266 1198
rect -286 1018 -230 1074
rect -162 1018 -106 1074
rect -38 1018 18 1074
rect 86 1018 142 1074
rect 210 1018 266 1074
rect -286 894 -230 950
rect -162 894 -106 950
rect -38 894 18 950
rect 86 894 142 950
rect 210 894 266 950
rect -286 770 -230 826
rect -162 770 -106 826
rect -38 770 18 826
rect 86 770 142 826
rect 210 770 266 826
rect -286 646 -230 702
rect -162 646 -106 702
rect -38 646 18 702
rect 86 646 142 702
rect 210 646 266 702
rect -286 522 -230 578
rect -162 522 -106 578
rect -38 522 18 578
rect 86 522 142 578
rect 210 522 266 578
rect 903 12254 959 12310
rect 1045 12254 1101 12310
rect 903 12112 959 12168
rect 1045 12112 1101 12168
rect 903 11970 959 12026
rect 1045 11970 1101 12026
rect 903 11828 959 11884
rect 1045 11828 1101 11884
rect 903 11686 959 11742
rect 1045 11686 1101 11742
rect 903 11544 959 11600
rect 1045 11544 1101 11600
rect 903 11402 959 11458
rect 1045 11402 1101 11458
rect 903 11260 959 11316
rect 1045 11260 1101 11316
rect 903 11118 959 11174
rect 1045 11118 1101 11174
rect 903 10976 959 11032
rect 1045 10976 1101 11032
rect 903 10834 959 10890
rect 1045 10834 1101 10890
rect 903 10692 959 10748
rect 1045 10692 1101 10748
rect 903 10550 959 10606
rect 1045 10550 1101 10606
rect 903 10408 959 10464
rect 1045 10408 1101 10464
rect 903 10266 959 10322
rect 1045 10266 1101 10322
rect 903 10124 959 10180
rect 1045 10124 1101 10180
rect 903 9982 959 10038
rect 1045 9982 1101 10038
rect 903 9840 959 9896
rect 1045 9840 1101 9896
rect 903 9698 959 9754
rect 1045 9698 1101 9754
rect 903 9556 959 9612
rect 1045 9556 1101 9612
rect 903 9414 959 9470
rect 1045 9414 1101 9470
rect 903 9272 959 9328
rect 1045 9272 1101 9328
rect 903 9130 959 9186
rect 1045 9130 1101 9186
rect 903 8988 959 9044
rect 1045 8988 1101 9044
rect 903 8846 959 8902
rect 1045 8846 1101 8902
rect 903 8704 959 8760
rect 1045 8704 1101 8760
rect 903 8562 959 8618
rect 1045 8562 1101 8618
rect 903 8420 959 8476
rect 1045 8420 1101 8476
rect 903 8278 959 8334
rect 1045 8278 1101 8334
rect 903 8136 959 8192
rect 1045 8136 1101 8192
rect 903 7994 959 8050
rect 1045 7994 1101 8050
rect 903 7852 959 7908
rect 1045 7852 1101 7908
rect 903 7710 959 7766
rect 1045 7710 1101 7766
rect 903 7568 959 7624
rect 1045 7568 1101 7624
rect 903 7426 959 7482
rect 1045 7426 1101 7482
rect 903 7284 959 7340
rect 1045 7284 1101 7340
rect 903 7142 959 7198
rect 1045 7142 1101 7198
rect 903 7000 959 7056
rect 1045 7000 1101 7056
rect 903 6858 959 6914
rect 1045 6858 1101 6914
rect 903 6716 959 6772
rect 1045 6716 1101 6772
rect 903 6574 959 6630
rect 1045 6574 1101 6630
rect 903 6432 959 6488
rect 1045 6432 1101 6488
rect 903 6290 959 6346
rect 1045 6290 1101 6346
rect 903 6148 959 6204
rect 1045 6148 1101 6204
rect 903 6006 959 6062
rect 1045 6006 1101 6062
rect 903 5864 959 5920
rect 1045 5864 1101 5920
rect 903 5722 959 5778
rect 1045 5722 1101 5778
rect 903 5580 959 5636
rect 1045 5580 1101 5636
rect 903 5438 959 5494
rect 1045 5438 1101 5494
rect 903 5296 959 5352
rect 1045 5296 1101 5352
rect 903 5154 959 5210
rect 1045 5154 1101 5210
rect 903 5012 959 5068
rect 1045 5012 1101 5068
rect 903 4870 959 4926
rect 1045 4870 1101 4926
rect 903 4728 959 4784
rect 1045 4728 1101 4784
rect 903 4586 959 4642
rect 1045 4586 1101 4642
rect 903 4444 959 4500
rect 1045 4444 1101 4500
rect 903 4302 959 4358
rect 1045 4302 1101 4358
rect 903 4160 959 4216
rect 1045 4160 1101 4216
rect 903 4018 959 4074
rect 1045 4018 1101 4074
rect 903 3876 959 3932
rect 1045 3876 1101 3932
rect 903 3734 959 3790
rect 1045 3734 1101 3790
rect 903 3592 959 3648
rect 1045 3592 1101 3648
rect 903 3450 959 3506
rect 1045 3450 1101 3506
rect 903 3308 959 3364
rect 1045 3308 1101 3364
rect 903 3166 959 3222
rect 1045 3166 1101 3222
rect 903 3024 959 3080
rect 1045 3024 1101 3080
rect 903 2882 959 2938
rect 1045 2882 1101 2938
rect 903 2740 959 2796
rect 1045 2740 1101 2796
rect 903 2598 959 2654
rect 1045 2598 1101 2654
rect 903 2456 959 2512
rect 1045 2456 1101 2512
rect 903 2314 959 2370
rect 1045 2314 1101 2370
rect 903 2172 959 2228
rect 1045 2172 1101 2228
rect 903 2030 959 2086
rect 1045 2030 1101 2086
rect 903 1888 959 1944
rect 1045 1888 1101 1944
rect 903 1746 959 1802
rect 1045 1746 1101 1802
rect 903 1604 959 1660
rect 1045 1604 1101 1660
rect 903 1462 959 1518
rect 1045 1462 1101 1518
rect 903 1320 959 1376
rect 1045 1320 1101 1376
rect 903 1178 959 1234
rect 1045 1178 1101 1234
rect 903 1036 959 1092
rect 1045 1036 1101 1092
rect 903 894 959 950
rect 1045 894 1101 950
rect 903 752 959 808
rect 1045 752 1101 808
rect 903 610 959 666
rect 1045 610 1101 666
rect 903 468 959 524
rect 1045 468 1101 524
rect 1444 12254 1500 12310
rect 1586 12254 1642 12310
rect 1444 12112 1500 12168
rect 1586 12112 1642 12168
rect 1444 11970 1500 12026
rect 1586 11970 1642 12026
rect 1444 11828 1500 11884
rect 1586 11828 1642 11884
rect 1444 11686 1500 11742
rect 1586 11686 1642 11742
rect 1444 11544 1500 11600
rect 1586 11544 1642 11600
rect 1444 11402 1500 11458
rect 1586 11402 1642 11458
rect 1444 11260 1500 11316
rect 1586 11260 1642 11316
rect 1444 11118 1500 11174
rect 1586 11118 1642 11174
rect 1444 10976 1500 11032
rect 1586 10976 1642 11032
rect 1444 10834 1500 10890
rect 1586 10834 1642 10890
rect 1444 10692 1500 10748
rect 1586 10692 1642 10748
rect 1444 10550 1500 10606
rect 1586 10550 1642 10606
rect 1444 10408 1500 10464
rect 1586 10408 1642 10464
rect 1444 10266 1500 10322
rect 1586 10266 1642 10322
rect 1444 10124 1500 10180
rect 1586 10124 1642 10180
rect 1444 9982 1500 10038
rect 1586 9982 1642 10038
rect 1444 9840 1500 9896
rect 1586 9840 1642 9896
rect 1444 9698 1500 9754
rect 1586 9698 1642 9754
rect 1444 9556 1500 9612
rect 1586 9556 1642 9612
rect 1444 9414 1500 9470
rect 1586 9414 1642 9470
rect 1444 9272 1500 9328
rect 1586 9272 1642 9328
rect 1444 9130 1500 9186
rect 1586 9130 1642 9186
rect 1444 8988 1500 9044
rect 1586 8988 1642 9044
rect 1444 8846 1500 8902
rect 1586 8846 1642 8902
rect 1444 8704 1500 8760
rect 1586 8704 1642 8760
rect 1444 8562 1500 8618
rect 1586 8562 1642 8618
rect 1444 8420 1500 8476
rect 1586 8420 1642 8476
rect 1444 8278 1500 8334
rect 1586 8278 1642 8334
rect 1444 8136 1500 8192
rect 1586 8136 1642 8192
rect 1444 7994 1500 8050
rect 1586 7994 1642 8050
rect 1444 7852 1500 7908
rect 1586 7852 1642 7908
rect 1444 7710 1500 7766
rect 1586 7710 1642 7766
rect 1444 7568 1500 7624
rect 1586 7568 1642 7624
rect 1444 7426 1500 7482
rect 1586 7426 1642 7482
rect 1444 7284 1500 7340
rect 1586 7284 1642 7340
rect 1444 7142 1500 7198
rect 1586 7142 1642 7198
rect 1444 7000 1500 7056
rect 1586 7000 1642 7056
rect 1444 6858 1500 6914
rect 1586 6858 1642 6914
rect 1444 6716 1500 6772
rect 1586 6716 1642 6772
rect 1444 6574 1500 6630
rect 1586 6574 1642 6630
rect 1444 6432 1500 6488
rect 1586 6432 1642 6488
rect 1444 6290 1500 6346
rect 1586 6290 1642 6346
rect 1444 6148 1500 6204
rect 1586 6148 1642 6204
rect 1444 6006 1500 6062
rect 1586 6006 1642 6062
rect 1444 5864 1500 5920
rect 1586 5864 1642 5920
rect 1444 5722 1500 5778
rect 1586 5722 1642 5778
rect 1444 5580 1500 5636
rect 1586 5580 1642 5636
rect 1444 5438 1500 5494
rect 1586 5438 1642 5494
rect 1444 5296 1500 5352
rect 1586 5296 1642 5352
rect 1444 5154 1500 5210
rect 1586 5154 1642 5210
rect 1444 5012 1500 5068
rect 1586 5012 1642 5068
rect 1444 4870 1500 4926
rect 1586 4870 1642 4926
rect 1444 4728 1500 4784
rect 1586 4728 1642 4784
rect 1444 4586 1500 4642
rect 1586 4586 1642 4642
rect 1444 4444 1500 4500
rect 1586 4444 1642 4500
rect 1444 4302 1500 4358
rect 1586 4302 1642 4358
rect 1444 4160 1500 4216
rect 1586 4160 1642 4216
rect 1444 4018 1500 4074
rect 1586 4018 1642 4074
rect 1444 3876 1500 3932
rect 1586 3876 1642 3932
rect 1444 3734 1500 3790
rect 1586 3734 1642 3790
rect 1444 3592 1500 3648
rect 1586 3592 1642 3648
rect 1444 3450 1500 3506
rect 1586 3450 1642 3506
rect 1444 3308 1500 3364
rect 1586 3308 1642 3364
rect 1444 3166 1500 3222
rect 1586 3166 1642 3222
rect 1444 3024 1500 3080
rect 1586 3024 1642 3080
rect 1444 2882 1500 2938
rect 1586 2882 1642 2938
rect 1444 2740 1500 2796
rect 1586 2740 1642 2796
rect 1444 2598 1500 2654
rect 1586 2598 1642 2654
rect 1444 2456 1500 2512
rect 1586 2456 1642 2512
rect 1444 2314 1500 2370
rect 1586 2314 1642 2370
rect 1444 2172 1500 2228
rect 1586 2172 1642 2228
rect 1444 2030 1500 2086
rect 1586 2030 1642 2086
rect 1444 1888 1500 1944
rect 1586 1888 1642 1944
rect 1444 1746 1500 1802
rect 1586 1746 1642 1802
rect 1444 1604 1500 1660
rect 1586 1604 1642 1660
rect 1444 1462 1500 1518
rect 1586 1462 1642 1518
rect 1444 1320 1500 1376
rect 1586 1320 1642 1376
rect 1444 1178 1500 1234
rect 1586 1178 1642 1234
rect 1444 1036 1500 1092
rect 1586 1036 1642 1092
rect 1444 894 1500 950
rect 1586 894 1642 950
rect 1444 752 1500 808
rect 1586 752 1642 808
rect 1444 610 1500 666
rect 1586 610 1642 666
rect 1444 468 1500 524
rect 1586 468 1642 524
rect 1984 12254 2040 12310
rect 2126 12254 2182 12310
rect 1984 12112 2040 12168
rect 2126 12112 2182 12168
rect 1984 11970 2040 12026
rect 2126 11970 2182 12026
rect 1984 11828 2040 11884
rect 2126 11828 2182 11884
rect 1984 11686 2040 11742
rect 2126 11686 2182 11742
rect 1984 11544 2040 11600
rect 2126 11544 2182 11600
rect 1984 11402 2040 11458
rect 2126 11402 2182 11458
rect 1984 11260 2040 11316
rect 2126 11260 2182 11316
rect 1984 11118 2040 11174
rect 2126 11118 2182 11174
rect 1984 10976 2040 11032
rect 2126 10976 2182 11032
rect 1984 10834 2040 10890
rect 2126 10834 2182 10890
rect 1984 10692 2040 10748
rect 2126 10692 2182 10748
rect 1984 10550 2040 10606
rect 2126 10550 2182 10606
rect 1984 10408 2040 10464
rect 2126 10408 2182 10464
rect 1984 10266 2040 10322
rect 2126 10266 2182 10322
rect 1984 10124 2040 10180
rect 2126 10124 2182 10180
rect 1984 9982 2040 10038
rect 2126 9982 2182 10038
rect 1984 9840 2040 9896
rect 2126 9840 2182 9896
rect 1984 9698 2040 9754
rect 2126 9698 2182 9754
rect 1984 9556 2040 9612
rect 2126 9556 2182 9612
rect 1984 9414 2040 9470
rect 2126 9414 2182 9470
rect 1984 9272 2040 9328
rect 2126 9272 2182 9328
rect 1984 9130 2040 9186
rect 2126 9130 2182 9186
rect 1984 8988 2040 9044
rect 2126 8988 2182 9044
rect 1984 8846 2040 8902
rect 2126 8846 2182 8902
rect 1984 8704 2040 8760
rect 2126 8704 2182 8760
rect 1984 8562 2040 8618
rect 2126 8562 2182 8618
rect 1984 8420 2040 8476
rect 2126 8420 2182 8476
rect 1984 8278 2040 8334
rect 2126 8278 2182 8334
rect 1984 8136 2040 8192
rect 2126 8136 2182 8192
rect 1984 7994 2040 8050
rect 2126 7994 2182 8050
rect 1984 7852 2040 7908
rect 2126 7852 2182 7908
rect 1984 7710 2040 7766
rect 2126 7710 2182 7766
rect 1984 7568 2040 7624
rect 2126 7568 2182 7624
rect 1984 7426 2040 7482
rect 2126 7426 2182 7482
rect 1984 7284 2040 7340
rect 2126 7284 2182 7340
rect 1984 7142 2040 7198
rect 2126 7142 2182 7198
rect 1984 7000 2040 7056
rect 2126 7000 2182 7056
rect 1984 6858 2040 6914
rect 2126 6858 2182 6914
rect 1984 6716 2040 6772
rect 2126 6716 2182 6772
rect 1984 6574 2040 6630
rect 2126 6574 2182 6630
rect 1984 6432 2040 6488
rect 2126 6432 2182 6488
rect 1984 6290 2040 6346
rect 2126 6290 2182 6346
rect 1984 6148 2040 6204
rect 2126 6148 2182 6204
rect 1984 6006 2040 6062
rect 2126 6006 2182 6062
rect 1984 5864 2040 5920
rect 2126 5864 2182 5920
rect 1984 5722 2040 5778
rect 2126 5722 2182 5778
rect 1984 5580 2040 5636
rect 2126 5580 2182 5636
rect 1984 5438 2040 5494
rect 2126 5438 2182 5494
rect 1984 5296 2040 5352
rect 2126 5296 2182 5352
rect 1984 5154 2040 5210
rect 2126 5154 2182 5210
rect 1984 5012 2040 5068
rect 2126 5012 2182 5068
rect 1984 4870 2040 4926
rect 2126 4870 2182 4926
rect 1984 4728 2040 4784
rect 2126 4728 2182 4784
rect 1984 4586 2040 4642
rect 2126 4586 2182 4642
rect 1984 4444 2040 4500
rect 2126 4444 2182 4500
rect 1984 4302 2040 4358
rect 2126 4302 2182 4358
rect 1984 4160 2040 4216
rect 2126 4160 2182 4216
rect 1984 4018 2040 4074
rect 2126 4018 2182 4074
rect 1984 3876 2040 3932
rect 2126 3876 2182 3932
rect 1984 3734 2040 3790
rect 2126 3734 2182 3790
rect 1984 3592 2040 3648
rect 2126 3592 2182 3648
rect 1984 3450 2040 3506
rect 2126 3450 2182 3506
rect 1984 3308 2040 3364
rect 2126 3308 2182 3364
rect 1984 3166 2040 3222
rect 2126 3166 2182 3222
rect 1984 3024 2040 3080
rect 2126 3024 2182 3080
rect 1984 2882 2040 2938
rect 2126 2882 2182 2938
rect 1984 2740 2040 2796
rect 2126 2740 2182 2796
rect 1984 2598 2040 2654
rect 2126 2598 2182 2654
rect 1984 2456 2040 2512
rect 2126 2456 2182 2512
rect 1984 2314 2040 2370
rect 2126 2314 2182 2370
rect 1984 2172 2040 2228
rect 2126 2172 2182 2228
rect 1984 2030 2040 2086
rect 2126 2030 2182 2086
rect 1984 1888 2040 1944
rect 2126 1888 2182 1944
rect 1984 1746 2040 1802
rect 2126 1746 2182 1802
rect 1984 1604 2040 1660
rect 2126 1604 2182 1660
rect 1984 1462 2040 1518
rect 2126 1462 2182 1518
rect 1984 1320 2040 1376
rect 2126 1320 2182 1376
rect 1984 1178 2040 1234
rect 2126 1178 2182 1234
rect 1984 1036 2040 1092
rect 2126 1036 2182 1092
rect 1984 894 2040 950
rect 2126 894 2182 950
rect 1984 752 2040 808
rect 2126 752 2182 808
rect 1984 610 2040 666
rect 2126 610 2182 666
rect 1984 468 2040 524
rect 2126 468 2182 524
rect 2521 12254 2577 12310
rect 2663 12254 2719 12310
rect 2521 12112 2577 12168
rect 2663 12112 2719 12168
rect 2521 11970 2577 12026
rect 2663 11970 2719 12026
rect 2521 11828 2577 11884
rect 2663 11828 2719 11884
rect 2521 11686 2577 11742
rect 2663 11686 2719 11742
rect 2521 11544 2577 11600
rect 2663 11544 2719 11600
rect 2521 11402 2577 11458
rect 2663 11402 2719 11458
rect 2521 11260 2577 11316
rect 2663 11260 2719 11316
rect 2521 11118 2577 11174
rect 2663 11118 2719 11174
rect 2521 10976 2577 11032
rect 2663 10976 2719 11032
rect 2521 10834 2577 10890
rect 2663 10834 2719 10890
rect 2521 10692 2577 10748
rect 2663 10692 2719 10748
rect 2521 10550 2577 10606
rect 2663 10550 2719 10606
rect 2521 10408 2577 10464
rect 2663 10408 2719 10464
rect 2521 10266 2577 10322
rect 2663 10266 2719 10322
rect 2521 10124 2577 10180
rect 2663 10124 2719 10180
rect 2521 9982 2577 10038
rect 2663 9982 2719 10038
rect 2521 9840 2577 9896
rect 2663 9840 2719 9896
rect 2521 9698 2577 9754
rect 2663 9698 2719 9754
rect 2521 9556 2577 9612
rect 2663 9556 2719 9612
rect 2521 9414 2577 9470
rect 2663 9414 2719 9470
rect 2521 9272 2577 9328
rect 2663 9272 2719 9328
rect 2521 9130 2577 9186
rect 2663 9130 2719 9186
rect 2521 8988 2577 9044
rect 2663 8988 2719 9044
rect 2521 8846 2577 8902
rect 2663 8846 2719 8902
rect 2521 8704 2577 8760
rect 2663 8704 2719 8760
rect 2521 8562 2577 8618
rect 2663 8562 2719 8618
rect 2521 8420 2577 8476
rect 2663 8420 2719 8476
rect 2521 8278 2577 8334
rect 2663 8278 2719 8334
rect 2521 8136 2577 8192
rect 2663 8136 2719 8192
rect 2521 7994 2577 8050
rect 2663 7994 2719 8050
rect 2521 7852 2577 7908
rect 2663 7852 2719 7908
rect 2521 7710 2577 7766
rect 2663 7710 2719 7766
rect 2521 7568 2577 7624
rect 2663 7568 2719 7624
rect 2521 7426 2577 7482
rect 2663 7426 2719 7482
rect 2521 7284 2577 7340
rect 2663 7284 2719 7340
rect 2521 7142 2577 7198
rect 2663 7142 2719 7198
rect 2521 7000 2577 7056
rect 2663 7000 2719 7056
rect 2521 6858 2577 6914
rect 2663 6858 2719 6914
rect 2521 6716 2577 6772
rect 2663 6716 2719 6772
rect 2521 6574 2577 6630
rect 2663 6574 2719 6630
rect 2521 6432 2577 6488
rect 2663 6432 2719 6488
rect 2521 6290 2577 6346
rect 2663 6290 2719 6346
rect 2521 6148 2577 6204
rect 2663 6148 2719 6204
rect 2521 6006 2577 6062
rect 2663 6006 2719 6062
rect 2521 5864 2577 5920
rect 2663 5864 2719 5920
rect 2521 5722 2577 5778
rect 2663 5722 2719 5778
rect 2521 5580 2577 5636
rect 2663 5580 2719 5636
rect 2521 5438 2577 5494
rect 2663 5438 2719 5494
rect 2521 5296 2577 5352
rect 2663 5296 2719 5352
rect 2521 5154 2577 5210
rect 2663 5154 2719 5210
rect 2521 5012 2577 5068
rect 2663 5012 2719 5068
rect 2521 4870 2577 4926
rect 2663 4870 2719 4926
rect 2521 4728 2577 4784
rect 2663 4728 2719 4784
rect 2521 4586 2577 4642
rect 2663 4586 2719 4642
rect 2521 4444 2577 4500
rect 2663 4444 2719 4500
rect 2521 4302 2577 4358
rect 2663 4302 2719 4358
rect 2521 4160 2577 4216
rect 2663 4160 2719 4216
rect 2521 4018 2577 4074
rect 2663 4018 2719 4074
rect 2521 3876 2577 3932
rect 2663 3876 2719 3932
rect 2521 3734 2577 3790
rect 2663 3734 2719 3790
rect 2521 3592 2577 3648
rect 2663 3592 2719 3648
rect 2521 3450 2577 3506
rect 2663 3450 2719 3506
rect 2521 3308 2577 3364
rect 2663 3308 2719 3364
rect 2521 3166 2577 3222
rect 2663 3166 2719 3222
rect 2521 3024 2577 3080
rect 2663 3024 2719 3080
rect 2521 2882 2577 2938
rect 2663 2882 2719 2938
rect 2521 2740 2577 2796
rect 2663 2740 2719 2796
rect 2521 2598 2577 2654
rect 2663 2598 2719 2654
rect 2521 2456 2577 2512
rect 2663 2456 2719 2512
rect 2521 2314 2577 2370
rect 2663 2314 2719 2370
rect 2521 2172 2577 2228
rect 2663 2172 2719 2228
rect 2521 2030 2577 2086
rect 2663 2030 2719 2086
rect 2521 1888 2577 1944
rect 2663 1888 2719 1944
rect 2521 1746 2577 1802
rect 2663 1746 2719 1802
rect 2521 1604 2577 1660
rect 2663 1604 2719 1660
rect 2521 1462 2577 1518
rect 2663 1462 2719 1518
rect 2521 1320 2577 1376
rect 2663 1320 2719 1376
rect 2521 1178 2577 1234
rect 2663 1178 2719 1234
rect 2521 1036 2577 1092
rect 2663 1036 2719 1092
rect 2521 894 2577 950
rect 2663 894 2719 950
rect 2521 752 2577 808
rect 2663 752 2719 808
rect 2521 610 2577 666
rect 2663 610 2719 666
rect 2521 468 2577 524
rect 2663 468 2719 524
rect 3058 12254 3114 12310
rect 3200 12254 3256 12310
rect 3058 12112 3114 12168
rect 3200 12112 3256 12168
rect 3058 11970 3114 12026
rect 3200 11970 3256 12026
rect 3058 11828 3114 11884
rect 3200 11828 3256 11884
rect 3058 11686 3114 11742
rect 3200 11686 3256 11742
rect 3058 11544 3114 11600
rect 3200 11544 3256 11600
rect 3058 11402 3114 11458
rect 3200 11402 3256 11458
rect 3058 11260 3114 11316
rect 3200 11260 3256 11316
rect 3058 11118 3114 11174
rect 3200 11118 3256 11174
rect 3058 10976 3114 11032
rect 3200 10976 3256 11032
rect 3058 10834 3114 10890
rect 3200 10834 3256 10890
rect 3058 10692 3114 10748
rect 3200 10692 3256 10748
rect 3058 10550 3114 10606
rect 3200 10550 3256 10606
rect 3058 10408 3114 10464
rect 3200 10408 3256 10464
rect 3058 10266 3114 10322
rect 3200 10266 3256 10322
rect 3058 10124 3114 10180
rect 3200 10124 3256 10180
rect 3058 9982 3114 10038
rect 3200 9982 3256 10038
rect 3058 9840 3114 9896
rect 3200 9840 3256 9896
rect 3058 9698 3114 9754
rect 3200 9698 3256 9754
rect 3058 9556 3114 9612
rect 3200 9556 3256 9612
rect 3058 9414 3114 9470
rect 3200 9414 3256 9470
rect 3058 9272 3114 9328
rect 3200 9272 3256 9328
rect 3058 9130 3114 9186
rect 3200 9130 3256 9186
rect 3058 8988 3114 9044
rect 3200 8988 3256 9044
rect 3058 8846 3114 8902
rect 3200 8846 3256 8902
rect 3058 8704 3114 8760
rect 3200 8704 3256 8760
rect 3058 8562 3114 8618
rect 3200 8562 3256 8618
rect 3058 8420 3114 8476
rect 3200 8420 3256 8476
rect 3058 8278 3114 8334
rect 3200 8278 3256 8334
rect 3058 8136 3114 8192
rect 3200 8136 3256 8192
rect 3058 7994 3114 8050
rect 3200 7994 3256 8050
rect 3058 7852 3114 7908
rect 3200 7852 3256 7908
rect 3058 7710 3114 7766
rect 3200 7710 3256 7766
rect 3058 7568 3114 7624
rect 3200 7568 3256 7624
rect 3058 7426 3114 7482
rect 3200 7426 3256 7482
rect 3058 7284 3114 7340
rect 3200 7284 3256 7340
rect 3058 7142 3114 7198
rect 3200 7142 3256 7198
rect 3058 7000 3114 7056
rect 3200 7000 3256 7056
rect 3058 6858 3114 6914
rect 3200 6858 3256 6914
rect 3058 6716 3114 6772
rect 3200 6716 3256 6772
rect 3058 6574 3114 6630
rect 3200 6574 3256 6630
rect 3058 6432 3114 6488
rect 3200 6432 3256 6488
rect 3058 6290 3114 6346
rect 3200 6290 3256 6346
rect 3058 6148 3114 6204
rect 3200 6148 3256 6204
rect 3058 6006 3114 6062
rect 3200 6006 3256 6062
rect 3058 5864 3114 5920
rect 3200 5864 3256 5920
rect 3058 5722 3114 5778
rect 3200 5722 3256 5778
rect 3058 5580 3114 5636
rect 3200 5580 3256 5636
rect 3058 5438 3114 5494
rect 3200 5438 3256 5494
rect 3058 5296 3114 5352
rect 3200 5296 3256 5352
rect 3058 5154 3114 5210
rect 3200 5154 3256 5210
rect 3058 5012 3114 5068
rect 3200 5012 3256 5068
rect 3058 4870 3114 4926
rect 3200 4870 3256 4926
rect 3058 4728 3114 4784
rect 3200 4728 3256 4784
rect 3058 4586 3114 4642
rect 3200 4586 3256 4642
rect 3058 4444 3114 4500
rect 3200 4444 3256 4500
rect 3058 4302 3114 4358
rect 3200 4302 3256 4358
rect 3058 4160 3114 4216
rect 3200 4160 3256 4216
rect 3058 4018 3114 4074
rect 3200 4018 3256 4074
rect 3058 3876 3114 3932
rect 3200 3876 3256 3932
rect 3058 3734 3114 3790
rect 3200 3734 3256 3790
rect 3058 3592 3114 3648
rect 3200 3592 3256 3648
rect 3058 3450 3114 3506
rect 3200 3450 3256 3506
rect 3058 3308 3114 3364
rect 3200 3308 3256 3364
rect 3058 3166 3114 3222
rect 3200 3166 3256 3222
rect 3058 3024 3114 3080
rect 3200 3024 3256 3080
rect 3058 2882 3114 2938
rect 3200 2882 3256 2938
rect 3058 2740 3114 2796
rect 3200 2740 3256 2796
rect 3058 2598 3114 2654
rect 3200 2598 3256 2654
rect 3058 2456 3114 2512
rect 3200 2456 3256 2512
rect 3058 2314 3114 2370
rect 3200 2314 3256 2370
rect 3058 2172 3114 2228
rect 3200 2172 3256 2228
rect 3058 2030 3114 2086
rect 3200 2030 3256 2086
rect 3058 1888 3114 1944
rect 3200 1888 3256 1944
rect 3058 1746 3114 1802
rect 3200 1746 3256 1802
rect 3058 1604 3114 1660
rect 3200 1604 3256 1660
rect 3058 1462 3114 1518
rect 3200 1462 3256 1518
rect 3058 1320 3114 1376
rect 3200 1320 3256 1376
rect 3058 1178 3114 1234
rect 3200 1178 3256 1234
rect 3058 1036 3114 1092
rect 3200 1036 3256 1092
rect 3058 894 3114 950
rect 3200 894 3256 950
rect 3058 752 3114 808
rect 3200 752 3256 808
rect 3058 610 3114 666
rect 3200 610 3256 666
rect 3058 468 3114 524
rect 3200 468 3256 524
rect 3602 12254 3658 12310
rect 3744 12254 3800 12310
rect 3602 12112 3658 12168
rect 3744 12112 3800 12168
rect 3602 11970 3658 12026
rect 3744 11970 3800 12026
rect 3602 11828 3658 11884
rect 3744 11828 3800 11884
rect 3602 11686 3658 11742
rect 3744 11686 3800 11742
rect 3602 11544 3658 11600
rect 3744 11544 3800 11600
rect 3602 11402 3658 11458
rect 3744 11402 3800 11458
rect 3602 11260 3658 11316
rect 3744 11260 3800 11316
rect 3602 11118 3658 11174
rect 3744 11118 3800 11174
rect 3602 10976 3658 11032
rect 3744 10976 3800 11032
rect 3602 10834 3658 10890
rect 3744 10834 3800 10890
rect 3602 10692 3658 10748
rect 3744 10692 3800 10748
rect 3602 10550 3658 10606
rect 3744 10550 3800 10606
rect 3602 10408 3658 10464
rect 3744 10408 3800 10464
rect 3602 10266 3658 10322
rect 3744 10266 3800 10322
rect 3602 10124 3658 10180
rect 3744 10124 3800 10180
rect 3602 9982 3658 10038
rect 3744 9982 3800 10038
rect 3602 9840 3658 9896
rect 3744 9840 3800 9896
rect 3602 9698 3658 9754
rect 3744 9698 3800 9754
rect 3602 9556 3658 9612
rect 3744 9556 3800 9612
rect 3602 9414 3658 9470
rect 3744 9414 3800 9470
rect 3602 9272 3658 9328
rect 3744 9272 3800 9328
rect 3602 9130 3658 9186
rect 3744 9130 3800 9186
rect 3602 8988 3658 9044
rect 3744 8988 3800 9044
rect 3602 8846 3658 8902
rect 3744 8846 3800 8902
rect 3602 8704 3658 8760
rect 3744 8704 3800 8760
rect 3602 8562 3658 8618
rect 3744 8562 3800 8618
rect 3602 8420 3658 8476
rect 3744 8420 3800 8476
rect 3602 8278 3658 8334
rect 3744 8278 3800 8334
rect 3602 8136 3658 8192
rect 3744 8136 3800 8192
rect 3602 7994 3658 8050
rect 3744 7994 3800 8050
rect 3602 7852 3658 7908
rect 3744 7852 3800 7908
rect 3602 7710 3658 7766
rect 3744 7710 3800 7766
rect 3602 7568 3658 7624
rect 3744 7568 3800 7624
rect 3602 7426 3658 7482
rect 3744 7426 3800 7482
rect 3602 7284 3658 7340
rect 3744 7284 3800 7340
rect 3602 7142 3658 7198
rect 3744 7142 3800 7198
rect 3602 7000 3658 7056
rect 3744 7000 3800 7056
rect 3602 6858 3658 6914
rect 3744 6858 3800 6914
rect 3602 6716 3658 6772
rect 3744 6716 3800 6772
rect 3602 6574 3658 6630
rect 3744 6574 3800 6630
rect 3602 6432 3658 6488
rect 3744 6432 3800 6488
rect 3602 6290 3658 6346
rect 3744 6290 3800 6346
rect 3602 6148 3658 6204
rect 3744 6148 3800 6204
rect 3602 6006 3658 6062
rect 3744 6006 3800 6062
rect 3602 5864 3658 5920
rect 3744 5864 3800 5920
rect 3602 5722 3658 5778
rect 3744 5722 3800 5778
rect 3602 5580 3658 5636
rect 3744 5580 3800 5636
rect 3602 5438 3658 5494
rect 3744 5438 3800 5494
rect 3602 5296 3658 5352
rect 3744 5296 3800 5352
rect 3602 5154 3658 5210
rect 3744 5154 3800 5210
rect 3602 5012 3658 5068
rect 3744 5012 3800 5068
rect 3602 4870 3658 4926
rect 3744 4870 3800 4926
rect 3602 4728 3658 4784
rect 3744 4728 3800 4784
rect 3602 4586 3658 4642
rect 3744 4586 3800 4642
rect 3602 4444 3658 4500
rect 3744 4444 3800 4500
rect 3602 4302 3658 4358
rect 3744 4302 3800 4358
rect 3602 4160 3658 4216
rect 3744 4160 3800 4216
rect 3602 4018 3658 4074
rect 3744 4018 3800 4074
rect 3602 3876 3658 3932
rect 3744 3876 3800 3932
rect 3602 3734 3658 3790
rect 3744 3734 3800 3790
rect 3602 3592 3658 3648
rect 3744 3592 3800 3648
rect 3602 3450 3658 3506
rect 3744 3450 3800 3506
rect 3602 3308 3658 3364
rect 3744 3308 3800 3364
rect 3602 3166 3658 3222
rect 3744 3166 3800 3222
rect 3602 3024 3658 3080
rect 3744 3024 3800 3080
rect 3602 2882 3658 2938
rect 3744 2882 3800 2938
rect 3602 2740 3658 2796
rect 3744 2740 3800 2796
rect 3602 2598 3658 2654
rect 3744 2598 3800 2654
rect 3602 2456 3658 2512
rect 3744 2456 3800 2512
rect 3602 2314 3658 2370
rect 3744 2314 3800 2370
rect 3602 2172 3658 2228
rect 3744 2172 3800 2228
rect 3602 2030 3658 2086
rect 3744 2030 3800 2086
rect 3602 1888 3658 1944
rect 3744 1888 3800 1944
rect 3602 1746 3658 1802
rect 3744 1746 3800 1802
rect 3602 1604 3658 1660
rect 3744 1604 3800 1660
rect 3602 1462 3658 1518
rect 3744 1462 3800 1518
rect 3602 1320 3658 1376
rect 3744 1320 3800 1376
rect 3602 1178 3658 1234
rect 3744 1178 3800 1234
rect 3602 1036 3658 1092
rect 3744 1036 3800 1092
rect 3602 894 3658 950
rect 3744 894 3800 950
rect 3602 752 3658 808
rect 3744 752 3800 808
rect 3602 610 3658 666
rect 3744 610 3800 666
rect 3602 468 3658 524
rect 3744 468 3800 524
rect 4138 12254 4194 12310
rect 4280 12254 4336 12310
rect 4138 12112 4194 12168
rect 4280 12112 4336 12168
rect 4138 11970 4194 12026
rect 4280 11970 4336 12026
rect 4138 11828 4194 11884
rect 4280 11828 4336 11884
rect 4138 11686 4194 11742
rect 4280 11686 4336 11742
rect 4138 11544 4194 11600
rect 4280 11544 4336 11600
rect 4138 11402 4194 11458
rect 4280 11402 4336 11458
rect 4138 11260 4194 11316
rect 4280 11260 4336 11316
rect 4138 11118 4194 11174
rect 4280 11118 4336 11174
rect 4138 10976 4194 11032
rect 4280 10976 4336 11032
rect 4138 10834 4194 10890
rect 4280 10834 4336 10890
rect 4138 10692 4194 10748
rect 4280 10692 4336 10748
rect 4138 10550 4194 10606
rect 4280 10550 4336 10606
rect 4138 10408 4194 10464
rect 4280 10408 4336 10464
rect 4138 10266 4194 10322
rect 4280 10266 4336 10322
rect 4138 10124 4194 10180
rect 4280 10124 4336 10180
rect 4138 9982 4194 10038
rect 4280 9982 4336 10038
rect 4138 9840 4194 9896
rect 4280 9840 4336 9896
rect 4138 9698 4194 9754
rect 4280 9698 4336 9754
rect 4138 9556 4194 9612
rect 4280 9556 4336 9612
rect 4138 9414 4194 9470
rect 4280 9414 4336 9470
rect 4138 9272 4194 9328
rect 4280 9272 4336 9328
rect 4138 9130 4194 9186
rect 4280 9130 4336 9186
rect 4138 8988 4194 9044
rect 4280 8988 4336 9044
rect 4138 8846 4194 8902
rect 4280 8846 4336 8902
rect 4138 8704 4194 8760
rect 4280 8704 4336 8760
rect 4138 8562 4194 8618
rect 4280 8562 4336 8618
rect 4138 8420 4194 8476
rect 4280 8420 4336 8476
rect 4138 8278 4194 8334
rect 4280 8278 4336 8334
rect 4138 8136 4194 8192
rect 4280 8136 4336 8192
rect 4138 7994 4194 8050
rect 4280 7994 4336 8050
rect 4138 7852 4194 7908
rect 4280 7852 4336 7908
rect 4138 7710 4194 7766
rect 4280 7710 4336 7766
rect 4138 7568 4194 7624
rect 4280 7568 4336 7624
rect 4138 7426 4194 7482
rect 4280 7426 4336 7482
rect 4138 7284 4194 7340
rect 4280 7284 4336 7340
rect 4138 7142 4194 7198
rect 4280 7142 4336 7198
rect 4138 7000 4194 7056
rect 4280 7000 4336 7056
rect 4138 6858 4194 6914
rect 4280 6858 4336 6914
rect 4138 6716 4194 6772
rect 4280 6716 4336 6772
rect 4138 6574 4194 6630
rect 4280 6574 4336 6630
rect 4138 6432 4194 6488
rect 4280 6432 4336 6488
rect 4138 6290 4194 6346
rect 4280 6290 4336 6346
rect 4138 6148 4194 6204
rect 4280 6148 4336 6204
rect 4138 6006 4194 6062
rect 4280 6006 4336 6062
rect 4138 5864 4194 5920
rect 4280 5864 4336 5920
rect 4138 5722 4194 5778
rect 4280 5722 4336 5778
rect 4138 5580 4194 5636
rect 4280 5580 4336 5636
rect 4138 5438 4194 5494
rect 4280 5438 4336 5494
rect 4138 5296 4194 5352
rect 4280 5296 4336 5352
rect 4138 5154 4194 5210
rect 4280 5154 4336 5210
rect 4138 5012 4194 5068
rect 4280 5012 4336 5068
rect 4138 4870 4194 4926
rect 4280 4870 4336 4926
rect 4138 4728 4194 4784
rect 4280 4728 4336 4784
rect 4138 4586 4194 4642
rect 4280 4586 4336 4642
rect 4138 4444 4194 4500
rect 4280 4444 4336 4500
rect 4138 4302 4194 4358
rect 4280 4302 4336 4358
rect 4138 4160 4194 4216
rect 4280 4160 4336 4216
rect 4138 4018 4194 4074
rect 4280 4018 4336 4074
rect 4138 3876 4194 3932
rect 4280 3876 4336 3932
rect 4138 3734 4194 3790
rect 4280 3734 4336 3790
rect 4138 3592 4194 3648
rect 4280 3592 4336 3648
rect 4138 3450 4194 3506
rect 4280 3450 4336 3506
rect 4138 3308 4194 3364
rect 4280 3308 4336 3364
rect 4138 3166 4194 3222
rect 4280 3166 4336 3222
rect 4138 3024 4194 3080
rect 4280 3024 4336 3080
rect 4138 2882 4194 2938
rect 4280 2882 4336 2938
rect 4138 2740 4194 2796
rect 4280 2740 4336 2796
rect 4138 2598 4194 2654
rect 4280 2598 4336 2654
rect 4138 2456 4194 2512
rect 4280 2456 4336 2512
rect 4138 2314 4194 2370
rect 4280 2314 4336 2370
rect 4138 2172 4194 2228
rect 4280 2172 4336 2228
rect 4138 2030 4194 2086
rect 4280 2030 4336 2086
rect 4138 1888 4194 1944
rect 4280 1888 4336 1944
rect 4138 1746 4194 1802
rect 4280 1746 4336 1802
rect 4138 1604 4194 1660
rect 4280 1604 4336 1660
rect 4138 1462 4194 1518
rect 4280 1462 4336 1518
rect 4138 1320 4194 1376
rect 4280 1320 4336 1376
rect 4138 1178 4194 1234
rect 4280 1178 4336 1234
rect 4138 1036 4194 1092
rect 4280 1036 4336 1092
rect 4138 894 4194 950
rect 4280 894 4336 950
rect 4138 752 4194 808
rect 4280 752 4336 808
rect 4138 610 4194 666
rect 4280 610 4336 666
rect 4138 468 4194 524
rect 4280 468 4336 524
rect 4678 12254 4734 12310
rect 4820 12254 4876 12310
rect 4678 12112 4734 12168
rect 4820 12112 4876 12168
rect 4678 11970 4734 12026
rect 4820 11970 4876 12026
rect 4678 11828 4734 11884
rect 4820 11828 4876 11884
rect 4678 11686 4734 11742
rect 4820 11686 4876 11742
rect 4678 11544 4734 11600
rect 4820 11544 4876 11600
rect 4678 11402 4734 11458
rect 4820 11402 4876 11458
rect 4678 11260 4734 11316
rect 4820 11260 4876 11316
rect 4678 11118 4734 11174
rect 4820 11118 4876 11174
rect 4678 10976 4734 11032
rect 4820 10976 4876 11032
rect 4678 10834 4734 10890
rect 4820 10834 4876 10890
rect 4678 10692 4734 10748
rect 4820 10692 4876 10748
rect 4678 10550 4734 10606
rect 4820 10550 4876 10606
rect 4678 10408 4734 10464
rect 4820 10408 4876 10464
rect 4678 10266 4734 10322
rect 4820 10266 4876 10322
rect 4678 10124 4734 10180
rect 4820 10124 4876 10180
rect 4678 9982 4734 10038
rect 4820 9982 4876 10038
rect 4678 9840 4734 9896
rect 4820 9840 4876 9896
rect 4678 9698 4734 9754
rect 4820 9698 4876 9754
rect 4678 9556 4734 9612
rect 4820 9556 4876 9612
rect 4678 9414 4734 9470
rect 4820 9414 4876 9470
rect 4678 9272 4734 9328
rect 4820 9272 4876 9328
rect 4678 9130 4734 9186
rect 4820 9130 4876 9186
rect 4678 8988 4734 9044
rect 4820 8988 4876 9044
rect 4678 8846 4734 8902
rect 4820 8846 4876 8902
rect 4678 8704 4734 8760
rect 4820 8704 4876 8760
rect 4678 8562 4734 8618
rect 4820 8562 4876 8618
rect 4678 8420 4734 8476
rect 4820 8420 4876 8476
rect 4678 8278 4734 8334
rect 4820 8278 4876 8334
rect 4678 8136 4734 8192
rect 4820 8136 4876 8192
rect 4678 7994 4734 8050
rect 4820 7994 4876 8050
rect 4678 7852 4734 7908
rect 4820 7852 4876 7908
rect 4678 7710 4734 7766
rect 4820 7710 4876 7766
rect 4678 7568 4734 7624
rect 4820 7568 4876 7624
rect 4678 7426 4734 7482
rect 4820 7426 4876 7482
rect 4678 7284 4734 7340
rect 4820 7284 4876 7340
rect 4678 7142 4734 7198
rect 4820 7142 4876 7198
rect 4678 7000 4734 7056
rect 4820 7000 4876 7056
rect 4678 6858 4734 6914
rect 4820 6858 4876 6914
rect 4678 6716 4734 6772
rect 4820 6716 4876 6772
rect 4678 6574 4734 6630
rect 4820 6574 4876 6630
rect 4678 6432 4734 6488
rect 4820 6432 4876 6488
rect 4678 6290 4734 6346
rect 4820 6290 4876 6346
rect 4678 6148 4734 6204
rect 4820 6148 4876 6204
rect 4678 6006 4734 6062
rect 4820 6006 4876 6062
rect 4678 5864 4734 5920
rect 4820 5864 4876 5920
rect 4678 5722 4734 5778
rect 4820 5722 4876 5778
rect 4678 5580 4734 5636
rect 4820 5580 4876 5636
rect 4678 5438 4734 5494
rect 4820 5438 4876 5494
rect 4678 5296 4734 5352
rect 4820 5296 4876 5352
rect 4678 5154 4734 5210
rect 4820 5154 4876 5210
rect 4678 5012 4734 5068
rect 4820 5012 4876 5068
rect 4678 4870 4734 4926
rect 4820 4870 4876 4926
rect 4678 4728 4734 4784
rect 4820 4728 4876 4784
rect 4678 4586 4734 4642
rect 4820 4586 4876 4642
rect 4678 4444 4734 4500
rect 4820 4444 4876 4500
rect 4678 4302 4734 4358
rect 4820 4302 4876 4358
rect 4678 4160 4734 4216
rect 4820 4160 4876 4216
rect 4678 4018 4734 4074
rect 4820 4018 4876 4074
rect 4678 3876 4734 3932
rect 4820 3876 4876 3932
rect 4678 3734 4734 3790
rect 4820 3734 4876 3790
rect 4678 3592 4734 3648
rect 4820 3592 4876 3648
rect 4678 3450 4734 3506
rect 4820 3450 4876 3506
rect 4678 3308 4734 3364
rect 4820 3308 4876 3364
rect 4678 3166 4734 3222
rect 4820 3166 4876 3222
rect 4678 3024 4734 3080
rect 4820 3024 4876 3080
rect 4678 2882 4734 2938
rect 4820 2882 4876 2938
rect 4678 2740 4734 2796
rect 4820 2740 4876 2796
rect 4678 2598 4734 2654
rect 4820 2598 4876 2654
rect 4678 2456 4734 2512
rect 4820 2456 4876 2512
rect 4678 2314 4734 2370
rect 4820 2314 4876 2370
rect 4678 2172 4734 2228
rect 4820 2172 4876 2228
rect 4678 2030 4734 2086
rect 4820 2030 4876 2086
rect 4678 1888 4734 1944
rect 4820 1888 4876 1944
rect 4678 1746 4734 1802
rect 4820 1746 4876 1802
rect 4678 1604 4734 1660
rect 4820 1604 4876 1660
rect 4678 1462 4734 1518
rect 4820 1462 4876 1518
rect 4678 1320 4734 1376
rect 4820 1320 4876 1376
rect 4678 1178 4734 1234
rect 4820 1178 4876 1234
rect 4678 1036 4734 1092
rect 4820 1036 4876 1092
rect 4678 894 4734 950
rect 4820 894 4876 950
rect 4678 752 4734 808
rect 4820 752 4876 808
rect 4678 610 4734 666
rect 4820 610 4876 666
rect 4678 468 4734 524
rect 4820 468 4876 524
rect 5215 12254 5271 12310
rect 5357 12254 5413 12310
rect 5215 12112 5271 12168
rect 5357 12112 5413 12168
rect 5215 11970 5271 12026
rect 5357 11970 5413 12026
rect 5215 11828 5271 11884
rect 5357 11828 5413 11884
rect 5215 11686 5271 11742
rect 5357 11686 5413 11742
rect 5215 11544 5271 11600
rect 5357 11544 5413 11600
rect 5215 11402 5271 11458
rect 5357 11402 5413 11458
rect 5215 11260 5271 11316
rect 5357 11260 5413 11316
rect 5215 11118 5271 11174
rect 5357 11118 5413 11174
rect 5215 10976 5271 11032
rect 5357 10976 5413 11032
rect 5215 10834 5271 10890
rect 5357 10834 5413 10890
rect 5215 10692 5271 10748
rect 5357 10692 5413 10748
rect 5215 10550 5271 10606
rect 5357 10550 5413 10606
rect 5215 10408 5271 10464
rect 5357 10408 5413 10464
rect 5215 10266 5271 10322
rect 5357 10266 5413 10322
rect 5215 10124 5271 10180
rect 5357 10124 5413 10180
rect 5215 9982 5271 10038
rect 5357 9982 5413 10038
rect 5215 9840 5271 9896
rect 5357 9840 5413 9896
rect 5215 9698 5271 9754
rect 5357 9698 5413 9754
rect 5215 9556 5271 9612
rect 5357 9556 5413 9612
rect 5215 9414 5271 9470
rect 5357 9414 5413 9470
rect 5215 9272 5271 9328
rect 5357 9272 5413 9328
rect 5215 9130 5271 9186
rect 5357 9130 5413 9186
rect 5215 8988 5271 9044
rect 5357 8988 5413 9044
rect 5215 8846 5271 8902
rect 5357 8846 5413 8902
rect 5215 8704 5271 8760
rect 5357 8704 5413 8760
rect 5215 8562 5271 8618
rect 5357 8562 5413 8618
rect 5215 8420 5271 8476
rect 5357 8420 5413 8476
rect 5215 8278 5271 8334
rect 5357 8278 5413 8334
rect 5215 8136 5271 8192
rect 5357 8136 5413 8192
rect 5215 7994 5271 8050
rect 5357 7994 5413 8050
rect 5215 7852 5271 7908
rect 5357 7852 5413 7908
rect 5215 7710 5271 7766
rect 5357 7710 5413 7766
rect 5215 7568 5271 7624
rect 5357 7568 5413 7624
rect 5215 7426 5271 7482
rect 5357 7426 5413 7482
rect 5215 7284 5271 7340
rect 5357 7284 5413 7340
rect 5215 7142 5271 7198
rect 5357 7142 5413 7198
rect 5215 7000 5271 7056
rect 5357 7000 5413 7056
rect 5215 6858 5271 6914
rect 5357 6858 5413 6914
rect 5215 6716 5271 6772
rect 5357 6716 5413 6772
rect 5215 6574 5271 6630
rect 5357 6574 5413 6630
rect 5215 6432 5271 6488
rect 5357 6432 5413 6488
rect 5215 6290 5271 6346
rect 5357 6290 5413 6346
rect 5215 6148 5271 6204
rect 5357 6148 5413 6204
rect 5215 6006 5271 6062
rect 5357 6006 5413 6062
rect 5215 5864 5271 5920
rect 5357 5864 5413 5920
rect 5215 5722 5271 5778
rect 5357 5722 5413 5778
rect 5215 5580 5271 5636
rect 5357 5580 5413 5636
rect 5215 5438 5271 5494
rect 5357 5438 5413 5494
rect 5215 5296 5271 5352
rect 5357 5296 5413 5352
rect 5215 5154 5271 5210
rect 5357 5154 5413 5210
rect 5215 5012 5271 5068
rect 5357 5012 5413 5068
rect 5215 4870 5271 4926
rect 5357 4870 5413 4926
rect 5215 4728 5271 4784
rect 5357 4728 5413 4784
rect 5215 4586 5271 4642
rect 5357 4586 5413 4642
rect 5215 4444 5271 4500
rect 5357 4444 5413 4500
rect 5215 4302 5271 4358
rect 5357 4302 5413 4358
rect 5215 4160 5271 4216
rect 5357 4160 5413 4216
rect 5215 4018 5271 4074
rect 5357 4018 5413 4074
rect 5215 3876 5271 3932
rect 5357 3876 5413 3932
rect 5215 3734 5271 3790
rect 5357 3734 5413 3790
rect 5215 3592 5271 3648
rect 5357 3592 5413 3648
rect 5215 3450 5271 3506
rect 5357 3450 5413 3506
rect 5215 3308 5271 3364
rect 5357 3308 5413 3364
rect 5215 3166 5271 3222
rect 5357 3166 5413 3222
rect 5215 3024 5271 3080
rect 5357 3024 5413 3080
rect 5215 2882 5271 2938
rect 5357 2882 5413 2938
rect 5215 2740 5271 2796
rect 5357 2740 5413 2796
rect 5215 2598 5271 2654
rect 5357 2598 5413 2654
rect 5215 2456 5271 2512
rect 5357 2456 5413 2512
rect 5215 2314 5271 2370
rect 5357 2314 5413 2370
rect 5215 2172 5271 2228
rect 5357 2172 5413 2228
rect 5215 2030 5271 2086
rect 5357 2030 5413 2086
rect 5215 1888 5271 1944
rect 5357 1888 5413 1944
rect 5215 1746 5271 1802
rect 5357 1746 5413 1802
rect 5215 1604 5271 1660
rect 5357 1604 5413 1660
rect 5215 1462 5271 1518
rect 5357 1462 5413 1518
rect 5215 1320 5271 1376
rect 5357 1320 5413 1376
rect 5215 1178 5271 1234
rect 5357 1178 5413 1234
rect 5215 1036 5271 1092
rect 5357 1036 5413 1092
rect 5215 894 5271 950
rect 5357 894 5413 950
rect 5215 752 5271 808
rect 5357 752 5413 808
rect 5215 610 5271 666
rect 5357 610 5413 666
rect 5215 468 5271 524
rect 5357 468 5413 524
rect 5760 12254 5816 12310
rect 5902 12254 5958 12310
rect 5760 12112 5816 12168
rect 5902 12112 5958 12168
rect 5760 11970 5816 12026
rect 5902 11970 5958 12026
rect 5760 11828 5816 11884
rect 5902 11828 5958 11884
rect 5760 11686 5816 11742
rect 5902 11686 5958 11742
rect 5760 11544 5816 11600
rect 5902 11544 5958 11600
rect 5760 11402 5816 11458
rect 5902 11402 5958 11458
rect 5760 11260 5816 11316
rect 5902 11260 5958 11316
rect 5760 11118 5816 11174
rect 5902 11118 5958 11174
rect 5760 10976 5816 11032
rect 5902 10976 5958 11032
rect 5760 10834 5816 10890
rect 5902 10834 5958 10890
rect 5760 10692 5816 10748
rect 5902 10692 5958 10748
rect 5760 10550 5816 10606
rect 5902 10550 5958 10606
rect 5760 10408 5816 10464
rect 5902 10408 5958 10464
rect 5760 10266 5816 10322
rect 5902 10266 5958 10322
rect 5760 10124 5816 10180
rect 5902 10124 5958 10180
rect 5760 9982 5816 10038
rect 5902 9982 5958 10038
rect 5760 9840 5816 9896
rect 5902 9840 5958 9896
rect 5760 9698 5816 9754
rect 5902 9698 5958 9754
rect 5760 9556 5816 9612
rect 5902 9556 5958 9612
rect 5760 9414 5816 9470
rect 5902 9414 5958 9470
rect 5760 9272 5816 9328
rect 5902 9272 5958 9328
rect 5760 9130 5816 9186
rect 5902 9130 5958 9186
rect 5760 8988 5816 9044
rect 5902 8988 5958 9044
rect 5760 8846 5816 8902
rect 5902 8846 5958 8902
rect 5760 8704 5816 8760
rect 5902 8704 5958 8760
rect 5760 8562 5816 8618
rect 5902 8562 5958 8618
rect 5760 8420 5816 8476
rect 5902 8420 5958 8476
rect 5760 8278 5816 8334
rect 5902 8278 5958 8334
rect 5760 8136 5816 8192
rect 5902 8136 5958 8192
rect 5760 7994 5816 8050
rect 5902 7994 5958 8050
rect 5760 7852 5816 7908
rect 5902 7852 5958 7908
rect 5760 7710 5816 7766
rect 5902 7710 5958 7766
rect 5760 7568 5816 7624
rect 5902 7568 5958 7624
rect 5760 7426 5816 7482
rect 5902 7426 5958 7482
rect 5760 7284 5816 7340
rect 5902 7284 5958 7340
rect 5760 7142 5816 7198
rect 5902 7142 5958 7198
rect 5760 7000 5816 7056
rect 5902 7000 5958 7056
rect 5760 6858 5816 6914
rect 5902 6858 5958 6914
rect 5760 6716 5816 6772
rect 5902 6716 5958 6772
rect 5760 6574 5816 6630
rect 5902 6574 5958 6630
rect 5760 6432 5816 6488
rect 5902 6432 5958 6488
rect 5760 6290 5816 6346
rect 5902 6290 5958 6346
rect 5760 6148 5816 6204
rect 5902 6148 5958 6204
rect 5760 6006 5816 6062
rect 5902 6006 5958 6062
rect 5760 5864 5816 5920
rect 5902 5864 5958 5920
rect 5760 5722 5816 5778
rect 5902 5722 5958 5778
rect 5760 5580 5816 5636
rect 5902 5580 5958 5636
rect 5760 5438 5816 5494
rect 5902 5438 5958 5494
rect 5760 5296 5816 5352
rect 5902 5296 5958 5352
rect 5760 5154 5816 5210
rect 5902 5154 5958 5210
rect 5760 5012 5816 5068
rect 5902 5012 5958 5068
rect 5760 4870 5816 4926
rect 5902 4870 5958 4926
rect 5760 4728 5816 4784
rect 5902 4728 5958 4784
rect 5760 4586 5816 4642
rect 5902 4586 5958 4642
rect 5760 4444 5816 4500
rect 5902 4444 5958 4500
rect 5760 4302 5816 4358
rect 5902 4302 5958 4358
rect 5760 4160 5816 4216
rect 5902 4160 5958 4216
rect 5760 4018 5816 4074
rect 5902 4018 5958 4074
rect 5760 3876 5816 3932
rect 5902 3876 5958 3932
rect 5760 3734 5816 3790
rect 5902 3734 5958 3790
rect 5760 3592 5816 3648
rect 5902 3592 5958 3648
rect 5760 3450 5816 3506
rect 5902 3450 5958 3506
rect 5760 3308 5816 3364
rect 5902 3308 5958 3364
rect 5760 3166 5816 3222
rect 5902 3166 5958 3222
rect 5760 3024 5816 3080
rect 5902 3024 5958 3080
rect 5760 2882 5816 2938
rect 5902 2882 5958 2938
rect 5760 2740 5816 2796
rect 5902 2740 5958 2796
rect 5760 2598 5816 2654
rect 5902 2598 5958 2654
rect 5760 2456 5816 2512
rect 5902 2456 5958 2512
rect 5760 2314 5816 2370
rect 5902 2314 5958 2370
rect 5760 2172 5816 2228
rect 5902 2172 5958 2228
rect 5760 2030 5816 2086
rect 5902 2030 5958 2086
rect 5760 1888 5816 1944
rect 5902 1888 5958 1944
rect 5760 1746 5816 1802
rect 5902 1746 5958 1802
rect 5760 1604 5816 1660
rect 5902 1604 5958 1660
rect 5760 1462 5816 1518
rect 5902 1462 5958 1518
rect 5760 1320 5816 1376
rect 5902 1320 5958 1376
rect 5760 1178 5816 1234
rect 5902 1178 5958 1234
rect 5760 1036 5816 1092
rect 5902 1036 5958 1092
rect 5760 894 5816 950
rect 5902 894 5958 950
rect 5760 752 5816 808
rect 5902 752 5958 808
rect 5760 610 5816 666
rect 5902 610 5958 666
rect 5760 468 5816 524
rect 5902 468 5958 524
rect 6300 12254 6356 12310
rect 6442 12254 6498 12310
rect 6300 12112 6356 12168
rect 6442 12112 6498 12168
rect 6300 11970 6356 12026
rect 6442 11970 6498 12026
rect 6300 11828 6356 11884
rect 6442 11828 6498 11884
rect 6300 11686 6356 11742
rect 6442 11686 6498 11742
rect 6300 11544 6356 11600
rect 6442 11544 6498 11600
rect 6300 11402 6356 11458
rect 6442 11402 6498 11458
rect 6300 11260 6356 11316
rect 6442 11260 6498 11316
rect 6300 11118 6356 11174
rect 6442 11118 6498 11174
rect 6300 10976 6356 11032
rect 6442 10976 6498 11032
rect 6300 10834 6356 10890
rect 6442 10834 6498 10890
rect 6300 10692 6356 10748
rect 6442 10692 6498 10748
rect 6300 10550 6356 10606
rect 6442 10550 6498 10606
rect 6300 10408 6356 10464
rect 6442 10408 6498 10464
rect 6300 10266 6356 10322
rect 6442 10266 6498 10322
rect 6300 10124 6356 10180
rect 6442 10124 6498 10180
rect 6300 9982 6356 10038
rect 6442 9982 6498 10038
rect 6300 9840 6356 9896
rect 6442 9840 6498 9896
rect 6300 9698 6356 9754
rect 6442 9698 6498 9754
rect 6300 9556 6356 9612
rect 6442 9556 6498 9612
rect 6300 9414 6356 9470
rect 6442 9414 6498 9470
rect 6300 9272 6356 9328
rect 6442 9272 6498 9328
rect 6300 9130 6356 9186
rect 6442 9130 6498 9186
rect 6300 8988 6356 9044
rect 6442 8988 6498 9044
rect 6300 8846 6356 8902
rect 6442 8846 6498 8902
rect 6300 8704 6356 8760
rect 6442 8704 6498 8760
rect 6300 8562 6356 8618
rect 6442 8562 6498 8618
rect 6300 8420 6356 8476
rect 6442 8420 6498 8476
rect 6300 8278 6356 8334
rect 6442 8278 6498 8334
rect 6300 8136 6356 8192
rect 6442 8136 6498 8192
rect 6300 7994 6356 8050
rect 6442 7994 6498 8050
rect 6300 7852 6356 7908
rect 6442 7852 6498 7908
rect 6300 7710 6356 7766
rect 6442 7710 6498 7766
rect 6300 7568 6356 7624
rect 6442 7568 6498 7624
rect 6300 7426 6356 7482
rect 6442 7426 6498 7482
rect 6300 7284 6356 7340
rect 6442 7284 6498 7340
rect 6300 7142 6356 7198
rect 6442 7142 6498 7198
rect 6300 7000 6356 7056
rect 6442 7000 6498 7056
rect 6300 6858 6356 6914
rect 6442 6858 6498 6914
rect 6300 6716 6356 6772
rect 6442 6716 6498 6772
rect 6300 6574 6356 6630
rect 6442 6574 6498 6630
rect 6300 6432 6356 6488
rect 6442 6432 6498 6488
rect 6300 6290 6356 6346
rect 6442 6290 6498 6346
rect 6300 6148 6356 6204
rect 6442 6148 6498 6204
rect 6300 6006 6356 6062
rect 6442 6006 6498 6062
rect 6300 5864 6356 5920
rect 6442 5864 6498 5920
rect 6300 5722 6356 5778
rect 6442 5722 6498 5778
rect 6300 5580 6356 5636
rect 6442 5580 6498 5636
rect 6300 5438 6356 5494
rect 6442 5438 6498 5494
rect 6300 5296 6356 5352
rect 6442 5296 6498 5352
rect 6300 5154 6356 5210
rect 6442 5154 6498 5210
rect 6300 5012 6356 5068
rect 6442 5012 6498 5068
rect 6300 4870 6356 4926
rect 6442 4870 6498 4926
rect 6300 4728 6356 4784
rect 6442 4728 6498 4784
rect 6300 4586 6356 4642
rect 6442 4586 6498 4642
rect 6300 4444 6356 4500
rect 6442 4444 6498 4500
rect 6300 4302 6356 4358
rect 6442 4302 6498 4358
rect 6300 4160 6356 4216
rect 6442 4160 6498 4216
rect 6300 4018 6356 4074
rect 6442 4018 6498 4074
rect 6300 3876 6356 3932
rect 6442 3876 6498 3932
rect 6300 3734 6356 3790
rect 6442 3734 6498 3790
rect 6300 3592 6356 3648
rect 6442 3592 6498 3648
rect 6300 3450 6356 3506
rect 6442 3450 6498 3506
rect 6300 3308 6356 3364
rect 6442 3308 6498 3364
rect 6300 3166 6356 3222
rect 6442 3166 6498 3222
rect 6300 3024 6356 3080
rect 6442 3024 6498 3080
rect 6300 2882 6356 2938
rect 6442 2882 6498 2938
rect 6300 2740 6356 2796
rect 6442 2740 6498 2796
rect 6300 2598 6356 2654
rect 6442 2598 6498 2654
rect 6300 2456 6356 2512
rect 6442 2456 6498 2512
rect 6300 2314 6356 2370
rect 6442 2314 6498 2370
rect 6300 2172 6356 2228
rect 6442 2172 6498 2228
rect 6300 2030 6356 2086
rect 6442 2030 6498 2086
rect 6300 1888 6356 1944
rect 6442 1888 6498 1944
rect 6300 1746 6356 1802
rect 6442 1746 6498 1802
rect 6300 1604 6356 1660
rect 6442 1604 6498 1660
rect 6300 1462 6356 1518
rect 6442 1462 6498 1518
rect 6300 1320 6356 1376
rect 6442 1320 6498 1376
rect 6300 1178 6356 1234
rect 6442 1178 6498 1234
rect 6300 1036 6356 1092
rect 6442 1036 6498 1092
rect 6300 894 6356 950
rect 6442 894 6498 950
rect 6300 752 6356 808
rect 6442 752 6498 808
rect 6300 610 6356 666
rect 6442 610 6498 666
rect 6300 468 6356 524
rect 6442 468 6498 524
rect 6845 12254 6901 12310
rect 6987 12254 7043 12310
rect 6845 12112 6901 12168
rect 6987 12112 7043 12168
rect 6845 11970 6901 12026
rect 6987 11970 7043 12026
rect 6845 11828 6901 11884
rect 6987 11828 7043 11884
rect 6845 11686 6901 11742
rect 6987 11686 7043 11742
rect 6845 11544 6901 11600
rect 6987 11544 7043 11600
rect 6845 11402 6901 11458
rect 6987 11402 7043 11458
rect 6845 11260 6901 11316
rect 6987 11260 7043 11316
rect 6845 11118 6901 11174
rect 6987 11118 7043 11174
rect 6845 10976 6901 11032
rect 6987 10976 7043 11032
rect 6845 10834 6901 10890
rect 6987 10834 7043 10890
rect 6845 10692 6901 10748
rect 6987 10692 7043 10748
rect 6845 10550 6901 10606
rect 6987 10550 7043 10606
rect 6845 10408 6901 10464
rect 6987 10408 7043 10464
rect 6845 10266 6901 10322
rect 6987 10266 7043 10322
rect 6845 10124 6901 10180
rect 6987 10124 7043 10180
rect 6845 9982 6901 10038
rect 6987 9982 7043 10038
rect 6845 9840 6901 9896
rect 6987 9840 7043 9896
rect 6845 9698 6901 9754
rect 6987 9698 7043 9754
rect 6845 9556 6901 9612
rect 6987 9556 7043 9612
rect 6845 9414 6901 9470
rect 6987 9414 7043 9470
rect 6845 9272 6901 9328
rect 6987 9272 7043 9328
rect 6845 9130 6901 9186
rect 6987 9130 7043 9186
rect 6845 8988 6901 9044
rect 6987 8988 7043 9044
rect 6845 8846 6901 8902
rect 6987 8846 7043 8902
rect 6845 8704 6901 8760
rect 6987 8704 7043 8760
rect 6845 8562 6901 8618
rect 6987 8562 7043 8618
rect 6845 8420 6901 8476
rect 6987 8420 7043 8476
rect 6845 8278 6901 8334
rect 6987 8278 7043 8334
rect 6845 8136 6901 8192
rect 6987 8136 7043 8192
rect 6845 7994 6901 8050
rect 6987 7994 7043 8050
rect 6845 7852 6901 7908
rect 6987 7852 7043 7908
rect 6845 7710 6901 7766
rect 6987 7710 7043 7766
rect 6845 7568 6901 7624
rect 6987 7568 7043 7624
rect 6845 7426 6901 7482
rect 6987 7426 7043 7482
rect 6845 7284 6901 7340
rect 6987 7284 7043 7340
rect 6845 7142 6901 7198
rect 6987 7142 7043 7198
rect 6845 7000 6901 7056
rect 6987 7000 7043 7056
rect 6845 6858 6901 6914
rect 6987 6858 7043 6914
rect 6845 6716 6901 6772
rect 6987 6716 7043 6772
rect 6845 6574 6901 6630
rect 6987 6574 7043 6630
rect 6845 6432 6901 6488
rect 6987 6432 7043 6488
rect 6845 6290 6901 6346
rect 6987 6290 7043 6346
rect 6845 6148 6901 6204
rect 6987 6148 7043 6204
rect 6845 6006 6901 6062
rect 6987 6006 7043 6062
rect 6845 5864 6901 5920
rect 6987 5864 7043 5920
rect 6845 5722 6901 5778
rect 6987 5722 7043 5778
rect 6845 5580 6901 5636
rect 6987 5580 7043 5636
rect 6845 5438 6901 5494
rect 6987 5438 7043 5494
rect 6845 5296 6901 5352
rect 6987 5296 7043 5352
rect 6845 5154 6901 5210
rect 6987 5154 7043 5210
rect 6845 5012 6901 5068
rect 6987 5012 7043 5068
rect 6845 4870 6901 4926
rect 6987 4870 7043 4926
rect 6845 4728 6901 4784
rect 6987 4728 7043 4784
rect 6845 4586 6901 4642
rect 6987 4586 7043 4642
rect 6845 4444 6901 4500
rect 6987 4444 7043 4500
rect 6845 4302 6901 4358
rect 6987 4302 7043 4358
rect 6845 4160 6901 4216
rect 6987 4160 7043 4216
rect 6845 4018 6901 4074
rect 6987 4018 7043 4074
rect 6845 3876 6901 3932
rect 6987 3876 7043 3932
rect 6845 3734 6901 3790
rect 6987 3734 7043 3790
rect 6845 3592 6901 3648
rect 6987 3592 7043 3648
rect 6845 3450 6901 3506
rect 6987 3450 7043 3506
rect 6845 3308 6901 3364
rect 6987 3308 7043 3364
rect 6845 3166 6901 3222
rect 6987 3166 7043 3222
rect 6845 3024 6901 3080
rect 6987 3024 7043 3080
rect 6845 2882 6901 2938
rect 6987 2882 7043 2938
rect 6845 2740 6901 2796
rect 6987 2740 7043 2796
rect 6845 2598 6901 2654
rect 6987 2598 7043 2654
rect 6845 2456 6901 2512
rect 6987 2456 7043 2512
rect 6845 2314 6901 2370
rect 6987 2314 7043 2370
rect 6845 2172 6901 2228
rect 6987 2172 7043 2228
rect 6845 2030 6901 2086
rect 6987 2030 7043 2086
rect 6845 1888 6901 1944
rect 6987 1888 7043 1944
rect 6845 1746 6901 1802
rect 6987 1746 7043 1802
rect 6845 1604 6901 1660
rect 6987 1604 7043 1660
rect 6845 1462 6901 1518
rect 6987 1462 7043 1518
rect 6845 1320 6901 1376
rect 6987 1320 7043 1376
rect 6845 1178 6901 1234
rect 6987 1178 7043 1234
rect 6845 1036 6901 1092
rect 6987 1036 7043 1092
rect 6845 894 6901 950
rect 6987 894 7043 950
rect 6845 752 6901 808
rect 6987 752 7043 808
rect 6845 610 6901 666
rect 6987 610 7043 666
rect 6845 468 6901 524
rect 6987 468 7043 524
rect 7382 12254 7438 12310
rect 7524 12254 7580 12310
rect 7382 12112 7438 12168
rect 7524 12112 7580 12168
rect 7382 11970 7438 12026
rect 7524 11970 7580 12026
rect 7382 11828 7438 11884
rect 7524 11828 7580 11884
rect 7382 11686 7438 11742
rect 7524 11686 7580 11742
rect 7382 11544 7438 11600
rect 7524 11544 7580 11600
rect 7382 11402 7438 11458
rect 7524 11402 7580 11458
rect 7382 11260 7438 11316
rect 7524 11260 7580 11316
rect 7382 11118 7438 11174
rect 7524 11118 7580 11174
rect 7382 10976 7438 11032
rect 7524 10976 7580 11032
rect 7382 10834 7438 10890
rect 7524 10834 7580 10890
rect 7382 10692 7438 10748
rect 7524 10692 7580 10748
rect 7382 10550 7438 10606
rect 7524 10550 7580 10606
rect 7382 10408 7438 10464
rect 7524 10408 7580 10464
rect 7382 10266 7438 10322
rect 7524 10266 7580 10322
rect 7382 10124 7438 10180
rect 7524 10124 7580 10180
rect 7382 9982 7438 10038
rect 7524 9982 7580 10038
rect 7382 9840 7438 9896
rect 7524 9840 7580 9896
rect 7382 9698 7438 9754
rect 7524 9698 7580 9754
rect 7382 9556 7438 9612
rect 7524 9556 7580 9612
rect 7382 9414 7438 9470
rect 7524 9414 7580 9470
rect 7382 9272 7438 9328
rect 7524 9272 7580 9328
rect 7382 9130 7438 9186
rect 7524 9130 7580 9186
rect 7382 8988 7438 9044
rect 7524 8988 7580 9044
rect 7382 8846 7438 8902
rect 7524 8846 7580 8902
rect 7382 8704 7438 8760
rect 7524 8704 7580 8760
rect 7382 8562 7438 8618
rect 7524 8562 7580 8618
rect 7382 8420 7438 8476
rect 7524 8420 7580 8476
rect 7382 8278 7438 8334
rect 7524 8278 7580 8334
rect 7382 8136 7438 8192
rect 7524 8136 7580 8192
rect 7382 7994 7438 8050
rect 7524 7994 7580 8050
rect 7382 7852 7438 7908
rect 7524 7852 7580 7908
rect 7382 7710 7438 7766
rect 7524 7710 7580 7766
rect 7382 7568 7438 7624
rect 7524 7568 7580 7624
rect 7382 7426 7438 7482
rect 7524 7426 7580 7482
rect 7382 7284 7438 7340
rect 7524 7284 7580 7340
rect 7382 7142 7438 7198
rect 7524 7142 7580 7198
rect 7382 7000 7438 7056
rect 7524 7000 7580 7056
rect 7382 6858 7438 6914
rect 7524 6858 7580 6914
rect 7382 6716 7438 6772
rect 7524 6716 7580 6772
rect 7382 6574 7438 6630
rect 7524 6574 7580 6630
rect 7382 6432 7438 6488
rect 7524 6432 7580 6488
rect 7382 6290 7438 6346
rect 7524 6290 7580 6346
rect 7382 6148 7438 6204
rect 7524 6148 7580 6204
rect 7382 6006 7438 6062
rect 7524 6006 7580 6062
rect 7382 5864 7438 5920
rect 7524 5864 7580 5920
rect 7382 5722 7438 5778
rect 7524 5722 7580 5778
rect 7382 5580 7438 5636
rect 7524 5580 7580 5636
rect 7382 5438 7438 5494
rect 7524 5438 7580 5494
rect 7382 5296 7438 5352
rect 7524 5296 7580 5352
rect 7382 5154 7438 5210
rect 7524 5154 7580 5210
rect 7382 5012 7438 5068
rect 7524 5012 7580 5068
rect 7382 4870 7438 4926
rect 7524 4870 7580 4926
rect 7382 4728 7438 4784
rect 7524 4728 7580 4784
rect 7382 4586 7438 4642
rect 7524 4586 7580 4642
rect 7382 4444 7438 4500
rect 7524 4444 7580 4500
rect 7382 4302 7438 4358
rect 7524 4302 7580 4358
rect 7382 4160 7438 4216
rect 7524 4160 7580 4216
rect 7382 4018 7438 4074
rect 7524 4018 7580 4074
rect 7382 3876 7438 3932
rect 7524 3876 7580 3932
rect 7382 3734 7438 3790
rect 7524 3734 7580 3790
rect 7382 3592 7438 3648
rect 7524 3592 7580 3648
rect 7382 3450 7438 3506
rect 7524 3450 7580 3506
rect 7382 3308 7438 3364
rect 7524 3308 7580 3364
rect 7382 3166 7438 3222
rect 7524 3166 7580 3222
rect 7382 3024 7438 3080
rect 7524 3024 7580 3080
rect 7382 2882 7438 2938
rect 7524 2882 7580 2938
rect 7382 2740 7438 2796
rect 7524 2740 7580 2796
rect 7382 2598 7438 2654
rect 7524 2598 7580 2654
rect 7382 2456 7438 2512
rect 7524 2456 7580 2512
rect 7382 2314 7438 2370
rect 7524 2314 7580 2370
rect 7382 2172 7438 2228
rect 7524 2172 7580 2228
rect 7382 2030 7438 2086
rect 7524 2030 7580 2086
rect 7382 1888 7438 1944
rect 7524 1888 7580 1944
rect 7382 1746 7438 1802
rect 7524 1746 7580 1802
rect 7382 1604 7438 1660
rect 7524 1604 7580 1660
rect 7382 1462 7438 1518
rect 7524 1462 7580 1518
rect 7382 1320 7438 1376
rect 7524 1320 7580 1376
rect 7382 1178 7438 1234
rect 7524 1178 7580 1234
rect 7382 1036 7438 1092
rect 7524 1036 7580 1092
rect 7382 894 7438 950
rect 7524 894 7580 950
rect 7382 752 7438 808
rect 7524 752 7580 808
rect 7382 610 7438 666
rect 7524 610 7580 666
rect 7382 468 7438 524
rect 7524 468 7580 524
rect 7919 12254 7975 12310
rect 8061 12254 8117 12310
rect 7919 12112 7975 12168
rect 8061 12112 8117 12168
rect 7919 11970 7975 12026
rect 8061 11970 8117 12026
rect 7919 11828 7975 11884
rect 8061 11828 8117 11884
rect 7919 11686 7975 11742
rect 8061 11686 8117 11742
rect 7919 11544 7975 11600
rect 8061 11544 8117 11600
rect 7919 11402 7975 11458
rect 8061 11402 8117 11458
rect 7919 11260 7975 11316
rect 8061 11260 8117 11316
rect 7919 11118 7975 11174
rect 8061 11118 8117 11174
rect 7919 10976 7975 11032
rect 8061 10976 8117 11032
rect 7919 10834 7975 10890
rect 8061 10834 8117 10890
rect 7919 10692 7975 10748
rect 8061 10692 8117 10748
rect 7919 10550 7975 10606
rect 8061 10550 8117 10606
rect 7919 10408 7975 10464
rect 8061 10408 8117 10464
rect 7919 10266 7975 10322
rect 8061 10266 8117 10322
rect 7919 10124 7975 10180
rect 8061 10124 8117 10180
rect 7919 9982 7975 10038
rect 8061 9982 8117 10038
rect 7919 9840 7975 9896
rect 8061 9840 8117 9896
rect 7919 9698 7975 9754
rect 8061 9698 8117 9754
rect 7919 9556 7975 9612
rect 8061 9556 8117 9612
rect 7919 9414 7975 9470
rect 8061 9414 8117 9470
rect 7919 9272 7975 9328
rect 8061 9272 8117 9328
rect 7919 9130 7975 9186
rect 8061 9130 8117 9186
rect 7919 8988 7975 9044
rect 8061 8988 8117 9044
rect 7919 8846 7975 8902
rect 8061 8846 8117 8902
rect 7919 8704 7975 8760
rect 8061 8704 8117 8760
rect 7919 8562 7975 8618
rect 8061 8562 8117 8618
rect 7919 8420 7975 8476
rect 8061 8420 8117 8476
rect 7919 8278 7975 8334
rect 8061 8278 8117 8334
rect 7919 8136 7975 8192
rect 8061 8136 8117 8192
rect 7919 7994 7975 8050
rect 8061 7994 8117 8050
rect 7919 7852 7975 7908
rect 8061 7852 8117 7908
rect 7919 7710 7975 7766
rect 8061 7710 8117 7766
rect 7919 7568 7975 7624
rect 8061 7568 8117 7624
rect 7919 7426 7975 7482
rect 8061 7426 8117 7482
rect 7919 7284 7975 7340
rect 8061 7284 8117 7340
rect 7919 7142 7975 7198
rect 8061 7142 8117 7198
rect 7919 7000 7975 7056
rect 8061 7000 8117 7056
rect 7919 6858 7975 6914
rect 8061 6858 8117 6914
rect 7919 6716 7975 6772
rect 8061 6716 8117 6772
rect 7919 6574 7975 6630
rect 8061 6574 8117 6630
rect 7919 6432 7975 6488
rect 8061 6432 8117 6488
rect 7919 6290 7975 6346
rect 8061 6290 8117 6346
rect 7919 6148 7975 6204
rect 8061 6148 8117 6204
rect 7919 6006 7975 6062
rect 8061 6006 8117 6062
rect 7919 5864 7975 5920
rect 8061 5864 8117 5920
rect 7919 5722 7975 5778
rect 8061 5722 8117 5778
rect 7919 5580 7975 5636
rect 8061 5580 8117 5636
rect 7919 5438 7975 5494
rect 8061 5438 8117 5494
rect 7919 5296 7975 5352
rect 8061 5296 8117 5352
rect 7919 5154 7975 5210
rect 8061 5154 8117 5210
rect 7919 5012 7975 5068
rect 8061 5012 8117 5068
rect 7919 4870 7975 4926
rect 8061 4870 8117 4926
rect 7919 4728 7975 4784
rect 8061 4728 8117 4784
rect 7919 4586 7975 4642
rect 8061 4586 8117 4642
rect 7919 4444 7975 4500
rect 8061 4444 8117 4500
rect 7919 4302 7975 4358
rect 8061 4302 8117 4358
rect 7919 4160 7975 4216
rect 8061 4160 8117 4216
rect 7919 4018 7975 4074
rect 8061 4018 8117 4074
rect 7919 3876 7975 3932
rect 8061 3876 8117 3932
rect 7919 3734 7975 3790
rect 8061 3734 8117 3790
rect 7919 3592 7975 3648
rect 8061 3592 8117 3648
rect 7919 3450 7975 3506
rect 8061 3450 8117 3506
rect 7919 3308 7975 3364
rect 8061 3308 8117 3364
rect 7919 3166 7975 3222
rect 8061 3166 8117 3222
rect 7919 3024 7975 3080
rect 8061 3024 8117 3080
rect 7919 2882 7975 2938
rect 8061 2882 8117 2938
rect 7919 2740 7975 2796
rect 8061 2740 8117 2796
rect 7919 2598 7975 2654
rect 8061 2598 8117 2654
rect 7919 2456 7975 2512
rect 8061 2456 8117 2512
rect 7919 2314 7975 2370
rect 8061 2314 8117 2370
rect 7919 2172 7975 2228
rect 8061 2172 8117 2228
rect 7919 2030 7975 2086
rect 8061 2030 8117 2086
rect 7919 1888 7975 1944
rect 8061 1888 8117 1944
rect 7919 1746 7975 1802
rect 8061 1746 8117 1802
rect 7919 1604 7975 1660
rect 8061 1604 8117 1660
rect 7919 1462 7975 1518
rect 8061 1462 8117 1518
rect 7919 1320 7975 1376
rect 8061 1320 8117 1376
rect 7919 1178 7975 1234
rect 8061 1178 8117 1234
rect 7919 1036 7975 1092
rect 8061 1036 8117 1092
rect 7919 894 7975 950
rect 8061 894 8117 950
rect 7919 752 7975 808
rect 8061 752 8117 808
rect 7919 610 7975 666
rect 8061 610 8117 666
rect 7919 468 7975 524
rect 8061 468 8117 524
rect 8462 12254 8518 12310
rect 8604 12254 8660 12310
rect 8462 12112 8518 12168
rect 8604 12112 8660 12168
rect 8462 11970 8518 12026
rect 8604 11970 8660 12026
rect 8462 11828 8518 11884
rect 8604 11828 8660 11884
rect 8462 11686 8518 11742
rect 8604 11686 8660 11742
rect 8462 11544 8518 11600
rect 8604 11544 8660 11600
rect 8462 11402 8518 11458
rect 8604 11402 8660 11458
rect 8462 11260 8518 11316
rect 8604 11260 8660 11316
rect 8462 11118 8518 11174
rect 8604 11118 8660 11174
rect 8462 10976 8518 11032
rect 8604 10976 8660 11032
rect 8462 10834 8518 10890
rect 8604 10834 8660 10890
rect 8462 10692 8518 10748
rect 8604 10692 8660 10748
rect 8462 10550 8518 10606
rect 8604 10550 8660 10606
rect 8462 10408 8518 10464
rect 8604 10408 8660 10464
rect 8462 10266 8518 10322
rect 8604 10266 8660 10322
rect 8462 10124 8518 10180
rect 8604 10124 8660 10180
rect 8462 9982 8518 10038
rect 8604 9982 8660 10038
rect 8462 9840 8518 9896
rect 8604 9840 8660 9896
rect 8462 9698 8518 9754
rect 8604 9698 8660 9754
rect 8462 9556 8518 9612
rect 8604 9556 8660 9612
rect 8462 9414 8518 9470
rect 8604 9414 8660 9470
rect 8462 9272 8518 9328
rect 8604 9272 8660 9328
rect 8462 9130 8518 9186
rect 8604 9130 8660 9186
rect 8462 8988 8518 9044
rect 8604 8988 8660 9044
rect 8462 8846 8518 8902
rect 8604 8846 8660 8902
rect 8462 8704 8518 8760
rect 8604 8704 8660 8760
rect 8462 8562 8518 8618
rect 8604 8562 8660 8618
rect 8462 8420 8518 8476
rect 8604 8420 8660 8476
rect 8462 8278 8518 8334
rect 8604 8278 8660 8334
rect 8462 8136 8518 8192
rect 8604 8136 8660 8192
rect 8462 7994 8518 8050
rect 8604 7994 8660 8050
rect 8462 7852 8518 7908
rect 8604 7852 8660 7908
rect 8462 7710 8518 7766
rect 8604 7710 8660 7766
rect 8462 7568 8518 7624
rect 8604 7568 8660 7624
rect 8462 7426 8518 7482
rect 8604 7426 8660 7482
rect 8462 7284 8518 7340
rect 8604 7284 8660 7340
rect 8462 7142 8518 7198
rect 8604 7142 8660 7198
rect 8462 7000 8518 7056
rect 8604 7000 8660 7056
rect 8462 6858 8518 6914
rect 8604 6858 8660 6914
rect 8462 6716 8518 6772
rect 8604 6716 8660 6772
rect 8462 6574 8518 6630
rect 8604 6574 8660 6630
rect 8462 6432 8518 6488
rect 8604 6432 8660 6488
rect 8462 6290 8518 6346
rect 8604 6290 8660 6346
rect 8462 6148 8518 6204
rect 8604 6148 8660 6204
rect 8462 6006 8518 6062
rect 8604 6006 8660 6062
rect 8462 5864 8518 5920
rect 8604 5864 8660 5920
rect 8462 5722 8518 5778
rect 8604 5722 8660 5778
rect 8462 5580 8518 5636
rect 8604 5580 8660 5636
rect 8462 5438 8518 5494
rect 8604 5438 8660 5494
rect 8462 5296 8518 5352
rect 8604 5296 8660 5352
rect 8462 5154 8518 5210
rect 8604 5154 8660 5210
rect 8462 5012 8518 5068
rect 8604 5012 8660 5068
rect 8462 4870 8518 4926
rect 8604 4870 8660 4926
rect 8462 4728 8518 4784
rect 8604 4728 8660 4784
rect 8462 4586 8518 4642
rect 8604 4586 8660 4642
rect 8462 4444 8518 4500
rect 8604 4444 8660 4500
rect 8462 4302 8518 4358
rect 8604 4302 8660 4358
rect 8462 4160 8518 4216
rect 8604 4160 8660 4216
rect 8462 4018 8518 4074
rect 8604 4018 8660 4074
rect 8462 3876 8518 3932
rect 8604 3876 8660 3932
rect 8462 3734 8518 3790
rect 8604 3734 8660 3790
rect 8462 3592 8518 3648
rect 8604 3592 8660 3648
rect 8462 3450 8518 3506
rect 8604 3450 8660 3506
rect 8462 3308 8518 3364
rect 8604 3308 8660 3364
rect 8462 3166 8518 3222
rect 8604 3166 8660 3222
rect 8462 3024 8518 3080
rect 8604 3024 8660 3080
rect 8462 2882 8518 2938
rect 8604 2882 8660 2938
rect 8462 2740 8518 2796
rect 8604 2740 8660 2796
rect 8462 2598 8518 2654
rect 8604 2598 8660 2654
rect 8462 2456 8518 2512
rect 8604 2456 8660 2512
rect 8462 2314 8518 2370
rect 8604 2314 8660 2370
rect 8462 2172 8518 2228
rect 8604 2172 8660 2228
rect 8462 2030 8518 2086
rect 8604 2030 8660 2086
rect 8462 1888 8518 1944
rect 8604 1888 8660 1944
rect 8462 1746 8518 1802
rect 8604 1746 8660 1802
rect 8462 1604 8518 1660
rect 8604 1604 8660 1660
rect 8462 1462 8518 1518
rect 8604 1462 8660 1518
rect 8462 1320 8518 1376
rect 8604 1320 8660 1376
rect 8462 1178 8518 1234
rect 8604 1178 8660 1234
rect 8462 1036 8518 1092
rect 8604 1036 8660 1092
rect 8462 894 8518 950
rect 8604 894 8660 950
rect 8462 752 8518 808
rect 8604 752 8660 808
rect 8462 610 8518 666
rect 8604 610 8660 666
rect 8462 468 8518 524
rect 8604 468 8660 524
rect 9004 12254 9060 12310
rect 9146 12254 9202 12310
rect 9004 12112 9060 12168
rect 9146 12112 9202 12168
rect 9004 11970 9060 12026
rect 9146 11970 9202 12026
rect 9004 11828 9060 11884
rect 9146 11828 9202 11884
rect 9004 11686 9060 11742
rect 9146 11686 9202 11742
rect 9004 11544 9060 11600
rect 9146 11544 9202 11600
rect 9004 11402 9060 11458
rect 9146 11402 9202 11458
rect 9004 11260 9060 11316
rect 9146 11260 9202 11316
rect 9004 11118 9060 11174
rect 9146 11118 9202 11174
rect 9004 10976 9060 11032
rect 9146 10976 9202 11032
rect 9004 10834 9060 10890
rect 9146 10834 9202 10890
rect 9004 10692 9060 10748
rect 9146 10692 9202 10748
rect 9004 10550 9060 10606
rect 9146 10550 9202 10606
rect 9004 10408 9060 10464
rect 9146 10408 9202 10464
rect 9004 10266 9060 10322
rect 9146 10266 9202 10322
rect 9004 10124 9060 10180
rect 9146 10124 9202 10180
rect 9004 9982 9060 10038
rect 9146 9982 9202 10038
rect 9004 9840 9060 9896
rect 9146 9840 9202 9896
rect 9004 9698 9060 9754
rect 9146 9698 9202 9754
rect 9004 9556 9060 9612
rect 9146 9556 9202 9612
rect 9004 9414 9060 9470
rect 9146 9414 9202 9470
rect 9004 9272 9060 9328
rect 9146 9272 9202 9328
rect 9004 9130 9060 9186
rect 9146 9130 9202 9186
rect 9004 8988 9060 9044
rect 9146 8988 9202 9044
rect 9004 8846 9060 8902
rect 9146 8846 9202 8902
rect 9004 8704 9060 8760
rect 9146 8704 9202 8760
rect 9004 8562 9060 8618
rect 9146 8562 9202 8618
rect 9004 8420 9060 8476
rect 9146 8420 9202 8476
rect 9004 8278 9060 8334
rect 9146 8278 9202 8334
rect 9004 8136 9060 8192
rect 9146 8136 9202 8192
rect 9004 7994 9060 8050
rect 9146 7994 9202 8050
rect 9004 7852 9060 7908
rect 9146 7852 9202 7908
rect 9004 7710 9060 7766
rect 9146 7710 9202 7766
rect 9004 7568 9060 7624
rect 9146 7568 9202 7624
rect 9004 7426 9060 7482
rect 9146 7426 9202 7482
rect 9004 7284 9060 7340
rect 9146 7284 9202 7340
rect 9004 7142 9060 7198
rect 9146 7142 9202 7198
rect 9004 7000 9060 7056
rect 9146 7000 9202 7056
rect 9004 6858 9060 6914
rect 9146 6858 9202 6914
rect 9004 6716 9060 6772
rect 9146 6716 9202 6772
rect 9004 6574 9060 6630
rect 9146 6574 9202 6630
rect 9004 6432 9060 6488
rect 9146 6432 9202 6488
rect 9004 6290 9060 6346
rect 9146 6290 9202 6346
rect 9004 6148 9060 6204
rect 9146 6148 9202 6204
rect 9004 6006 9060 6062
rect 9146 6006 9202 6062
rect 9004 5864 9060 5920
rect 9146 5864 9202 5920
rect 9004 5722 9060 5778
rect 9146 5722 9202 5778
rect 9004 5580 9060 5636
rect 9146 5580 9202 5636
rect 9004 5438 9060 5494
rect 9146 5438 9202 5494
rect 9004 5296 9060 5352
rect 9146 5296 9202 5352
rect 9004 5154 9060 5210
rect 9146 5154 9202 5210
rect 9004 5012 9060 5068
rect 9146 5012 9202 5068
rect 9004 4870 9060 4926
rect 9146 4870 9202 4926
rect 9004 4728 9060 4784
rect 9146 4728 9202 4784
rect 9004 4586 9060 4642
rect 9146 4586 9202 4642
rect 9004 4444 9060 4500
rect 9146 4444 9202 4500
rect 9004 4302 9060 4358
rect 9146 4302 9202 4358
rect 9004 4160 9060 4216
rect 9146 4160 9202 4216
rect 9004 4018 9060 4074
rect 9146 4018 9202 4074
rect 9004 3876 9060 3932
rect 9146 3876 9202 3932
rect 9004 3734 9060 3790
rect 9146 3734 9202 3790
rect 9004 3592 9060 3648
rect 9146 3592 9202 3648
rect 9004 3450 9060 3506
rect 9146 3450 9202 3506
rect 9004 3308 9060 3364
rect 9146 3308 9202 3364
rect 9004 3166 9060 3222
rect 9146 3166 9202 3222
rect 9004 3024 9060 3080
rect 9146 3024 9202 3080
rect 9004 2882 9060 2938
rect 9146 2882 9202 2938
rect 9004 2740 9060 2796
rect 9146 2740 9202 2796
rect 9004 2598 9060 2654
rect 9146 2598 9202 2654
rect 9004 2456 9060 2512
rect 9146 2456 9202 2512
rect 9004 2314 9060 2370
rect 9146 2314 9202 2370
rect 9004 2172 9060 2228
rect 9146 2172 9202 2228
rect 9004 2030 9060 2086
rect 9146 2030 9202 2086
rect 9004 1888 9060 1944
rect 9146 1888 9202 1944
rect 9004 1746 9060 1802
rect 9146 1746 9202 1802
rect 9004 1604 9060 1660
rect 9146 1604 9202 1660
rect 9004 1462 9060 1518
rect 9146 1462 9202 1518
rect 9004 1320 9060 1376
rect 9146 1320 9202 1376
rect 9004 1178 9060 1234
rect 9146 1178 9202 1234
rect 9004 1036 9060 1092
rect 9146 1036 9202 1092
rect 9004 894 9060 950
rect 9146 894 9202 950
rect 9004 752 9060 808
rect 9146 752 9202 808
rect 9004 610 9060 666
rect 9146 610 9202 666
rect 9004 468 9060 524
rect 9146 468 9202 524
rect 9547 12254 9603 12310
rect 9689 12254 9745 12310
rect 9547 12112 9603 12168
rect 9689 12112 9745 12168
rect 9547 11970 9603 12026
rect 9689 11970 9745 12026
rect 9547 11828 9603 11884
rect 9689 11828 9745 11884
rect 9547 11686 9603 11742
rect 9689 11686 9745 11742
rect 9547 11544 9603 11600
rect 9689 11544 9745 11600
rect 9547 11402 9603 11458
rect 9689 11402 9745 11458
rect 9547 11260 9603 11316
rect 9689 11260 9745 11316
rect 9547 11118 9603 11174
rect 9689 11118 9745 11174
rect 9547 10976 9603 11032
rect 9689 10976 9745 11032
rect 9547 10834 9603 10890
rect 9689 10834 9745 10890
rect 9547 10692 9603 10748
rect 9689 10692 9745 10748
rect 9547 10550 9603 10606
rect 9689 10550 9745 10606
rect 9547 10408 9603 10464
rect 9689 10408 9745 10464
rect 9547 10266 9603 10322
rect 9689 10266 9745 10322
rect 9547 10124 9603 10180
rect 9689 10124 9745 10180
rect 9547 9982 9603 10038
rect 9689 9982 9745 10038
rect 9547 9840 9603 9896
rect 9689 9840 9745 9896
rect 9547 9698 9603 9754
rect 9689 9698 9745 9754
rect 9547 9556 9603 9612
rect 9689 9556 9745 9612
rect 9547 9414 9603 9470
rect 9689 9414 9745 9470
rect 9547 9272 9603 9328
rect 9689 9272 9745 9328
rect 9547 9130 9603 9186
rect 9689 9130 9745 9186
rect 9547 8988 9603 9044
rect 9689 8988 9745 9044
rect 9547 8846 9603 8902
rect 9689 8846 9745 8902
rect 9547 8704 9603 8760
rect 9689 8704 9745 8760
rect 9547 8562 9603 8618
rect 9689 8562 9745 8618
rect 9547 8420 9603 8476
rect 9689 8420 9745 8476
rect 9547 8278 9603 8334
rect 9689 8278 9745 8334
rect 9547 8136 9603 8192
rect 9689 8136 9745 8192
rect 9547 7994 9603 8050
rect 9689 7994 9745 8050
rect 9547 7852 9603 7908
rect 9689 7852 9745 7908
rect 9547 7710 9603 7766
rect 9689 7710 9745 7766
rect 9547 7568 9603 7624
rect 9689 7568 9745 7624
rect 9547 7426 9603 7482
rect 9689 7426 9745 7482
rect 9547 7284 9603 7340
rect 9689 7284 9745 7340
rect 9547 7142 9603 7198
rect 9689 7142 9745 7198
rect 9547 7000 9603 7056
rect 9689 7000 9745 7056
rect 9547 6858 9603 6914
rect 9689 6858 9745 6914
rect 9547 6716 9603 6772
rect 9689 6716 9745 6772
rect 9547 6574 9603 6630
rect 9689 6574 9745 6630
rect 9547 6432 9603 6488
rect 9689 6432 9745 6488
rect 9547 6290 9603 6346
rect 9689 6290 9745 6346
rect 9547 6148 9603 6204
rect 9689 6148 9745 6204
rect 9547 6006 9603 6062
rect 9689 6006 9745 6062
rect 9547 5864 9603 5920
rect 9689 5864 9745 5920
rect 9547 5722 9603 5778
rect 9689 5722 9745 5778
rect 9547 5580 9603 5636
rect 9689 5580 9745 5636
rect 9547 5438 9603 5494
rect 9689 5438 9745 5494
rect 9547 5296 9603 5352
rect 9689 5296 9745 5352
rect 9547 5154 9603 5210
rect 9689 5154 9745 5210
rect 9547 5012 9603 5068
rect 9689 5012 9745 5068
rect 9547 4870 9603 4926
rect 9689 4870 9745 4926
rect 9547 4728 9603 4784
rect 9689 4728 9745 4784
rect 9547 4586 9603 4642
rect 9689 4586 9745 4642
rect 9547 4444 9603 4500
rect 9689 4444 9745 4500
rect 9547 4302 9603 4358
rect 9689 4302 9745 4358
rect 9547 4160 9603 4216
rect 9689 4160 9745 4216
rect 9547 4018 9603 4074
rect 9689 4018 9745 4074
rect 9547 3876 9603 3932
rect 9689 3876 9745 3932
rect 9547 3734 9603 3790
rect 9689 3734 9745 3790
rect 9547 3592 9603 3648
rect 9689 3592 9745 3648
rect 9547 3450 9603 3506
rect 9689 3450 9745 3506
rect 9547 3308 9603 3364
rect 9689 3308 9745 3364
rect 9547 3166 9603 3222
rect 9689 3166 9745 3222
rect 9547 3024 9603 3080
rect 9689 3024 9745 3080
rect 9547 2882 9603 2938
rect 9689 2882 9745 2938
rect 9547 2740 9603 2796
rect 9689 2740 9745 2796
rect 9547 2598 9603 2654
rect 9689 2598 9745 2654
rect 9547 2456 9603 2512
rect 9689 2456 9745 2512
rect 9547 2314 9603 2370
rect 9689 2314 9745 2370
rect 9547 2172 9603 2228
rect 9689 2172 9745 2228
rect 9547 2030 9603 2086
rect 9689 2030 9745 2086
rect 9547 1888 9603 1944
rect 9689 1888 9745 1944
rect 9547 1746 9603 1802
rect 9689 1746 9745 1802
rect 9547 1604 9603 1660
rect 9689 1604 9745 1660
rect 9547 1462 9603 1518
rect 9689 1462 9745 1518
rect 9547 1320 9603 1376
rect 9689 1320 9745 1376
rect 9547 1178 9603 1234
rect 9689 1178 9745 1234
rect 9547 1036 9603 1092
rect 9689 1036 9745 1092
rect 9547 894 9603 950
rect 9689 894 9745 950
rect 9547 752 9603 808
rect 9689 752 9745 808
rect 9547 610 9603 666
rect 9689 610 9745 666
rect 9547 468 9603 524
rect 9689 468 9745 524
rect 10081 12254 10137 12310
rect 10223 12254 10279 12310
rect 10081 12112 10137 12168
rect 10223 12112 10279 12168
rect 10081 11970 10137 12026
rect 10223 11970 10279 12026
rect 10081 11828 10137 11884
rect 10223 11828 10279 11884
rect 10081 11686 10137 11742
rect 10223 11686 10279 11742
rect 10081 11544 10137 11600
rect 10223 11544 10279 11600
rect 10081 11402 10137 11458
rect 10223 11402 10279 11458
rect 10081 11260 10137 11316
rect 10223 11260 10279 11316
rect 10081 11118 10137 11174
rect 10223 11118 10279 11174
rect 10081 10976 10137 11032
rect 10223 10976 10279 11032
rect 10081 10834 10137 10890
rect 10223 10834 10279 10890
rect 10081 10692 10137 10748
rect 10223 10692 10279 10748
rect 10081 10550 10137 10606
rect 10223 10550 10279 10606
rect 10081 10408 10137 10464
rect 10223 10408 10279 10464
rect 10081 10266 10137 10322
rect 10223 10266 10279 10322
rect 10081 10124 10137 10180
rect 10223 10124 10279 10180
rect 10081 9982 10137 10038
rect 10223 9982 10279 10038
rect 10081 9840 10137 9896
rect 10223 9840 10279 9896
rect 10081 9698 10137 9754
rect 10223 9698 10279 9754
rect 10081 9556 10137 9612
rect 10223 9556 10279 9612
rect 10081 9414 10137 9470
rect 10223 9414 10279 9470
rect 10081 9272 10137 9328
rect 10223 9272 10279 9328
rect 10081 9130 10137 9186
rect 10223 9130 10279 9186
rect 10081 8988 10137 9044
rect 10223 8988 10279 9044
rect 10081 8846 10137 8902
rect 10223 8846 10279 8902
rect 10081 8704 10137 8760
rect 10223 8704 10279 8760
rect 10081 8562 10137 8618
rect 10223 8562 10279 8618
rect 10081 8420 10137 8476
rect 10223 8420 10279 8476
rect 10081 8278 10137 8334
rect 10223 8278 10279 8334
rect 10081 8136 10137 8192
rect 10223 8136 10279 8192
rect 10081 7994 10137 8050
rect 10223 7994 10279 8050
rect 10081 7852 10137 7908
rect 10223 7852 10279 7908
rect 10081 7710 10137 7766
rect 10223 7710 10279 7766
rect 10081 7568 10137 7624
rect 10223 7568 10279 7624
rect 10081 7426 10137 7482
rect 10223 7426 10279 7482
rect 10081 7284 10137 7340
rect 10223 7284 10279 7340
rect 10081 7142 10137 7198
rect 10223 7142 10279 7198
rect 10081 7000 10137 7056
rect 10223 7000 10279 7056
rect 10081 6858 10137 6914
rect 10223 6858 10279 6914
rect 10081 6716 10137 6772
rect 10223 6716 10279 6772
rect 10081 6574 10137 6630
rect 10223 6574 10279 6630
rect 10081 6432 10137 6488
rect 10223 6432 10279 6488
rect 10081 6290 10137 6346
rect 10223 6290 10279 6346
rect 10081 6148 10137 6204
rect 10223 6148 10279 6204
rect 10081 6006 10137 6062
rect 10223 6006 10279 6062
rect 10081 5864 10137 5920
rect 10223 5864 10279 5920
rect 10081 5722 10137 5778
rect 10223 5722 10279 5778
rect 10081 5580 10137 5636
rect 10223 5580 10279 5636
rect 10081 5438 10137 5494
rect 10223 5438 10279 5494
rect 10081 5296 10137 5352
rect 10223 5296 10279 5352
rect 10081 5154 10137 5210
rect 10223 5154 10279 5210
rect 10081 5012 10137 5068
rect 10223 5012 10279 5068
rect 10081 4870 10137 4926
rect 10223 4870 10279 4926
rect 10081 4728 10137 4784
rect 10223 4728 10279 4784
rect 10081 4586 10137 4642
rect 10223 4586 10279 4642
rect 10081 4444 10137 4500
rect 10223 4444 10279 4500
rect 10081 4302 10137 4358
rect 10223 4302 10279 4358
rect 10081 4160 10137 4216
rect 10223 4160 10279 4216
rect 10081 4018 10137 4074
rect 10223 4018 10279 4074
rect 10081 3876 10137 3932
rect 10223 3876 10279 3932
rect 10081 3734 10137 3790
rect 10223 3734 10279 3790
rect 10081 3592 10137 3648
rect 10223 3592 10279 3648
rect 10081 3450 10137 3506
rect 10223 3450 10279 3506
rect 10081 3308 10137 3364
rect 10223 3308 10279 3364
rect 10081 3166 10137 3222
rect 10223 3166 10279 3222
rect 10081 3024 10137 3080
rect 10223 3024 10279 3080
rect 10081 2882 10137 2938
rect 10223 2882 10279 2938
rect 10081 2740 10137 2796
rect 10223 2740 10279 2796
rect 10081 2598 10137 2654
rect 10223 2598 10279 2654
rect 10081 2456 10137 2512
rect 10223 2456 10279 2512
rect 10081 2314 10137 2370
rect 10223 2314 10279 2370
rect 10081 2172 10137 2228
rect 10223 2172 10279 2228
rect 10081 2030 10137 2086
rect 10223 2030 10279 2086
rect 10081 1888 10137 1944
rect 10223 1888 10279 1944
rect 10081 1746 10137 1802
rect 10223 1746 10279 1802
rect 10081 1604 10137 1660
rect 10223 1604 10279 1660
rect 10081 1462 10137 1518
rect 10223 1462 10279 1518
rect 10081 1320 10137 1376
rect 10223 1320 10279 1376
rect 10081 1178 10137 1234
rect 10223 1178 10279 1234
rect 10081 1036 10137 1092
rect 10223 1036 10279 1092
rect 10081 894 10137 950
rect 10223 894 10279 950
rect 10081 752 10137 808
rect 10223 752 10279 808
rect 10081 610 10137 666
rect 10223 610 10279 666
rect 10081 468 10137 524
rect 10223 468 10279 524
rect 10622 12254 10678 12310
rect 10764 12254 10820 12310
rect 10622 12112 10678 12168
rect 10764 12112 10820 12168
rect 10622 11970 10678 12026
rect 10764 11970 10820 12026
rect 10622 11828 10678 11884
rect 10764 11828 10820 11884
rect 10622 11686 10678 11742
rect 10764 11686 10820 11742
rect 10622 11544 10678 11600
rect 10764 11544 10820 11600
rect 10622 11402 10678 11458
rect 10764 11402 10820 11458
rect 10622 11260 10678 11316
rect 10764 11260 10820 11316
rect 10622 11118 10678 11174
rect 10764 11118 10820 11174
rect 10622 10976 10678 11032
rect 10764 10976 10820 11032
rect 10622 10834 10678 10890
rect 10764 10834 10820 10890
rect 10622 10692 10678 10748
rect 10764 10692 10820 10748
rect 10622 10550 10678 10606
rect 10764 10550 10820 10606
rect 10622 10408 10678 10464
rect 10764 10408 10820 10464
rect 10622 10266 10678 10322
rect 10764 10266 10820 10322
rect 10622 10124 10678 10180
rect 10764 10124 10820 10180
rect 10622 9982 10678 10038
rect 10764 9982 10820 10038
rect 10622 9840 10678 9896
rect 10764 9840 10820 9896
rect 10622 9698 10678 9754
rect 10764 9698 10820 9754
rect 10622 9556 10678 9612
rect 10764 9556 10820 9612
rect 10622 9414 10678 9470
rect 10764 9414 10820 9470
rect 10622 9272 10678 9328
rect 10764 9272 10820 9328
rect 10622 9130 10678 9186
rect 10764 9130 10820 9186
rect 10622 8988 10678 9044
rect 10764 8988 10820 9044
rect 10622 8846 10678 8902
rect 10764 8846 10820 8902
rect 10622 8704 10678 8760
rect 10764 8704 10820 8760
rect 10622 8562 10678 8618
rect 10764 8562 10820 8618
rect 10622 8420 10678 8476
rect 10764 8420 10820 8476
rect 10622 8278 10678 8334
rect 10764 8278 10820 8334
rect 10622 8136 10678 8192
rect 10764 8136 10820 8192
rect 10622 7994 10678 8050
rect 10764 7994 10820 8050
rect 10622 7852 10678 7908
rect 10764 7852 10820 7908
rect 10622 7710 10678 7766
rect 10764 7710 10820 7766
rect 10622 7568 10678 7624
rect 10764 7568 10820 7624
rect 10622 7426 10678 7482
rect 10764 7426 10820 7482
rect 10622 7284 10678 7340
rect 10764 7284 10820 7340
rect 10622 7142 10678 7198
rect 10764 7142 10820 7198
rect 10622 7000 10678 7056
rect 10764 7000 10820 7056
rect 10622 6858 10678 6914
rect 10764 6858 10820 6914
rect 10622 6716 10678 6772
rect 10764 6716 10820 6772
rect 10622 6574 10678 6630
rect 10764 6574 10820 6630
rect 10622 6432 10678 6488
rect 10764 6432 10820 6488
rect 10622 6290 10678 6346
rect 10764 6290 10820 6346
rect 10622 6148 10678 6204
rect 10764 6148 10820 6204
rect 10622 6006 10678 6062
rect 10764 6006 10820 6062
rect 10622 5864 10678 5920
rect 10764 5864 10820 5920
rect 10622 5722 10678 5778
rect 10764 5722 10820 5778
rect 10622 5580 10678 5636
rect 10764 5580 10820 5636
rect 10622 5438 10678 5494
rect 10764 5438 10820 5494
rect 10622 5296 10678 5352
rect 10764 5296 10820 5352
rect 10622 5154 10678 5210
rect 10764 5154 10820 5210
rect 10622 5012 10678 5068
rect 10764 5012 10820 5068
rect 10622 4870 10678 4926
rect 10764 4870 10820 4926
rect 10622 4728 10678 4784
rect 10764 4728 10820 4784
rect 10622 4586 10678 4642
rect 10764 4586 10820 4642
rect 10622 4444 10678 4500
rect 10764 4444 10820 4500
rect 10622 4302 10678 4358
rect 10764 4302 10820 4358
rect 10622 4160 10678 4216
rect 10764 4160 10820 4216
rect 10622 4018 10678 4074
rect 10764 4018 10820 4074
rect 10622 3876 10678 3932
rect 10764 3876 10820 3932
rect 10622 3734 10678 3790
rect 10764 3734 10820 3790
rect 10622 3592 10678 3648
rect 10764 3592 10820 3648
rect 10622 3450 10678 3506
rect 10764 3450 10820 3506
rect 10622 3308 10678 3364
rect 10764 3308 10820 3364
rect 10622 3166 10678 3222
rect 10764 3166 10820 3222
rect 10622 3024 10678 3080
rect 10764 3024 10820 3080
rect 10622 2882 10678 2938
rect 10764 2882 10820 2938
rect 10622 2740 10678 2796
rect 10764 2740 10820 2796
rect 10622 2598 10678 2654
rect 10764 2598 10820 2654
rect 10622 2456 10678 2512
rect 10764 2456 10820 2512
rect 10622 2314 10678 2370
rect 10764 2314 10820 2370
rect 10622 2172 10678 2228
rect 10764 2172 10820 2228
rect 10622 2030 10678 2086
rect 10764 2030 10820 2086
rect 10622 1888 10678 1944
rect 10764 1888 10820 1944
rect 10622 1746 10678 1802
rect 10764 1746 10820 1802
rect 10622 1604 10678 1660
rect 10764 1604 10820 1660
rect 10622 1462 10678 1518
rect 10764 1462 10820 1518
rect 10622 1320 10678 1376
rect 10764 1320 10820 1376
rect 10622 1178 10678 1234
rect 10764 1178 10820 1234
rect 10622 1036 10678 1092
rect 10764 1036 10820 1092
rect 10622 894 10678 950
rect 10764 894 10820 950
rect 10622 752 10678 808
rect 10764 752 10820 808
rect 10622 610 10678 666
rect 10764 610 10820 666
rect 10622 468 10678 524
rect 10764 468 10820 524
rect 11162 12254 11218 12310
rect 11304 12254 11360 12310
rect 11162 12112 11218 12168
rect 11304 12112 11360 12168
rect 11162 11970 11218 12026
rect 11304 11970 11360 12026
rect 11162 11828 11218 11884
rect 11304 11828 11360 11884
rect 11162 11686 11218 11742
rect 11304 11686 11360 11742
rect 11162 11544 11218 11600
rect 11304 11544 11360 11600
rect 11162 11402 11218 11458
rect 11304 11402 11360 11458
rect 11162 11260 11218 11316
rect 11304 11260 11360 11316
rect 11162 11118 11218 11174
rect 11304 11118 11360 11174
rect 11162 10976 11218 11032
rect 11304 10976 11360 11032
rect 11162 10834 11218 10890
rect 11304 10834 11360 10890
rect 11162 10692 11218 10748
rect 11304 10692 11360 10748
rect 11162 10550 11218 10606
rect 11304 10550 11360 10606
rect 11162 10408 11218 10464
rect 11304 10408 11360 10464
rect 11162 10266 11218 10322
rect 11304 10266 11360 10322
rect 11162 10124 11218 10180
rect 11304 10124 11360 10180
rect 11162 9982 11218 10038
rect 11304 9982 11360 10038
rect 11162 9840 11218 9896
rect 11304 9840 11360 9896
rect 11162 9698 11218 9754
rect 11304 9698 11360 9754
rect 11162 9556 11218 9612
rect 11304 9556 11360 9612
rect 11162 9414 11218 9470
rect 11304 9414 11360 9470
rect 11162 9272 11218 9328
rect 11304 9272 11360 9328
rect 11162 9130 11218 9186
rect 11304 9130 11360 9186
rect 11162 8988 11218 9044
rect 11304 8988 11360 9044
rect 11162 8846 11218 8902
rect 11304 8846 11360 8902
rect 11162 8704 11218 8760
rect 11304 8704 11360 8760
rect 11162 8562 11218 8618
rect 11304 8562 11360 8618
rect 11162 8420 11218 8476
rect 11304 8420 11360 8476
rect 11162 8278 11218 8334
rect 11304 8278 11360 8334
rect 11162 8136 11218 8192
rect 11304 8136 11360 8192
rect 11162 7994 11218 8050
rect 11304 7994 11360 8050
rect 11162 7852 11218 7908
rect 11304 7852 11360 7908
rect 11162 7710 11218 7766
rect 11304 7710 11360 7766
rect 11162 7568 11218 7624
rect 11304 7568 11360 7624
rect 11162 7426 11218 7482
rect 11304 7426 11360 7482
rect 11162 7284 11218 7340
rect 11304 7284 11360 7340
rect 11162 7142 11218 7198
rect 11304 7142 11360 7198
rect 11162 7000 11218 7056
rect 11304 7000 11360 7056
rect 11162 6858 11218 6914
rect 11304 6858 11360 6914
rect 11162 6716 11218 6772
rect 11304 6716 11360 6772
rect 11162 6574 11218 6630
rect 11304 6574 11360 6630
rect 11162 6432 11218 6488
rect 11304 6432 11360 6488
rect 11162 6290 11218 6346
rect 11304 6290 11360 6346
rect 11162 6148 11218 6204
rect 11304 6148 11360 6204
rect 11162 6006 11218 6062
rect 11304 6006 11360 6062
rect 11162 5864 11218 5920
rect 11304 5864 11360 5920
rect 11162 5722 11218 5778
rect 11304 5722 11360 5778
rect 11162 5580 11218 5636
rect 11304 5580 11360 5636
rect 11162 5438 11218 5494
rect 11304 5438 11360 5494
rect 11162 5296 11218 5352
rect 11304 5296 11360 5352
rect 11162 5154 11218 5210
rect 11304 5154 11360 5210
rect 11162 5012 11218 5068
rect 11304 5012 11360 5068
rect 11162 4870 11218 4926
rect 11304 4870 11360 4926
rect 11162 4728 11218 4784
rect 11304 4728 11360 4784
rect 11162 4586 11218 4642
rect 11304 4586 11360 4642
rect 11162 4444 11218 4500
rect 11304 4444 11360 4500
rect 11162 4302 11218 4358
rect 11304 4302 11360 4358
rect 11162 4160 11218 4216
rect 11304 4160 11360 4216
rect 11162 4018 11218 4074
rect 11304 4018 11360 4074
rect 11162 3876 11218 3932
rect 11304 3876 11360 3932
rect 11162 3734 11218 3790
rect 11304 3734 11360 3790
rect 11162 3592 11218 3648
rect 11304 3592 11360 3648
rect 11162 3450 11218 3506
rect 11304 3450 11360 3506
rect 11162 3308 11218 3364
rect 11304 3308 11360 3364
rect 11162 3166 11218 3222
rect 11304 3166 11360 3222
rect 11162 3024 11218 3080
rect 11304 3024 11360 3080
rect 11162 2882 11218 2938
rect 11304 2882 11360 2938
rect 11162 2740 11218 2796
rect 11304 2740 11360 2796
rect 11162 2598 11218 2654
rect 11304 2598 11360 2654
rect 11162 2456 11218 2512
rect 11304 2456 11360 2512
rect 11162 2314 11218 2370
rect 11304 2314 11360 2370
rect 11162 2172 11218 2228
rect 11304 2172 11360 2228
rect 11162 2030 11218 2086
rect 11304 2030 11360 2086
rect 11162 1888 11218 1944
rect 11304 1888 11360 1944
rect 11162 1746 11218 1802
rect 11304 1746 11360 1802
rect 11162 1604 11218 1660
rect 11304 1604 11360 1660
rect 11162 1462 11218 1518
rect 11304 1462 11360 1518
rect 11162 1320 11218 1376
rect 11304 1320 11360 1376
rect 11162 1178 11218 1234
rect 11304 1178 11360 1234
rect 11162 1036 11218 1092
rect 11304 1036 11360 1092
rect 11162 894 11218 950
rect 11304 894 11360 950
rect 11162 752 11218 808
rect 11304 752 11360 808
rect 11162 610 11218 666
rect 11304 610 11360 666
rect 11162 468 11218 524
rect 11304 468 11360 524
rect 11702 12254 11758 12310
rect 11844 12254 11900 12310
rect 11702 12112 11758 12168
rect 11844 12112 11900 12168
rect 11702 11970 11758 12026
rect 11844 11970 11900 12026
rect 11702 11828 11758 11884
rect 11844 11828 11900 11884
rect 11702 11686 11758 11742
rect 11844 11686 11900 11742
rect 11702 11544 11758 11600
rect 11844 11544 11900 11600
rect 11702 11402 11758 11458
rect 11844 11402 11900 11458
rect 11702 11260 11758 11316
rect 11844 11260 11900 11316
rect 11702 11118 11758 11174
rect 11844 11118 11900 11174
rect 11702 10976 11758 11032
rect 11844 10976 11900 11032
rect 11702 10834 11758 10890
rect 11844 10834 11900 10890
rect 11702 10692 11758 10748
rect 11844 10692 11900 10748
rect 11702 10550 11758 10606
rect 11844 10550 11900 10606
rect 11702 10408 11758 10464
rect 11844 10408 11900 10464
rect 11702 10266 11758 10322
rect 11844 10266 11900 10322
rect 11702 10124 11758 10180
rect 11844 10124 11900 10180
rect 11702 9982 11758 10038
rect 11844 9982 11900 10038
rect 11702 9840 11758 9896
rect 11844 9840 11900 9896
rect 11702 9698 11758 9754
rect 11844 9698 11900 9754
rect 11702 9556 11758 9612
rect 11844 9556 11900 9612
rect 11702 9414 11758 9470
rect 11844 9414 11900 9470
rect 11702 9272 11758 9328
rect 11844 9272 11900 9328
rect 11702 9130 11758 9186
rect 11844 9130 11900 9186
rect 11702 8988 11758 9044
rect 11844 8988 11900 9044
rect 11702 8846 11758 8902
rect 11844 8846 11900 8902
rect 11702 8704 11758 8760
rect 11844 8704 11900 8760
rect 11702 8562 11758 8618
rect 11844 8562 11900 8618
rect 11702 8420 11758 8476
rect 11844 8420 11900 8476
rect 11702 8278 11758 8334
rect 11844 8278 11900 8334
rect 11702 8136 11758 8192
rect 11844 8136 11900 8192
rect 11702 7994 11758 8050
rect 11844 7994 11900 8050
rect 11702 7852 11758 7908
rect 11844 7852 11900 7908
rect 11702 7710 11758 7766
rect 11844 7710 11900 7766
rect 11702 7568 11758 7624
rect 11844 7568 11900 7624
rect 11702 7426 11758 7482
rect 11844 7426 11900 7482
rect 11702 7284 11758 7340
rect 11844 7284 11900 7340
rect 11702 7142 11758 7198
rect 11844 7142 11900 7198
rect 11702 7000 11758 7056
rect 11844 7000 11900 7056
rect 11702 6858 11758 6914
rect 11844 6858 11900 6914
rect 11702 6716 11758 6772
rect 11844 6716 11900 6772
rect 11702 6574 11758 6630
rect 11844 6574 11900 6630
rect 11702 6432 11758 6488
rect 11844 6432 11900 6488
rect 11702 6290 11758 6346
rect 11844 6290 11900 6346
rect 11702 6148 11758 6204
rect 11844 6148 11900 6204
rect 11702 6006 11758 6062
rect 11844 6006 11900 6062
rect 11702 5864 11758 5920
rect 11844 5864 11900 5920
rect 11702 5722 11758 5778
rect 11844 5722 11900 5778
rect 11702 5580 11758 5636
rect 11844 5580 11900 5636
rect 11702 5438 11758 5494
rect 11844 5438 11900 5494
rect 11702 5296 11758 5352
rect 11844 5296 11900 5352
rect 11702 5154 11758 5210
rect 11844 5154 11900 5210
rect 11702 5012 11758 5068
rect 11844 5012 11900 5068
rect 11702 4870 11758 4926
rect 11844 4870 11900 4926
rect 11702 4728 11758 4784
rect 11844 4728 11900 4784
rect 11702 4586 11758 4642
rect 11844 4586 11900 4642
rect 11702 4444 11758 4500
rect 11844 4444 11900 4500
rect 11702 4302 11758 4358
rect 11844 4302 11900 4358
rect 11702 4160 11758 4216
rect 11844 4160 11900 4216
rect 11702 4018 11758 4074
rect 11844 4018 11900 4074
rect 11702 3876 11758 3932
rect 11844 3876 11900 3932
rect 11702 3734 11758 3790
rect 11844 3734 11900 3790
rect 11702 3592 11758 3648
rect 11844 3592 11900 3648
rect 11702 3450 11758 3506
rect 11844 3450 11900 3506
rect 11702 3308 11758 3364
rect 11844 3308 11900 3364
rect 11702 3166 11758 3222
rect 11844 3166 11900 3222
rect 11702 3024 11758 3080
rect 11844 3024 11900 3080
rect 11702 2882 11758 2938
rect 11844 2882 11900 2938
rect 11702 2740 11758 2796
rect 11844 2740 11900 2796
rect 11702 2598 11758 2654
rect 11844 2598 11900 2654
rect 11702 2456 11758 2512
rect 11844 2456 11900 2512
rect 11702 2314 11758 2370
rect 11844 2314 11900 2370
rect 11702 2172 11758 2228
rect 11844 2172 11900 2228
rect 11702 2030 11758 2086
rect 11844 2030 11900 2086
rect 11702 1888 11758 1944
rect 11844 1888 11900 1944
rect 11702 1746 11758 1802
rect 11844 1746 11900 1802
rect 11702 1604 11758 1660
rect 11844 1604 11900 1660
rect 11702 1462 11758 1518
rect 11844 1462 11900 1518
rect 11702 1320 11758 1376
rect 11844 1320 11900 1376
rect 11702 1178 11758 1234
rect 11844 1178 11900 1234
rect 11702 1036 11758 1092
rect 11844 1036 11900 1092
rect 11702 894 11758 950
rect 11844 894 11900 950
rect 11702 752 11758 808
rect 11844 752 11900 808
rect 11702 610 11758 666
rect 11844 610 11900 666
rect 11702 468 11758 524
rect 11844 468 11900 524
rect 12526 12302 12582 12358
rect 12650 12302 12706 12358
rect 12774 12302 12830 12358
rect 12898 12302 12954 12358
rect 13022 12302 13078 12358
rect 12526 12178 12582 12234
rect 12650 12178 12706 12234
rect 12774 12178 12830 12234
rect 12898 12178 12954 12234
rect 13022 12178 13078 12234
rect 12526 12054 12582 12110
rect 12650 12054 12706 12110
rect 12774 12054 12830 12110
rect 12898 12054 12954 12110
rect 13022 12054 13078 12110
rect 12526 11930 12582 11986
rect 12650 11930 12706 11986
rect 12774 11930 12830 11986
rect 12898 11930 12954 11986
rect 13022 11930 13078 11986
rect 12526 11806 12582 11862
rect 12650 11806 12706 11862
rect 12774 11806 12830 11862
rect 12898 11806 12954 11862
rect 13022 11806 13078 11862
rect 12526 11682 12582 11738
rect 12650 11682 12706 11738
rect 12774 11682 12830 11738
rect 12898 11682 12954 11738
rect 13022 11682 13078 11738
rect 12526 11558 12582 11614
rect 12650 11558 12706 11614
rect 12774 11558 12830 11614
rect 12898 11558 12954 11614
rect 13022 11558 13078 11614
rect 12526 11434 12582 11490
rect 12650 11434 12706 11490
rect 12774 11434 12830 11490
rect 12898 11434 12954 11490
rect 13022 11434 13078 11490
rect 12526 11310 12582 11366
rect 12650 11310 12706 11366
rect 12774 11310 12830 11366
rect 12898 11310 12954 11366
rect 13022 11310 13078 11366
rect 12526 11186 12582 11242
rect 12650 11186 12706 11242
rect 12774 11186 12830 11242
rect 12898 11186 12954 11242
rect 13022 11186 13078 11242
rect 12526 11062 12582 11118
rect 12650 11062 12706 11118
rect 12774 11062 12830 11118
rect 12898 11062 12954 11118
rect 13022 11062 13078 11118
rect 12526 10938 12582 10994
rect 12650 10938 12706 10994
rect 12774 10938 12830 10994
rect 12898 10938 12954 10994
rect 13022 10938 13078 10994
rect 12526 10814 12582 10870
rect 12650 10814 12706 10870
rect 12774 10814 12830 10870
rect 12898 10814 12954 10870
rect 13022 10814 13078 10870
rect 12526 10690 12582 10746
rect 12650 10690 12706 10746
rect 12774 10690 12830 10746
rect 12898 10690 12954 10746
rect 13022 10690 13078 10746
rect 12526 10566 12582 10622
rect 12650 10566 12706 10622
rect 12774 10566 12830 10622
rect 12898 10566 12954 10622
rect 13022 10566 13078 10622
rect 12526 10442 12582 10498
rect 12650 10442 12706 10498
rect 12774 10442 12830 10498
rect 12898 10442 12954 10498
rect 13022 10442 13078 10498
rect 12526 10318 12582 10374
rect 12650 10318 12706 10374
rect 12774 10318 12830 10374
rect 12898 10318 12954 10374
rect 13022 10318 13078 10374
rect 12526 10194 12582 10250
rect 12650 10194 12706 10250
rect 12774 10194 12830 10250
rect 12898 10194 12954 10250
rect 13022 10194 13078 10250
rect 12526 10070 12582 10126
rect 12650 10070 12706 10126
rect 12774 10070 12830 10126
rect 12898 10070 12954 10126
rect 13022 10070 13078 10126
rect 12526 9946 12582 10002
rect 12650 9946 12706 10002
rect 12774 9946 12830 10002
rect 12898 9946 12954 10002
rect 13022 9946 13078 10002
rect 12526 9822 12582 9878
rect 12650 9822 12706 9878
rect 12774 9822 12830 9878
rect 12898 9822 12954 9878
rect 13022 9822 13078 9878
rect 12526 9698 12582 9754
rect 12650 9698 12706 9754
rect 12774 9698 12830 9754
rect 12898 9698 12954 9754
rect 13022 9698 13078 9754
rect 12526 9574 12582 9630
rect 12650 9574 12706 9630
rect 12774 9574 12830 9630
rect 12898 9574 12954 9630
rect 13022 9574 13078 9630
rect 12526 9450 12582 9506
rect 12650 9450 12706 9506
rect 12774 9450 12830 9506
rect 12898 9450 12954 9506
rect 13022 9450 13078 9506
rect 12526 9326 12582 9382
rect 12650 9326 12706 9382
rect 12774 9326 12830 9382
rect 12898 9326 12954 9382
rect 13022 9326 13078 9382
rect 12526 9202 12582 9258
rect 12650 9202 12706 9258
rect 12774 9202 12830 9258
rect 12898 9202 12954 9258
rect 13022 9202 13078 9258
rect 12526 9078 12582 9134
rect 12650 9078 12706 9134
rect 12774 9078 12830 9134
rect 12898 9078 12954 9134
rect 13022 9078 13078 9134
rect 12526 8954 12582 9010
rect 12650 8954 12706 9010
rect 12774 8954 12830 9010
rect 12898 8954 12954 9010
rect 13022 8954 13078 9010
rect 12526 8830 12582 8886
rect 12650 8830 12706 8886
rect 12774 8830 12830 8886
rect 12898 8830 12954 8886
rect 13022 8830 13078 8886
rect 12526 8706 12582 8762
rect 12650 8706 12706 8762
rect 12774 8706 12830 8762
rect 12898 8706 12954 8762
rect 13022 8706 13078 8762
rect 12526 8582 12582 8638
rect 12650 8582 12706 8638
rect 12774 8582 12830 8638
rect 12898 8582 12954 8638
rect 13022 8582 13078 8638
rect 12526 8458 12582 8514
rect 12650 8458 12706 8514
rect 12774 8458 12830 8514
rect 12898 8458 12954 8514
rect 13022 8458 13078 8514
rect 12526 8334 12582 8390
rect 12650 8334 12706 8390
rect 12774 8334 12830 8390
rect 12898 8334 12954 8390
rect 13022 8334 13078 8390
rect 12526 8210 12582 8266
rect 12650 8210 12706 8266
rect 12774 8210 12830 8266
rect 12898 8210 12954 8266
rect 13022 8210 13078 8266
rect 12526 8086 12582 8142
rect 12650 8086 12706 8142
rect 12774 8086 12830 8142
rect 12898 8086 12954 8142
rect 13022 8086 13078 8142
rect 12526 7962 12582 8018
rect 12650 7962 12706 8018
rect 12774 7962 12830 8018
rect 12898 7962 12954 8018
rect 13022 7962 13078 8018
rect 12526 7838 12582 7894
rect 12650 7838 12706 7894
rect 12774 7838 12830 7894
rect 12898 7838 12954 7894
rect 13022 7838 13078 7894
rect 12526 7714 12582 7770
rect 12650 7714 12706 7770
rect 12774 7714 12830 7770
rect 12898 7714 12954 7770
rect 13022 7714 13078 7770
rect 12526 7590 12582 7646
rect 12650 7590 12706 7646
rect 12774 7590 12830 7646
rect 12898 7590 12954 7646
rect 13022 7590 13078 7646
rect 12526 7466 12582 7522
rect 12650 7466 12706 7522
rect 12774 7466 12830 7522
rect 12898 7466 12954 7522
rect 13022 7466 13078 7522
rect 12526 7342 12582 7398
rect 12650 7342 12706 7398
rect 12774 7342 12830 7398
rect 12898 7342 12954 7398
rect 13022 7342 13078 7398
rect 12526 7218 12582 7274
rect 12650 7218 12706 7274
rect 12774 7218 12830 7274
rect 12898 7218 12954 7274
rect 13022 7218 13078 7274
rect 12526 7094 12582 7150
rect 12650 7094 12706 7150
rect 12774 7094 12830 7150
rect 12898 7094 12954 7150
rect 13022 7094 13078 7150
rect 12526 6970 12582 7026
rect 12650 6970 12706 7026
rect 12774 6970 12830 7026
rect 12898 6970 12954 7026
rect 13022 6970 13078 7026
rect 12526 6846 12582 6902
rect 12650 6846 12706 6902
rect 12774 6846 12830 6902
rect 12898 6846 12954 6902
rect 13022 6846 13078 6902
rect 12526 6722 12582 6778
rect 12650 6722 12706 6778
rect 12774 6722 12830 6778
rect 12898 6722 12954 6778
rect 13022 6722 13078 6778
rect 12526 6598 12582 6654
rect 12650 6598 12706 6654
rect 12774 6598 12830 6654
rect 12898 6598 12954 6654
rect 13022 6598 13078 6654
rect 12526 6474 12582 6530
rect 12650 6474 12706 6530
rect 12774 6474 12830 6530
rect 12898 6474 12954 6530
rect 13022 6474 13078 6530
rect 12526 6350 12582 6406
rect 12650 6350 12706 6406
rect 12774 6350 12830 6406
rect 12898 6350 12954 6406
rect 13022 6350 13078 6406
rect 12526 6226 12582 6282
rect 12650 6226 12706 6282
rect 12774 6226 12830 6282
rect 12898 6226 12954 6282
rect 13022 6226 13078 6282
rect 12526 6102 12582 6158
rect 12650 6102 12706 6158
rect 12774 6102 12830 6158
rect 12898 6102 12954 6158
rect 13022 6102 13078 6158
rect 12526 5978 12582 6034
rect 12650 5978 12706 6034
rect 12774 5978 12830 6034
rect 12898 5978 12954 6034
rect 13022 5978 13078 6034
rect 12526 5854 12582 5910
rect 12650 5854 12706 5910
rect 12774 5854 12830 5910
rect 12898 5854 12954 5910
rect 13022 5854 13078 5910
rect 12526 5730 12582 5786
rect 12650 5730 12706 5786
rect 12774 5730 12830 5786
rect 12898 5730 12954 5786
rect 13022 5730 13078 5786
rect 12526 5606 12582 5662
rect 12650 5606 12706 5662
rect 12774 5606 12830 5662
rect 12898 5606 12954 5662
rect 13022 5606 13078 5662
rect 12526 5482 12582 5538
rect 12650 5482 12706 5538
rect 12774 5482 12830 5538
rect 12898 5482 12954 5538
rect 13022 5482 13078 5538
rect 12526 5358 12582 5414
rect 12650 5358 12706 5414
rect 12774 5358 12830 5414
rect 12898 5358 12954 5414
rect 13022 5358 13078 5414
rect 12526 5234 12582 5290
rect 12650 5234 12706 5290
rect 12774 5234 12830 5290
rect 12898 5234 12954 5290
rect 13022 5234 13078 5290
rect 12526 5110 12582 5166
rect 12650 5110 12706 5166
rect 12774 5110 12830 5166
rect 12898 5110 12954 5166
rect 13022 5110 13078 5166
rect 12526 4986 12582 5042
rect 12650 4986 12706 5042
rect 12774 4986 12830 5042
rect 12898 4986 12954 5042
rect 13022 4986 13078 5042
rect 12526 4862 12582 4918
rect 12650 4862 12706 4918
rect 12774 4862 12830 4918
rect 12898 4862 12954 4918
rect 13022 4862 13078 4918
rect 12526 4738 12582 4794
rect 12650 4738 12706 4794
rect 12774 4738 12830 4794
rect 12898 4738 12954 4794
rect 13022 4738 13078 4794
rect 12526 4614 12582 4670
rect 12650 4614 12706 4670
rect 12774 4614 12830 4670
rect 12898 4614 12954 4670
rect 13022 4614 13078 4670
rect 12526 4490 12582 4546
rect 12650 4490 12706 4546
rect 12774 4490 12830 4546
rect 12898 4490 12954 4546
rect 13022 4490 13078 4546
rect 12526 4366 12582 4422
rect 12650 4366 12706 4422
rect 12774 4366 12830 4422
rect 12898 4366 12954 4422
rect 13022 4366 13078 4422
rect 12526 4242 12582 4298
rect 12650 4242 12706 4298
rect 12774 4242 12830 4298
rect 12898 4242 12954 4298
rect 13022 4242 13078 4298
rect 12526 4118 12582 4174
rect 12650 4118 12706 4174
rect 12774 4118 12830 4174
rect 12898 4118 12954 4174
rect 13022 4118 13078 4174
rect 12526 3994 12582 4050
rect 12650 3994 12706 4050
rect 12774 3994 12830 4050
rect 12898 3994 12954 4050
rect 13022 3994 13078 4050
rect 12526 3870 12582 3926
rect 12650 3870 12706 3926
rect 12774 3870 12830 3926
rect 12898 3870 12954 3926
rect 13022 3870 13078 3926
rect 12526 3746 12582 3802
rect 12650 3746 12706 3802
rect 12774 3746 12830 3802
rect 12898 3746 12954 3802
rect 13022 3746 13078 3802
rect 12526 3622 12582 3678
rect 12650 3622 12706 3678
rect 12774 3622 12830 3678
rect 12898 3622 12954 3678
rect 13022 3622 13078 3678
rect 12526 3498 12582 3554
rect 12650 3498 12706 3554
rect 12774 3498 12830 3554
rect 12898 3498 12954 3554
rect 13022 3498 13078 3554
rect 12526 3374 12582 3430
rect 12650 3374 12706 3430
rect 12774 3374 12830 3430
rect 12898 3374 12954 3430
rect 13022 3374 13078 3430
rect 12526 3250 12582 3306
rect 12650 3250 12706 3306
rect 12774 3250 12830 3306
rect 12898 3250 12954 3306
rect 13022 3250 13078 3306
rect 12526 3126 12582 3182
rect 12650 3126 12706 3182
rect 12774 3126 12830 3182
rect 12898 3126 12954 3182
rect 13022 3126 13078 3182
rect 12526 3002 12582 3058
rect 12650 3002 12706 3058
rect 12774 3002 12830 3058
rect 12898 3002 12954 3058
rect 13022 3002 13078 3058
rect 12526 2878 12582 2934
rect 12650 2878 12706 2934
rect 12774 2878 12830 2934
rect 12898 2878 12954 2934
rect 13022 2878 13078 2934
rect 12526 2754 12582 2810
rect 12650 2754 12706 2810
rect 12774 2754 12830 2810
rect 12898 2754 12954 2810
rect 13022 2754 13078 2810
rect 12526 2630 12582 2686
rect 12650 2630 12706 2686
rect 12774 2630 12830 2686
rect 12898 2630 12954 2686
rect 13022 2630 13078 2686
rect 12526 2506 12582 2562
rect 12650 2506 12706 2562
rect 12774 2506 12830 2562
rect 12898 2506 12954 2562
rect 13022 2506 13078 2562
rect 12526 2382 12582 2438
rect 12650 2382 12706 2438
rect 12774 2382 12830 2438
rect 12898 2382 12954 2438
rect 13022 2382 13078 2438
rect 12526 2258 12582 2314
rect 12650 2258 12706 2314
rect 12774 2258 12830 2314
rect 12898 2258 12954 2314
rect 13022 2258 13078 2314
rect 12526 2134 12582 2190
rect 12650 2134 12706 2190
rect 12774 2134 12830 2190
rect 12898 2134 12954 2190
rect 13022 2134 13078 2190
rect 12526 2010 12582 2066
rect 12650 2010 12706 2066
rect 12774 2010 12830 2066
rect 12898 2010 12954 2066
rect 13022 2010 13078 2066
rect 12526 1886 12582 1942
rect 12650 1886 12706 1942
rect 12774 1886 12830 1942
rect 12898 1886 12954 1942
rect 13022 1886 13078 1942
rect 12526 1762 12582 1818
rect 12650 1762 12706 1818
rect 12774 1762 12830 1818
rect 12898 1762 12954 1818
rect 13022 1762 13078 1818
rect 12526 1638 12582 1694
rect 12650 1638 12706 1694
rect 12774 1638 12830 1694
rect 12898 1638 12954 1694
rect 13022 1638 13078 1694
rect 12526 1514 12582 1570
rect 12650 1514 12706 1570
rect 12774 1514 12830 1570
rect 12898 1514 12954 1570
rect 13022 1514 13078 1570
rect 12526 1390 12582 1446
rect 12650 1390 12706 1446
rect 12774 1390 12830 1446
rect 12898 1390 12954 1446
rect 13022 1390 13078 1446
rect 12526 1266 12582 1322
rect 12650 1266 12706 1322
rect 12774 1266 12830 1322
rect 12898 1266 12954 1322
rect 13022 1266 13078 1322
rect 12526 1142 12582 1198
rect 12650 1142 12706 1198
rect 12774 1142 12830 1198
rect 12898 1142 12954 1198
rect 13022 1142 13078 1198
rect 12526 1018 12582 1074
rect 12650 1018 12706 1074
rect 12774 1018 12830 1074
rect 12898 1018 12954 1074
rect 13022 1018 13078 1074
rect 12526 894 12582 950
rect 12650 894 12706 950
rect 12774 894 12830 950
rect 12898 894 12954 950
rect 13022 894 13078 950
rect 12526 770 12582 826
rect 12650 770 12706 826
rect 12774 770 12830 826
rect 12898 770 12954 826
rect 13022 770 13078 826
rect 12526 646 12582 702
rect 12650 646 12706 702
rect 12774 646 12830 702
rect 12898 646 12954 702
rect 13022 646 13078 702
rect 12526 522 12582 578
rect 12650 522 12706 578
rect 12774 522 12830 578
rect 12898 522 12954 578
rect 13022 522 13078 578
rect -286 398 -230 454
rect -162 398 -106 454
rect -38 398 18 454
rect 86 398 142 454
rect 210 398 266 454
rect 12526 398 12582 454
rect 12650 398 12706 454
rect 12774 398 12830 454
rect 12898 398 12954 454
rect 13022 398 13078 454
rect -286 274 -230 330
rect -162 274 -106 330
rect -38 274 18 330
rect 86 274 142 330
rect 210 274 266 330
rect 415 246 471 302
rect 557 246 613 302
rect 699 246 755 302
rect 841 246 897 302
rect 983 246 1039 302
rect 1125 246 1181 302
rect 1267 246 1323 302
rect 1409 246 1465 302
rect 1551 246 1607 302
rect 1693 246 1749 302
rect 1835 246 1891 302
rect 1977 246 2033 302
rect 2119 246 2175 302
rect 2261 246 2317 302
rect 2403 246 2459 302
rect 2545 246 2601 302
rect 2687 246 2743 302
rect 2829 246 2885 302
rect 2971 246 3027 302
rect 3113 246 3169 302
rect 3255 246 3311 302
rect 3397 246 3453 302
rect 3539 246 3595 302
rect 3681 246 3737 302
rect 3823 246 3879 302
rect 3965 246 4021 302
rect 4107 246 4163 302
rect 4249 246 4305 302
rect 4391 246 4447 302
rect 4533 246 4589 302
rect 4675 246 4731 302
rect 4817 246 4873 302
rect 4959 246 5015 302
rect 5101 246 5157 302
rect 5243 246 5299 302
rect 5385 246 5441 302
rect 5527 246 5583 302
rect 5669 246 5725 302
rect 5811 246 5867 302
rect 5953 246 6009 302
rect 6095 246 6151 302
rect 6237 246 6293 302
rect 6379 246 6435 302
rect 6521 246 6577 302
rect 6663 246 6719 302
rect 6805 246 6861 302
rect 6947 246 7003 302
rect 7089 246 7145 302
rect 7231 246 7287 302
rect 7373 246 7429 302
rect 7515 246 7571 302
rect 7657 246 7713 302
rect 7799 246 7855 302
rect 7941 246 7997 302
rect 8083 246 8139 302
rect 8225 246 8281 302
rect 8367 246 8423 302
rect 8509 246 8565 302
rect 8651 246 8707 302
rect 8793 246 8849 302
rect 8935 246 8991 302
rect 9077 246 9133 302
rect 9219 246 9275 302
rect 9361 246 9417 302
rect 9503 246 9559 302
rect 9645 246 9701 302
rect 9787 246 9843 302
rect 9929 246 9985 302
rect 10071 246 10127 302
rect 10213 246 10269 302
rect 10355 246 10411 302
rect 10497 246 10553 302
rect 10639 246 10695 302
rect 10781 246 10837 302
rect 10923 246 10979 302
rect 11065 246 11121 302
rect 11207 246 11263 302
rect 11349 246 11405 302
rect 11491 246 11547 302
rect 11633 246 11689 302
rect 11775 246 11831 302
rect 11917 246 11973 302
rect 12059 246 12115 302
rect 12201 246 12257 302
rect 12343 246 12399 302
rect 12526 274 12582 330
rect 12650 274 12706 330
rect 12774 274 12830 330
rect 12898 274 12954 330
rect 13022 274 13078 330
rect -286 150 -230 206
rect -162 150 -106 206
rect -38 150 18 206
rect 86 150 142 206
rect 210 150 266 206
rect 415 104 471 160
rect 557 104 613 160
rect 699 104 755 160
rect 841 104 897 160
rect 983 104 1039 160
rect 1125 104 1181 160
rect 1267 104 1323 160
rect 1409 104 1465 160
rect 1551 104 1607 160
rect 1693 104 1749 160
rect 1835 104 1891 160
rect 1977 104 2033 160
rect 2119 104 2175 160
rect 2261 104 2317 160
rect 2403 104 2459 160
rect 2545 104 2601 160
rect 2687 104 2743 160
rect 2829 104 2885 160
rect 2971 104 3027 160
rect 3113 104 3169 160
rect 3255 104 3311 160
rect 3397 104 3453 160
rect 3539 104 3595 160
rect 3681 104 3737 160
rect 3823 104 3879 160
rect 3965 104 4021 160
rect 4107 104 4163 160
rect 4249 104 4305 160
rect 4391 104 4447 160
rect 4533 104 4589 160
rect 4675 104 4731 160
rect 4817 104 4873 160
rect 4959 104 5015 160
rect 5101 104 5157 160
rect 5243 104 5299 160
rect 5385 104 5441 160
rect 5527 104 5583 160
rect 5669 104 5725 160
rect 5811 104 5867 160
rect 5953 104 6009 160
rect 6095 104 6151 160
rect 6237 104 6293 160
rect 6379 104 6435 160
rect 6521 104 6577 160
rect 6663 104 6719 160
rect 6805 104 6861 160
rect 6947 104 7003 160
rect 7089 104 7145 160
rect 7231 104 7287 160
rect 7373 104 7429 160
rect 7515 104 7571 160
rect 7657 104 7713 160
rect 7799 104 7855 160
rect 7941 104 7997 160
rect 8083 104 8139 160
rect 8225 104 8281 160
rect 8367 104 8423 160
rect 8509 104 8565 160
rect 8651 104 8707 160
rect 8793 104 8849 160
rect 8935 104 8991 160
rect 9077 104 9133 160
rect 9219 104 9275 160
rect 9361 104 9417 160
rect 9503 104 9559 160
rect 9645 104 9701 160
rect 9787 104 9843 160
rect 9929 104 9985 160
rect 10071 104 10127 160
rect 10213 104 10269 160
rect 10355 104 10411 160
rect 10497 104 10553 160
rect 10639 104 10695 160
rect 10781 104 10837 160
rect 10923 104 10979 160
rect 11065 104 11121 160
rect 11207 104 11263 160
rect 11349 104 11405 160
rect 11491 104 11547 160
rect 11633 104 11689 160
rect 11775 104 11831 160
rect 11917 104 11973 160
rect 12059 104 12115 160
rect 12201 104 12257 160
rect 12343 104 12399 160
rect 12526 150 12582 206
rect 12650 150 12706 206
rect 12774 150 12830 206
rect 12898 150 12954 206
rect 13022 150 13078 206
<< metal4 >>
rect -400 12949 13200 13065
rect -400 12893 -254 12949
rect -198 12893 -130 12949
rect -74 12893 -6 12949
rect 50 12893 118 12949
rect 174 12893 242 12949
rect 298 12893 366 12949
rect 422 12893 490 12949
rect 546 12893 614 12949
rect 670 12893 738 12949
rect 794 12893 862 12949
rect 918 12893 986 12949
rect 1042 12893 1110 12949
rect 1166 12893 1234 12949
rect 1290 12893 1358 12949
rect 1414 12893 1482 12949
rect 1538 12893 1606 12949
rect 1662 12893 1730 12949
rect 1786 12893 1854 12949
rect 1910 12893 1978 12949
rect 2034 12893 2102 12949
rect 2158 12893 2226 12949
rect 2282 12893 2350 12949
rect 2406 12893 2474 12949
rect 2530 12893 2598 12949
rect 2654 12893 2722 12949
rect 2778 12893 2846 12949
rect 2902 12893 2970 12949
rect 3026 12893 3094 12949
rect 3150 12893 3218 12949
rect 3274 12893 3342 12949
rect 3398 12893 3466 12949
rect 3522 12893 3590 12949
rect 3646 12893 3714 12949
rect 3770 12893 3838 12949
rect 3894 12893 3962 12949
rect 4018 12893 4086 12949
rect 4142 12893 4210 12949
rect 4266 12893 4334 12949
rect 4390 12893 4458 12949
rect 4514 12893 4582 12949
rect 4638 12893 4706 12949
rect 4762 12893 4830 12949
rect 4886 12893 4954 12949
rect 5010 12893 5078 12949
rect 5134 12893 5202 12949
rect 5258 12893 5326 12949
rect 5382 12893 5450 12949
rect 5506 12893 5574 12949
rect 5630 12893 5698 12949
rect 5754 12893 5822 12949
rect 5878 12893 5946 12949
rect 6002 12893 6070 12949
rect 6126 12893 6194 12949
rect 6250 12893 6318 12949
rect 6374 12893 6442 12949
rect 6498 12893 6566 12949
rect 6622 12893 6690 12949
rect 6746 12893 6814 12949
rect 6870 12893 6938 12949
rect 6994 12893 7062 12949
rect 7118 12893 7186 12949
rect 7242 12893 7310 12949
rect 7366 12893 7434 12949
rect 7490 12893 7558 12949
rect 7614 12893 7682 12949
rect 7738 12893 7806 12949
rect 7862 12893 7930 12949
rect 7986 12893 8054 12949
rect 8110 12893 8178 12949
rect 8234 12893 8302 12949
rect 8358 12893 8426 12949
rect 8482 12893 8550 12949
rect 8606 12893 8674 12949
rect 8730 12893 8798 12949
rect 8854 12893 8922 12949
rect 8978 12893 9046 12949
rect 9102 12893 9170 12949
rect 9226 12893 9294 12949
rect 9350 12893 9418 12949
rect 9474 12893 9542 12949
rect 9598 12893 9666 12949
rect 9722 12893 9790 12949
rect 9846 12893 9914 12949
rect 9970 12893 10038 12949
rect 10094 12893 10162 12949
rect 10218 12893 10286 12949
rect 10342 12893 10410 12949
rect 10466 12893 10534 12949
rect 10590 12893 10658 12949
rect 10714 12893 10782 12949
rect 10838 12893 10906 12949
rect 10962 12893 11030 12949
rect 11086 12893 11154 12949
rect 11210 12893 11278 12949
rect 11334 12893 11402 12949
rect 11458 12893 11526 12949
rect 11582 12893 11650 12949
rect 11706 12893 11774 12949
rect 11830 12893 11898 12949
rect 11954 12893 12022 12949
rect 12078 12893 12146 12949
rect 12202 12893 12270 12949
rect 12326 12893 12394 12949
rect 12450 12893 12518 12949
rect 12574 12893 12642 12949
rect 12698 12893 12766 12949
rect 12822 12893 12890 12949
rect 12946 12893 13014 12949
rect 13070 12893 13200 12949
rect -400 12825 13200 12893
rect -400 12769 -254 12825
rect -198 12769 -130 12825
rect -74 12769 -6 12825
rect 50 12769 118 12825
rect 174 12769 242 12825
rect 298 12769 366 12825
rect 422 12769 490 12825
rect 546 12769 614 12825
rect 670 12769 738 12825
rect 794 12769 862 12825
rect 918 12769 986 12825
rect 1042 12769 1110 12825
rect 1166 12769 1234 12825
rect 1290 12769 1358 12825
rect 1414 12769 1482 12825
rect 1538 12769 1606 12825
rect 1662 12769 1730 12825
rect 1786 12769 1854 12825
rect 1910 12769 1978 12825
rect 2034 12769 2102 12825
rect 2158 12769 2226 12825
rect 2282 12769 2350 12825
rect 2406 12769 2474 12825
rect 2530 12769 2598 12825
rect 2654 12769 2722 12825
rect 2778 12769 2846 12825
rect 2902 12769 2970 12825
rect 3026 12769 3094 12825
rect 3150 12769 3218 12825
rect 3274 12769 3342 12825
rect 3398 12769 3466 12825
rect 3522 12769 3590 12825
rect 3646 12769 3714 12825
rect 3770 12769 3838 12825
rect 3894 12769 3962 12825
rect 4018 12769 4086 12825
rect 4142 12769 4210 12825
rect 4266 12769 4334 12825
rect 4390 12769 4458 12825
rect 4514 12769 4582 12825
rect 4638 12769 4706 12825
rect 4762 12769 4830 12825
rect 4886 12769 4954 12825
rect 5010 12769 5078 12825
rect 5134 12769 5202 12825
rect 5258 12769 5326 12825
rect 5382 12769 5450 12825
rect 5506 12769 5574 12825
rect 5630 12769 5698 12825
rect 5754 12769 5822 12825
rect 5878 12769 5946 12825
rect 6002 12769 6070 12825
rect 6126 12769 6194 12825
rect 6250 12769 6318 12825
rect 6374 12769 6442 12825
rect 6498 12769 6566 12825
rect 6622 12769 6690 12825
rect 6746 12769 6814 12825
rect 6870 12769 6938 12825
rect 6994 12769 7062 12825
rect 7118 12769 7186 12825
rect 7242 12769 7310 12825
rect 7366 12769 7434 12825
rect 7490 12769 7558 12825
rect 7614 12769 7682 12825
rect 7738 12769 7806 12825
rect 7862 12769 7930 12825
rect 7986 12769 8054 12825
rect 8110 12769 8178 12825
rect 8234 12769 8302 12825
rect 8358 12769 8426 12825
rect 8482 12769 8550 12825
rect 8606 12769 8674 12825
rect 8730 12769 8798 12825
rect 8854 12769 8922 12825
rect 8978 12769 9046 12825
rect 9102 12769 9170 12825
rect 9226 12769 9294 12825
rect 9350 12769 9418 12825
rect 9474 12769 9542 12825
rect 9598 12769 9666 12825
rect 9722 12769 9790 12825
rect 9846 12769 9914 12825
rect 9970 12769 10038 12825
rect 10094 12769 10162 12825
rect 10218 12769 10286 12825
rect 10342 12769 10410 12825
rect 10466 12769 10534 12825
rect 10590 12769 10658 12825
rect 10714 12769 10782 12825
rect 10838 12769 10906 12825
rect 10962 12769 11030 12825
rect 11086 12769 11154 12825
rect 11210 12769 11278 12825
rect 11334 12769 11402 12825
rect 11458 12769 11526 12825
rect 11582 12769 11650 12825
rect 11706 12769 11774 12825
rect 11830 12769 11898 12825
rect 11954 12769 12022 12825
rect 12078 12769 12146 12825
rect 12202 12769 12270 12825
rect 12326 12769 12394 12825
rect 12450 12769 12518 12825
rect 12574 12769 12642 12825
rect 12698 12769 12766 12825
rect 12822 12769 12890 12825
rect 12946 12769 13014 12825
rect 13070 12769 13200 12825
rect -400 12701 13200 12769
rect -400 12645 -254 12701
rect -198 12645 -130 12701
rect -74 12645 -6 12701
rect 50 12645 118 12701
rect 174 12645 242 12701
rect 298 12645 366 12701
rect 422 12645 490 12701
rect 546 12645 614 12701
rect 670 12645 738 12701
rect 794 12645 862 12701
rect 918 12645 986 12701
rect 1042 12645 1110 12701
rect 1166 12645 1234 12701
rect 1290 12645 1358 12701
rect 1414 12645 1482 12701
rect 1538 12645 1606 12701
rect 1662 12645 1730 12701
rect 1786 12645 1854 12701
rect 1910 12645 1978 12701
rect 2034 12645 2102 12701
rect 2158 12645 2226 12701
rect 2282 12645 2350 12701
rect 2406 12645 2474 12701
rect 2530 12645 2598 12701
rect 2654 12645 2722 12701
rect 2778 12645 2846 12701
rect 2902 12645 2970 12701
rect 3026 12645 3094 12701
rect 3150 12645 3218 12701
rect 3274 12645 3342 12701
rect 3398 12645 3466 12701
rect 3522 12645 3590 12701
rect 3646 12645 3714 12701
rect 3770 12645 3838 12701
rect 3894 12645 3962 12701
rect 4018 12645 4086 12701
rect 4142 12645 4210 12701
rect 4266 12645 4334 12701
rect 4390 12645 4458 12701
rect 4514 12645 4582 12701
rect 4638 12645 4706 12701
rect 4762 12645 4830 12701
rect 4886 12645 4954 12701
rect 5010 12645 5078 12701
rect 5134 12645 5202 12701
rect 5258 12645 5326 12701
rect 5382 12645 5450 12701
rect 5506 12645 5574 12701
rect 5630 12645 5698 12701
rect 5754 12645 5822 12701
rect 5878 12645 5946 12701
rect 6002 12645 6070 12701
rect 6126 12645 6194 12701
rect 6250 12645 6318 12701
rect 6374 12645 6442 12701
rect 6498 12645 6566 12701
rect 6622 12645 6690 12701
rect 6746 12645 6814 12701
rect 6870 12645 6938 12701
rect 6994 12645 7062 12701
rect 7118 12645 7186 12701
rect 7242 12645 7310 12701
rect 7366 12645 7434 12701
rect 7490 12645 7558 12701
rect 7614 12645 7682 12701
rect 7738 12645 7806 12701
rect 7862 12645 7930 12701
rect 7986 12645 8054 12701
rect 8110 12645 8178 12701
rect 8234 12645 8302 12701
rect 8358 12645 8426 12701
rect 8482 12645 8550 12701
rect 8606 12645 8674 12701
rect 8730 12645 8798 12701
rect 8854 12645 8922 12701
rect 8978 12645 9046 12701
rect 9102 12645 9170 12701
rect 9226 12645 9294 12701
rect 9350 12645 9418 12701
rect 9474 12645 9542 12701
rect 9598 12645 9666 12701
rect 9722 12645 9790 12701
rect 9846 12645 9914 12701
rect 9970 12645 10038 12701
rect 10094 12645 10162 12701
rect 10218 12645 10286 12701
rect 10342 12645 10410 12701
rect 10466 12645 10534 12701
rect 10590 12645 10658 12701
rect 10714 12645 10782 12701
rect 10838 12645 10906 12701
rect 10962 12645 11030 12701
rect 11086 12645 11154 12701
rect 11210 12645 11278 12701
rect 11334 12645 11402 12701
rect 11458 12645 11526 12701
rect 11582 12645 11650 12701
rect 11706 12645 11774 12701
rect 11830 12645 11898 12701
rect 11954 12645 12022 12701
rect 12078 12645 12146 12701
rect 12202 12645 12270 12701
rect 12326 12645 12394 12701
rect 12450 12645 12518 12701
rect 12574 12645 12642 12701
rect 12698 12645 12766 12701
rect 12822 12645 12890 12701
rect 12946 12645 13014 12701
rect 13070 12645 13200 12701
rect -400 12577 13200 12645
rect -400 12521 -254 12577
rect -198 12521 -130 12577
rect -74 12521 -6 12577
rect 50 12521 118 12577
rect 174 12521 242 12577
rect 298 12521 366 12577
rect 422 12521 490 12577
rect 546 12521 614 12577
rect 670 12521 738 12577
rect 794 12521 862 12577
rect 918 12521 986 12577
rect 1042 12521 1110 12577
rect 1166 12521 1234 12577
rect 1290 12521 1358 12577
rect 1414 12521 1482 12577
rect 1538 12521 1606 12577
rect 1662 12521 1730 12577
rect 1786 12521 1854 12577
rect 1910 12521 1978 12577
rect 2034 12521 2102 12577
rect 2158 12521 2226 12577
rect 2282 12521 2350 12577
rect 2406 12521 2474 12577
rect 2530 12521 2598 12577
rect 2654 12521 2722 12577
rect 2778 12521 2846 12577
rect 2902 12521 2970 12577
rect 3026 12521 3094 12577
rect 3150 12521 3218 12577
rect 3274 12521 3342 12577
rect 3398 12521 3466 12577
rect 3522 12521 3590 12577
rect 3646 12521 3714 12577
rect 3770 12521 3838 12577
rect 3894 12521 3962 12577
rect 4018 12521 4086 12577
rect 4142 12521 4210 12577
rect 4266 12521 4334 12577
rect 4390 12521 4458 12577
rect 4514 12521 4582 12577
rect 4638 12521 4706 12577
rect 4762 12521 4830 12577
rect 4886 12521 4954 12577
rect 5010 12521 5078 12577
rect 5134 12521 5202 12577
rect 5258 12521 5326 12577
rect 5382 12521 5450 12577
rect 5506 12521 5574 12577
rect 5630 12521 5698 12577
rect 5754 12521 5822 12577
rect 5878 12521 5946 12577
rect 6002 12521 6070 12577
rect 6126 12521 6194 12577
rect 6250 12521 6318 12577
rect 6374 12521 6442 12577
rect 6498 12521 6566 12577
rect 6622 12521 6690 12577
rect 6746 12521 6814 12577
rect 6870 12521 6938 12577
rect 6994 12521 7062 12577
rect 7118 12521 7186 12577
rect 7242 12521 7310 12577
rect 7366 12521 7434 12577
rect 7490 12521 7558 12577
rect 7614 12521 7682 12577
rect 7738 12521 7806 12577
rect 7862 12521 7930 12577
rect 7986 12521 8054 12577
rect 8110 12521 8178 12577
rect 8234 12521 8302 12577
rect 8358 12521 8426 12577
rect 8482 12521 8550 12577
rect 8606 12521 8674 12577
rect 8730 12521 8798 12577
rect 8854 12521 8922 12577
rect 8978 12521 9046 12577
rect 9102 12521 9170 12577
rect 9226 12521 9294 12577
rect 9350 12521 9418 12577
rect 9474 12521 9542 12577
rect 9598 12521 9666 12577
rect 9722 12521 9790 12577
rect 9846 12521 9914 12577
rect 9970 12521 10038 12577
rect 10094 12521 10162 12577
rect 10218 12521 10286 12577
rect 10342 12521 10410 12577
rect 10466 12521 10534 12577
rect 10590 12521 10658 12577
rect 10714 12521 10782 12577
rect 10838 12521 10906 12577
rect 10962 12521 11030 12577
rect 11086 12521 11154 12577
rect 11210 12521 11278 12577
rect 11334 12521 11402 12577
rect 11458 12521 11526 12577
rect 11582 12521 11650 12577
rect 11706 12521 11774 12577
rect 11830 12521 11898 12577
rect 11954 12521 12022 12577
rect 12078 12521 12146 12577
rect 12202 12521 12270 12577
rect 12326 12521 12394 12577
rect 12450 12521 12518 12577
rect 12574 12521 12642 12577
rect 12698 12521 12766 12577
rect 12822 12521 12890 12577
rect 12946 12521 13014 12577
rect 13070 12521 13200 12577
rect -400 12358 13200 12521
rect -400 12302 -286 12358
rect -230 12302 -162 12358
rect -106 12302 -38 12358
rect 18 12302 86 12358
rect 142 12302 210 12358
rect 266 12320 12526 12358
rect 266 12302 400 12320
rect -400 12234 400 12302
rect -400 12178 -286 12234
rect -230 12178 -162 12234
rect -106 12178 -38 12234
rect 18 12178 86 12234
rect 142 12178 210 12234
rect 266 12178 400 12234
rect -400 12110 400 12178
rect -400 12054 -286 12110
rect -230 12054 -162 12110
rect -106 12054 -38 12110
rect 18 12054 86 12110
rect 142 12054 210 12110
rect 266 12054 400 12110
rect -400 11986 400 12054
rect -400 11930 -286 11986
rect -230 11930 -162 11986
rect -106 11930 -38 11986
rect 18 11930 86 11986
rect 142 11930 210 11986
rect 266 11930 400 11986
rect -400 11862 400 11930
rect -400 11806 -286 11862
rect -230 11806 -162 11862
rect -106 11806 -38 11862
rect 18 11806 86 11862
rect 142 11806 210 11862
rect 266 11806 400 11862
rect -400 11738 400 11806
rect -400 11682 -286 11738
rect -230 11682 -162 11738
rect -106 11682 -38 11738
rect 18 11682 86 11738
rect 142 11682 210 11738
rect 266 11682 400 11738
rect -400 11614 400 11682
rect -400 11558 -286 11614
rect -230 11558 -162 11614
rect -106 11558 -38 11614
rect 18 11558 86 11614
rect 142 11558 210 11614
rect 266 11558 400 11614
rect -400 11490 400 11558
rect -400 11434 -286 11490
rect -230 11434 -162 11490
rect -106 11434 -38 11490
rect 18 11434 86 11490
rect 142 11434 210 11490
rect 266 11434 400 11490
rect -400 11366 400 11434
rect -400 11310 -286 11366
rect -230 11310 -162 11366
rect -106 11310 -38 11366
rect 18 11310 86 11366
rect 142 11310 210 11366
rect 266 11310 400 11366
rect -400 11242 400 11310
rect -400 11186 -286 11242
rect -230 11186 -162 11242
rect -106 11186 -38 11242
rect 18 11186 86 11242
rect 142 11186 210 11242
rect 266 11186 400 11242
rect -400 11118 400 11186
rect -400 11062 -286 11118
rect -230 11062 -162 11118
rect -106 11062 -38 11118
rect 18 11062 86 11118
rect 142 11062 210 11118
rect 266 11062 400 11118
rect -400 10994 400 11062
rect -400 10938 -286 10994
rect -230 10938 -162 10994
rect -106 10938 -38 10994
rect 18 10938 86 10994
rect 142 10938 210 10994
rect 266 10938 400 10994
rect -400 10870 400 10938
rect -400 10814 -286 10870
rect -230 10814 -162 10870
rect -106 10814 -38 10870
rect 18 10814 86 10870
rect 142 10814 210 10870
rect 266 10814 400 10870
rect -400 10746 400 10814
rect -400 10690 -286 10746
rect -230 10690 -162 10746
rect -106 10690 -38 10746
rect 18 10690 86 10746
rect 142 10690 210 10746
rect 266 10690 400 10746
rect -400 10622 400 10690
rect -400 10566 -286 10622
rect -230 10566 -162 10622
rect -106 10566 -38 10622
rect 18 10566 86 10622
rect 142 10566 210 10622
rect 266 10566 400 10622
rect -400 10498 400 10566
rect -400 10442 -286 10498
rect -230 10442 -162 10498
rect -106 10442 -38 10498
rect 18 10442 86 10498
rect 142 10442 210 10498
rect 266 10442 400 10498
rect -400 10374 400 10442
rect -400 10318 -286 10374
rect -230 10318 -162 10374
rect -106 10318 -38 10374
rect 18 10318 86 10374
rect 142 10318 210 10374
rect 266 10318 400 10374
rect -400 10250 400 10318
rect -400 10194 -286 10250
rect -230 10194 -162 10250
rect -106 10194 -38 10250
rect 18 10194 86 10250
rect 142 10194 210 10250
rect 266 10194 400 10250
rect -400 10126 400 10194
rect -400 10070 -286 10126
rect -230 10070 -162 10126
rect -106 10070 -38 10126
rect 18 10070 86 10126
rect 142 10070 210 10126
rect 266 10070 400 10126
rect -400 10002 400 10070
rect -400 9946 -286 10002
rect -230 9946 -162 10002
rect -106 9946 -38 10002
rect 18 9946 86 10002
rect 142 9946 210 10002
rect 266 9946 400 10002
rect -400 9878 400 9946
rect -400 9822 -286 9878
rect -230 9822 -162 9878
rect -106 9822 -38 9878
rect 18 9822 86 9878
rect 142 9822 210 9878
rect 266 9822 400 9878
rect -400 9754 400 9822
rect -400 9698 -286 9754
rect -230 9698 -162 9754
rect -106 9698 -38 9754
rect 18 9698 86 9754
rect 142 9698 210 9754
rect 266 9698 400 9754
rect -400 9630 400 9698
rect -400 9574 -286 9630
rect -230 9574 -162 9630
rect -106 9574 -38 9630
rect 18 9574 86 9630
rect 142 9574 210 9630
rect 266 9574 400 9630
rect -400 9506 400 9574
rect -400 9450 -286 9506
rect -230 9450 -162 9506
rect -106 9450 -38 9506
rect 18 9450 86 9506
rect 142 9450 210 9506
rect 266 9450 400 9506
rect -400 9382 400 9450
rect -400 9326 -286 9382
rect -230 9326 -162 9382
rect -106 9326 -38 9382
rect 18 9326 86 9382
rect 142 9326 210 9382
rect 266 9326 400 9382
rect -400 9258 400 9326
rect -400 9202 -286 9258
rect -230 9202 -162 9258
rect -106 9202 -38 9258
rect 18 9202 86 9258
rect 142 9202 210 9258
rect 266 9202 400 9258
rect -400 9134 400 9202
rect -400 9078 -286 9134
rect -230 9078 -162 9134
rect -106 9078 -38 9134
rect 18 9078 86 9134
rect 142 9078 210 9134
rect 266 9078 400 9134
rect -400 9010 400 9078
rect -400 8954 -286 9010
rect -230 8954 -162 9010
rect -106 8954 -38 9010
rect 18 8954 86 9010
rect 142 8954 210 9010
rect 266 8954 400 9010
rect -400 8886 400 8954
rect -400 8830 -286 8886
rect -230 8830 -162 8886
rect -106 8830 -38 8886
rect 18 8830 86 8886
rect 142 8830 210 8886
rect 266 8830 400 8886
rect -400 8762 400 8830
rect -400 8706 -286 8762
rect -230 8706 -162 8762
rect -106 8706 -38 8762
rect 18 8706 86 8762
rect 142 8706 210 8762
rect 266 8706 400 8762
rect -400 8638 400 8706
rect -400 8582 -286 8638
rect -230 8582 -162 8638
rect -106 8582 -38 8638
rect 18 8582 86 8638
rect 142 8582 210 8638
rect 266 8582 400 8638
rect -400 8514 400 8582
rect -400 8458 -286 8514
rect -230 8458 -162 8514
rect -106 8458 -38 8514
rect 18 8458 86 8514
rect 142 8458 210 8514
rect 266 8458 400 8514
rect -400 8390 400 8458
rect -400 8334 -286 8390
rect -230 8334 -162 8390
rect -106 8334 -38 8390
rect 18 8334 86 8390
rect 142 8334 210 8390
rect 266 8334 400 8390
rect -400 8266 400 8334
rect -400 8210 -286 8266
rect -230 8210 -162 8266
rect -106 8210 -38 8266
rect 18 8210 86 8266
rect 142 8210 210 8266
rect 266 8210 400 8266
rect -400 8142 400 8210
rect -400 8086 -286 8142
rect -230 8086 -162 8142
rect -106 8086 -38 8142
rect 18 8086 86 8142
rect 142 8086 210 8142
rect 266 8086 400 8142
rect -400 8018 400 8086
rect -400 7962 -286 8018
rect -230 7962 -162 8018
rect -106 7962 -38 8018
rect 18 7962 86 8018
rect 142 7962 210 8018
rect 266 7962 400 8018
rect -400 7894 400 7962
rect -400 7838 -286 7894
rect -230 7838 -162 7894
rect -106 7838 -38 7894
rect 18 7838 86 7894
rect 142 7838 210 7894
rect 266 7838 400 7894
rect -400 7770 400 7838
rect -400 7714 -286 7770
rect -230 7714 -162 7770
rect -106 7714 -38 7770
rect 18 7714 86 7770
rect 142 7714 210 7770
rect 266 7714 400 7770
rect -400 7646 400 7714
rect -400 7590 -286 7646
rect -230 7590 -162 7646
rect -106 7590 -38 7646
rect 18 7590 86 7646
rect 142 7590 210 7646
rect 266 7590 400 7646
rect -400 7522 400 7590
rect -400 7466 -286 7522
rect -230 7466 -162 7522
rect -106 7466 -38 7522
rect 18 7466 86 7522
rect 142 7466 210 7522
rect 266 7466 400 7522
rect -400 7398 400 7466
rect -400 7342 -286 7398
rect -230 7342 -162 7398
rect -106 7342 -38 7398
rect 18 7342 86 7398
rect 142 7342 210 7398
rect 266 7342 400 7398
rect -400 7274 400 7342
rect -400 7218 -286 7274
rect -230 7218 -162 7274
rect -106 7218 -38 7274
rect 18 7218 86 7274
rect 142 7218 210 7274
rect 266 7218 400 7274
rect -400 7150 400 7218
rect -400 7094 -286 7150
rect -230 7094 -162 7150
rect -106 7094 -38 7150
rect 18 7094 86 7150
rect 142 7094 210 7150
rect 266 7094 400 7150
rect -400 7026 400 7094
rect -400 6970 -286 7026
rect -230 6970 -162 7026
rect -106 6970 -38 7026
rect 18 6970 86 7026
rect 142 6970 210 7026
rect 266 6970 400 7026
rect -400 6902 400 6970
rect -400 6846 -286 6902
rect -230 6846 -162 6902
rect -106 6846 -38 6902
rect 18 6846 86 6902
rect 142 6846 210 6902
rect 266 6846 400 6902
rect -400 6778 400 6846
rect -400 6722 -286 6778
rect -230 6722 -162 6778
rect -106 6722 -38 6778
rect 18 6722 86 6778
rect 142 6722 210 6778
rect 266 6722 400 6778
rect -400 6654 400 6722
rect -400 6598 -286 6654
rect -230 6598 -162 6654
rect -106 6598 -38 6654
rect 18 6598 86 6654
rect 142 6598 210 6654
rect 266 6598 400 6654
rect -400 6530 400 6598
rect -400 6474 -286 6530
rect -230 6474 -162 6530
rect -106 6474 -38 6530
rect 18 6474 86 6530
rect 142 6474 210 6530
rect 266 6474 400 6530
rect -400 6406 400 6474
rect -400 6350 -286 6406
rect -230 6350 -162 6406
rect -106 6350 -38 6406
rect 18 6350 86 6406
rect 142 6350 210 6406
rect 266 6350 400 6406
rect -400 6282 400 6350
rect -400 6226 -286 6282
rect -230 6226 -162 6282
rect -106 6226 -38 6282
rect 18 6226 86 6282
rect 142 6226 210 6282
rect 266 6226 400 6282
rect -400 6158 400 6226
rect -400 6102 -286 6158
rect -230 6102 -162 6158
rect -106 6102 -38 6158
rect 18 6102 86 6158
rect 142 6102 210 6158
rect 266 6102 400 6158
rect -400 6034 400 6102
rect -400 5978 -286 6034
rect -230 5978 -162 6034
rect -106 5978 -38 6034
rect 18 5978 86 6034
rect 142 5978 210 6034
rect 266 5978 400 6034
rect -400 5910 400 5978
rect -400 5854 -286 5910
rect -230 5854 -162 5910
rect -106 5854 -38 5910
rect 18 5854 86 5910
rect 142 5854 210 5910
rect 266 5854 400 5910
rect -400 5786 400 5854
rect -400 5730 -286 5786
rect -230 5730 -162 5786
rect -106 5730 -38 5786
rect 18 5730 86 5786
rect 142 5730 210 5786
rect 266 5730 400 5786
rect -400 5662 400 5730
rect -400 5606 -286 5662
rect -230 5606 -162 5662
rect -106 5606 -38 5662
rect 18 5606 86 5662
rect 142 5606 210 5662
rect 266 5606 400 5662
rect -400 5538 400 5606
rect -400 5482 -286 5538
rect -230 5482 -162 5538
rect -106 5482 -38 5538
rect 18 5482 86 5538
rect 142 5482 210 5538
rect 266 5482 400 5538
rect -400 5414 400 5482
rect -400 5358 -286 5414
rect -230 5358 -162 5414
rect -106 5358 -38 5414
rect 18 5358 86 5414
rect 142 5358 210 5414
rect 266 5358 400 5414
rect -400 5290 400 5358
rect -400 5234 -286 5290
rect -230 5234 -162 5290
rect -106 5234 -38 5290
rect 18 5234 86 5290
rect 142 5234 210 5290
rect 266 5234 400 5290
rect -400 5166 400 5234
rect -400 5110 -286 5166
rect -230 5110 -162 5166
rect -106 5110 -38 5166
rect 18 5110 86 5166
rect 142 5110 210 5166
rect 266 5110 400 5166
rect -400 5042 400 5110
rect -400 4986 -286 5042
rect -230 4986 -162 5042
rect -106 4986 -38 5042
rect 18 4986 86 5042
rect 142 4986 210 5042
rect 266 4986 400 5042
rect -400 4918 400 4986
rect -400 4862 -286 4918
rect -230 4862 -162 4918
rect -106 4862 -38 4918
rect 18 4862 86 4918
rect 142 4862 210 4918
rect 266 4862 400 4918
rect -400 4794 400 4862
rect -400 4738 -286 4794
rect -230 4738 -162 4794
rect -106 4738 -38 4794
rect 18 4738 86 4794
rect 142 4738 210 4794
rect 266 4738 400 4794
rect -400 4670 400 4738
rect -400 4614 -286 4670
rect -230 4614 -162 4670
rect -106 4614 -38 4670
rect 18 4614 86 4670
rect 142 4614 210 4670
rect 266 4614 400 4670
rect -400 4546 400 4614
rect -400 4490 -286 4546
rect -230 4490 -162 4546
rect -106 4490 -38 4546
rect 18 4490 86 4546
rect 142 4490 210 4546
rect 266 4490 400 4546
rect -400 4422 400 4490
rect -400 4366 -286 4422
rect -230 4366 -162 4422
rect -106 4366 -38 4422
rect 18 4366 86 4422
rect 142 4366 210 4422
rect 266 4366 400 4422
rect -400 4298 400 4366
rect -400 4242 -286 4298
rect -230 4242 -162 4298
rect -106 4242 -38 4298
rect 18 4242 86 4298
rect 142 4242 210 4298
rect 266 4242 400 4298
rect -400 4174 400 4242
rect -400 4118 -286 4174
rect -230 4118 -162 4174
rect -106 4118 -38 4174
rect 18 4118 86 4174
rect 142 4118 210 4174
rect 266 4118 400 4174
rect -400 4050 400 4118
rect -400 3994 -286 4050
rect -230 3994 -162 4050
rect -106 3994 -38 4050
rect 18 3994 86 4050
rect 142 3994 210 4050
rect 266 3994 400 4050
rect -400 3926 400 3994
rect -400 3870 -286 3926
rect -230 3870 -162 3926
rect -106 3870 -38 3926
rect 18 3870 86 3926
rect 142 3870 210 3926
rect 266 3870 400 3926
rect -400 3802 400 3870
rect -400 3746 -286 3802
rect -230 3746 -162 3802
rect -106 3746 -38 3802
rect 18 3746 86 3802
rect 142 3746 210 3802
rect 266 3746 400 3802
rect -400 3678 400 3746
rect -400 3622 -286 3678
rect -230 3622 -162 3678
rect -106 3622 -38 3678
rect 18 3622 86 3678
rect 142 3622 210 3678
rect 266 3622 400 3678
rect -400 3554 400 3622
rect -400 3498 -286 3554
rect -230 3498 -162 3554
rect -106 3498 -38 3554
rect 18 3498 86 3554
rect 142 3498 210 3554
rect 266 3498 400 3554
rect -400 3430 400 3498
rect -400 3374 -286 3430
rect -230 3374 -162 3430
rect -106 3374 -38 3430
rect 18 3374 86 3430
rect 142 3374 210 3430
rect 266 3374 400 3430
rect -400 3306 400 3374
rect -400 3250 -286 3306
rect -230 3250 -162 3306
rect -106 3250 -38 3306
rect 18 3250 86 3306
rect 142 3250 210 3306
rect 266 3250 400 3306
rect -400 3182 400 3250
rect -400 3126 -286 3182
rect -230 3126 -162 3182
rect -106 3126 -38 3182
rect 18 3126 86 3182
rect 142 3126 210 3182
rect 266 3126 400 3182
rect -400 3058 400 3126
rect -400 3002 -286 3058
rect -230 3002 -162 3058
rect -106 3002 -38 3058
rect 18 3002 86 3058
rect 142 3002 210 3058
rect 266 3002 400 3058
rect -400 2934 400 3002
rect -400 2878 -286 2934
rect -230 2878 -162 2934
rect -106 2878 -38 2934
rect 18 2878 86 2934
rect 142 2878 210 2934
rect 266 2878 400 2934
rect -400 2810 400 2878
rect -400 2754 -286 2810
rect -230 2754 -162 2810
rect -106 2754 -38 2810
rect 18 2754 86 2810
rect 142 2754 210 2810
rect 266 2754 400 2810
rect -400 2686 400 2754
rect -400 2630 -286 2686
rect -230 2630 -162 2686
rect -106 2630 -38 2686
rect 18 2630 86 2686
rect 142 2630 210 2686
rect 266 2630 400 2686
rect -400 2562 400 2630
rect -400 2506 -286 2562
rect -230 2506 -162 2562
rect -106 2506 -38 2562
rect 18 2506 86 2562
rect 142 2506 210 2562
rect 266 2506 400 2562
rect -400 2438 400 2506
rect -400 2382 -286 2438
rect -230 2382 -162 2438
rect -106 2382 -38 2438
rect 18 2382 86 2438
rect 142 2382 210 2438
rect 266 2382 400 2438
rect -400 2314 400 2382
rect -400 2258 -286 2314
rect -230 2258 -162 2314
rect -106 2258 -38 2314
rect 18 2258 86 2314
rect 142 2258 210 2314
rect 266 2258 400 2314
rect -400 2190 400 2258
rect -400 2134 -286 2190
rect -230 2134 -162 2190
rect -106 2134 -38 2190
rect 18 2134 86 2190
rect 142 2134 210 2190
rect 266 2134 400 2190
rect -400 2066 400 2134
rect -400 2010 -286 2066
rect -230 2010 -162 2066
rect -106 2010 -38 2066
rect 18 2010 86 2066
rect 142 2010 210 2066
rect 266 2010 400 2066
rect -400 1942 400 2010
rect -400 1886 -286 1942
rect -230 1886 -162 1942
rect -106 1886 -38 1942
rect 18 1886 86 1942
rect 142 1886 210 1942
rect 266 1886 400 1942
rect -400 1818 400 1886
rect -400 1762 -286 1818
rect -230 1762 -162 1818
rect -106 1762 -38 1818
rect 18 1762 86 1818
rect 142 1762 210 1818
rect 266 1762 400 1818
rect -400 1694 400 1762
rect -400 1638 -286 1694
rect -230 1638 -162 1694
rect -106 1638 -38 1694
rect 18 1638 86 1694
rect 142 1638 210 1694
rect 266 1638 400 1694
rect -400 1570 400 1638
rect -400 1514 -286 1570
rect -230 1514 -162 1570
rect -106 1514 -38 1570
rect 18 1514 86 1570
rect 142 1514 210 1570
rect 266 1514 400 1570
rect -400 1446 400 1514
rect -400 1390 -286 1446
rect -230 1390 -162 1446
rect -106 1390 -38 1446
rect 18 1390 86 1446
rect 142 1390 210 1446
rect 266 1390 400 1446
rect -400 1322 400 1390
rect -400 1266 -286 1322
rect -230 1266 -162 1322
rect -106 1266 -38 1322
rect 18 1266 86 1322
rect 142 1266 210 1322
rect 266 1266 400 1322
rect -400 1198 400 1266
rect -400 1142 -286 1198
rect -230 1142 -162 1198
rect -106 1142 -38 1198
rect 18 1142 86 1198
rect 142 1142 210 1198
rect 266 1142 400 1198
rect -400 1074 400 1142
rect -400 1018 -286 1074
rect -230 1018 -162 1074
rect -106 1018 -38 1074
rect 18 1018 86 1074
rect 142 1018 210 1074
rect 266 1018 400 1074
rect -400 950 400 1018
rect -400 894 -286 950
rect -230 894 -162 950
rect -106 894 -38 950
rect 18 894 86 950
rect 142 894 210 950
rect 266 894 400 950
rect -400 826 400 894
rect -400 770 -286 826
rect -230 770 -162 826
rect -106 770 -38 826
rect 18 770 86 826
rect 142 770 210 826
rect 266 770 400 826
rect -400 702 400 770
rect -400 646 -286 702
rect -230 646 -162 702
rect -106 646 -38 702
rect 18 646 86 702
rect 142 646 210 702
rect 266 646 400 702
rect -400 578 400 646
rect -400 522 -286 578
rect -230 522 -162 578
rect -106 522 -38 578
rect 18 522 86 578
rect 142 522 210 578
rect 266 522 400 578
rect -400 458 400 522
rect 830 12310 1170 12320
rect 830 12254 903 12310
rect 959 12254 1045 12310
rect 1101 12254 1170 12310
rect 830 12168 1170 12254
rect 830 12112 903 12168
rect 959 12112 1045 12168
rect 1101 12112 1170 12168
rect 830 12026 1170 12112
rect 830 11970 903 12026
rect 959 11970 1045 12026
rect 1101 11970 1170 12026
rect 830 11884 1170 11970
rect 830 11828 903 11884
rect 959 11828 1045 11884
rect 1101 11828 1170 11884
rect 830 11742 1170 11828
rect 830 11686 903 11742
rect 959 11686 1045 11742
rect 1101 11686 1170 11742
rect 830 11600 1170 11686
rect 830 11544 903 11600
rect 959 11544 1045 11600
rect 1101 11544 1170 11600
rect 830 11458 1170 11544
rect 830 11402 903 11458
rect 959 11402 1045 11458
rect 1101 11402 1170 11458
rect 830 11316 1170 11402
rect 830 11260 903 11316
rect 959 11260 1045 11316
rect 1101 11260 1170 11316
rect 830 11174 1170 11260
rect 830 11118 903 11174
rect 959 11118 1045 11174
rect 1101 11118 1170 11174
rect 830 11032 1170 11118
rect 830 10976 903 11032
rect 959 10976 1045 11032
rect 1101 10976 1170 11032
rect 830 10890 1170 10976
rect 830 10834 903 10890
rect 959 10834 1045 10890
rect 1101 10834 1170 10890
rect 830 10748 1170 10834
rect 830 10692 903 10748
rect 959 10692 1045 10748
rect 1101 10692 1170 10748
rect 830 10606 1170 10692
rect 830 10550 903 10606
rect 959 10550 1045 10606
rect 1101 10550 1170 10606
rect 830 10464 1170 10550
rect 830 10408 903 10464
rect 959 10408 1045 10464
rect 1101 10408 1170 10464
rect 830 10322 1170 10408
rect 830 10266 903 10322
rect 959 10266 1045 10322
rect 1101 10266 1170 10322
rect 830 10180 1170 10266
rect 830 10124 903 10180
rect 959 10124 1045 10180
rect 1101 10124 1170 10180
rect 830 10038 1170 10124
rect 830 9982 903 10038
rect 959 9982 1045 10038
rect 1101 9982 1170 10038
rect 830 9896 1170 9982
rect 830 9840 903 9896
rect 959 9840 1045 9896
rect 1101 9840 1170 9896
rect 830 9754 1170 9840
rect 830 9698 903 9754
rect 959 9698 1045 9754
rect 1101 9698 1170 9754
rect 830 9612 1170 9698
rect 830 9556 903 9612
rect 959 9556 1045 9612
rect 1101 9556 1170 9612
rect 830 9470 1170 9556
rect 830 9414 903 9470
rect 959 9414 1045 9470
rect 1101 9414 1170 9470
rect 830 9328 1170 9414
rect 830 9272 903 9328
rect 959 9272 1045 9328
rect 1101 9272 1170 9328
rect 830 9186 1170 9272
rect 830 9130 903 9186
rect 959 9130 1045 9186
rect 1101 9130 1170 9186
rect 830 9044 1170 9130
rect 830 8988 903 9044
rect 959 8988 1045 9044
rect 1101 8988 1170 9044
rect 830 8902 1170 8988
rect 830 8846 903 8902
rect 959 8846 1045 8902
rect 1101 8846 1170 8902
rect 830 8760 1170 8846
rect 830 8704 903 8760
rect 959 8704 1045 8760
rect 1101 8704 1170 8760
rect 830 8618 1170 8704
rect 830 8562 903 8618
rect 959 8562 1045 8618
rect 1101 8562 1170 8618
rect 830 8476 1170 8562
rect 830 8420 903 8476
rect 959 8420 1045 8476
rect 1101 8420 1170 8476
rect 830 8334 1170 8420
rect 830 8278 903 8334
rect 959 8278 1045 8334
rect 1101 8278 1170 8334
rect 830 8192 1170 8278
rect 830 8136 903 8192
rect 959 8136 1045 8192
rect 1101 8136 1170 8192
rect 830 8050 1170 8136
rect 830 7994 903 8050
rect 959 7994 1045 8050
rect 1101 7994 1170 8050
rect 830 7908 1170 7994
rect 830 7852 903 7908
rect 959 7852 1045 7908
rect 1101 7852 1170 7908
rect 830 7766 1170 7852
rect 830 7710 903 7766
rect 959 7710 1045 7766
rect 1101 7710 1170 7766
rect 830 7624 1170 7710
rect 830 7568 903 7624
rect 959 7568 1045 7624
rect 1101 7568 1170 7624
rect 830 7482 1170 7568
rect 830 7426 903 7482
rect 959 7426 1045 7482
rect 1101 7426 1170 7482
rect 830 7340 1170 7426
rect 830 7284 903 7340
rect 959 7284 1045 7340
rect 1101 7284 1170 7340
rect 830 7198 1170 7284
rect 830 7142 903 7198
rect 959 7142 1045 7198
rect 1101 7142 1170 7198
rect 830 7056 1170 7142
rect 830 7000 903 7056
rect 959 7000 1045 7056
rect 1101 7000 1170 7056
rect 830 6914 1170 7000
rect 830 6858 903 6914
rect 959 6858 1045 6914
rect 1101 6858 1170 6914
rect 830 6772 1170 6858
rect 830 6716 903 6772
rect 959 6716 1045 6772
rect 1101 6716 1170 6772
rect 830 6630 1170 6716
rect 830 6574 903 6630
rect 959 6574 1045 6630
rect 1101 6574 1170 6630
rect 830 6488 1170 6574
rect 830 6432 903 6488
rect 959 6432 1045 6488
rect 1101 6432 1170 6488
rect 830 6346 1170 6432
rect 830 6290 903 6346
rect 959 6290 1045 6346
rect 1101 6290 1170 6346
rect 830 6204 1170 6290
rect 830 6148 903 6204
rect 959 6148 1045 6204
rect 1101 6148 1170 6204
rect 830 6062 1170 6148
rect 830 6006 903 6062
rect 959 6006 1045 6062
rect 1101 6006 1170 6062
rect 830 5920 1170 6006
rect 830 5864 903 5920
rect 959 5864 1045 5920
rect 1101 5864 1170 5920
rect 830 5778 1170 5864
rect 830 5722 903 5778
rect 959 5722 1045 5778
rect 1101 5722 1170 5778
rect 830 5636 1170 5722
rect 830 5580 903 5636
rect 959 5580 1045 5636
rect 1101 5580 1170 5636
rect 830 5494 1170 5580
rect 830 5438 903 5494
rect 959 5438 1045 5494
rect 1101 5438 1170 5494
rect 830 5352 1170 5438
rect 830 5296 903 5352
rect 959 5296 1045 5352
rect 1101 5296 1170 5352
rect 830 5210 1170 5296
rect 830 5154 903 5210
rect 959 5154 1045 5210
rect 1101 5154 1170 5210
rect 830 5068 1170 5154
rect 830 5012 903 5068
rect 959 5012 1045 5068
rect 1101 5012 1170 5068
rect 830 4926 1170 5012
rect 830 4870 903 4926
rect 959 4870 1045 4926
rect 1101 4870 1170 4926
rect 830 4784 1170 4870
rect 830 4728 903 4784
rect 959 4728 1045 4784
rect 1101 4728 1170 4784
rect 830 4642 1170 4728
rect 830 4586 903 4642
rect 959 4586 1045 4642
rect 1101 4586 1170 4642
rect 830 4500 1170 4586
rect 830 4444 903 4500
rect 959 4444 1045 4500
rect 1101 4444 1170 4500
rect 830 4358 1170 4444
rect 830 4302 903 4358
rect 959 4302 1045 4358
rect 1101 4302 1170 4358
rect 830 4216 1170 4302
rect 830 4160 903 4216
rect 959 4160 1045 4216
rect 1101 4160 1170 4216
rect 830 4074 1170 4160
rect 830 4018 903 4074
rect 959 4018 1045 4074
rect 1101 4018 1170 4074
rect 830 3932 1170 4018
rect 830 3876 903 3932
rect 959 3876 1045 3932
rect 1101 3876 1170 3932
rect 830 3790 1170 3876
rect 830 3734 903 3790
rect 959 3734 1045 3790
rect 1101 3734 1170 3790
rect 830 3648 1170 3734
rect 830 3592 903 3648
rect 959 3592 1045 3648
rect 1101 3592 1170 3648
rect 830 3506 1170 3592
rect 830 3450 903 3506
rect 959 3450 1045 3506
rect 1101 3450 1170 3506
rect 830 3364 1170 3450
rect 830 3308 903 3364
rect 959 3308 1045 3364
rect 1101 3308 1170 3364
rect 830 3222 1170 3308
rect 830 3166 903 3222
rect 959 3166 1045 3222
rect 1101 3166 1170 3222
rect 830 3080 1170 3166
rect 830 3024 903 3080
rect 959 3024 1045 3080
rect 1101 3024 1170 3080
rect 830 2938 1170 3024
rect 830 2882 903 2938
rect 959 2882 1045 2938
rect 1101 2882 1170 2938
rect 830 2796 1170 2882
rect 830 2740 903 2796
rect 959 2740 1045 2796
rect 1101 2740 1170 2796
rect 830 2654 1170 2740
rect 830 2598 903 2654
rect 959 2598 1045 2654
rect 1101 2598 1170 2654
rect 830 2512 1170 2598
rect 830 2456 903 2512
rect 959 2456 1045 2512
rect 1101 2456 1170 2512
rect 830 2370 1170 2456
rect 830 2314 903 2370
rect 959 2314 1045 2370
rect 1101 2314 1170 2370
rect 830 2228 1170 2314
rect 830 2172 903 2228
rect 959 2172 1045 2228
rect 1101 2172 1170 2228
rect 830 2086 1170 2172
rect 830 2030 903 2086
rect 959 2030 1045 2086
rect 1101 2030 1170 2086
rect 830 1944 1170 2030
rect 830 1888 903 1944
rect 959 1888 1045 1944
rect 1101 1888 1170 1944
rect 830 1802 1170 1888
rect 830 1746 903 1802
rect 959 1746 1045 1802
rect 1101 1746 1170 1802
rect 830 1660 1170 1746
rect 830 1604 903 1660
rect 959 1604 1045 1660
rect 1101 1604 1170 1660
rect 830 1518 1170 1604
rect 830 1462 903 1518
rect 959 1462 1045 1518
rect 1101 1462 1170 1518
rect 830 1376 1170 1462
rect 830 1320 903 1376
rect 959 1320 1045 1376
rect 1101 1320 1170 1376
rect 830 1234 1170 1320
rect 830 1178 903 1234
rect 959 1178 1045 1234
rect 1101 1178 1170 1234
rect 830 1092 1170 1178
rect 830 1036 903 1092
rect 959 1036 1045 1092
rect 1101 1036 1170 1092
rect 830 950 1170 1036
rect 830 894 903 950
rect 959 894 1045 950
rect 1101 894 1170 950
rect 830 808 1170 894
rect 830 752 903 808
rect 959 752 1045 808
rect 1101 752 1170 808
rect 830 666 1170 752
rect 830 610 903 666
rect 959 610 1045 666
rect 1101 610 1170 666
rect 830 524 1170 610
rect 830 468 903 524
rect 959 468 1045 524
rect 1101 468 1170 524
rect 830 458 1170 468
rect 1370 12310 1710 12320
rect 1370 12254 1444 12310
rect 1500 12254 1586 12310
rect 1642 12254 1710 12310
rect 1370 12168 1710 12254
rect 1370 12112 1444 12168
rect 1500 12112 1586 12168
rect 1642 12112 1710 12168
rect 1370 12026 1710 12112
rect 1370 11970 1444 12026
rect 1500 11970 1586 12026
rect 1642 11970 1710 12026
rect 1370 11884 1710 11970
rect 1370 11828 1444 11884
rect 1500 11828 1586 11884
rect 1642 11828 1710 11884
rect 1370 11742 1710 11828
rect 1370 11686 1444 11742
rect 1500 11686 1586 11742
rect 1642 11686 1710 11742
rect 1370 11600 1710 11686
rect 1370 11544 1444 11600
rect 1500 11544 1586 11600
rect 1642 11544 1710 11600
rect 1370 11458 1710 11544
rect 1370 11402 1444 11458
rect 1500 11402 1586 11458
rect 1642 11402 1710 11458
rect 1370 11316 1710 11402
rect 1370 11260 1444 11316
rect 1500 11260 1586 11316
rect 1642 11260 1710 11316
rect 1370 11174 1710 11260
rect 1370 11118 1444 11174
rect 1500 11118 1586 11174
rect 1642 11118 1710 11174
rect 1370 11032 1710 11118
rect 1370 10976 1444 11032
rect 1500 10976 1586 11032
rect 1642 10976 1710 11032
rect 1370 10890 1710 10976
rect 1370 10834 1444 10890
rect 1500 10834 1586 10890
rect 1642 10834 1710 10890
rect 1370 10748 1710 10834
rect 1370 10692 1444 10748
rect 1500 10692 1586 10748
rect 1642 10692 1710 10748
rect 1370 10606 1710 10692
rect 1370 10550 1444 10606
rect 1500 10550 1586 10606
rect 1642 10550 1710 10606
rect 1370 10464 1710 10550
rect 1370 10408 1444 10464
rect 1500 10408 1586 10464
rect 1642 10408 1710 10464
rect 1370 10322 1710 10408
rect 1370 10266 1444 10322
rect 1500 10266 1586 10322
rect 1642 10266 1710 10322
rect 1370 10180 1710 10266
rect 1370 10124 1444 10180
rect 1500 10124 1586 10180
rect 1642 10124 1710 10180
rect 1370 10038 1710 10124
rect 1370 9982 1444 10038
rect 1500 9982 1586 10038
rect 1642 9982 1710 10038
rect 1370 9896 1710 9982
rect 1370 9840 1444 9896
rect 1500 9840 1586 9896
rect 1642 9840 1710 9896
rect 1370 9754 1710 9840
rect 1370 9698 1444 9754
rect 1500 9698 1586 9754
rect 1642 9698 1710 9754
rect 1370 9612 1710 9698
rect 1370 9556 1444 9612
rect 1500 9556 1586 9612
rect 1642 9556 1710 9612
rect 1370 9470 1710 9556
rect 1370 9414 1444 9470
rect 1500 9414 1586 9470
rect 1642 9414 1710 9470
rect 1370 9328 1710 9414
rect 1370 9272 1444 9328
rect 1500 9272 1586 9328
rect 1642 9272 1710 9328
rect 1370 9186 1710 9272
rect 1370 9130 1444 9186
rect 1500 9130 1586 9186
rect 1642 9130 1710 9186
rect 1370 9044 1710 9130
rect 1370 8988 1444 9044
rect 1500 8988 1586 9044
rect 1642 8988 1710 9044
rect 1370 8902 1710 8988
rect 1370 8846 1444 8902
rect 1500 8846 1586 8902
rect 1642 8846 1710 8902
rect 1370 8760 1710 8846
rect 1370 8704 1444 8760
rect 1500 8704 1586 8760
rect 1642 8704 1710 8760
rect 1370 8618 1710 8704
rect 1370 8562 1444 8618
rect 1500 8562 1586 8618
rect 1642 8562 1710 8618
rect 1370 8476 1710 8562
rect 1370 8420 1444 8476
rect 1500 8420 1586 8476
rect 1642 8420 1710 8476
rect 1370 8334 1710 8420
rect 1370 8278 1444 8334
rect 1500 8278 1586 8334
rect 1642 8278 1710 8334
rect 1370 8192 1710 8278
rect 1370 8136 1444 8192
rect 1500 8136 1586 8192
rect 1642 8136 1710 8192
rect 1370 8050 1710 8136
rect 1370 7994 1444 8050
rect 1500 7994 1586 8050
rect 1642 7994 1710 8050
rect 1370 7908 1710 7994
rect 1370 7852 1444 7908
rect 1500 7852 1586 7908
rect 1642 7852 1710 7908
rect 1370 7766 1710 7852
rect 1370 7710 1444 7766
rect 1500 7710 1586 7766
rect 1642 7710 1710 7766
rect 1370 7624 1710 7710
rect 1370 7568 1444 7624
rect 1500 7568 1586 7624
rect 1642 7568 1710 7624
rect 1370 7482 1710 7568
rect 1370 7426 1444 7482
rect 1500 7426 1586 7482
rect 1642 7426 1710 7482
rect 1370 7340 1710 7426
rect 1370 7284 1444 7340
rect 1500 7284 1586 7340
rect 1642 7284 1710 7340
rect 1370 7198 1710 7284
rect 1370 7142 1444 7198
rect 1500 7142 1586 7198
rect 1642 7142 1710 7198
rect 1370 7056 1710 7142
rect 1370 7000 1444 7056
rect 1500 7000 1586 7056
rect 1642 7000 1710 7056
rect 1370 6914 1710 7000
rect 1370 6858 1444 6914
rect 1500 6858 1586 6914
rect 1642 6858 1710 6914
rect 1370 6772 1710 6858
rect 1370 6716 1444 6772
rect 1500 6716 1586 6772
rect 1642 6716 1710 6772
rect 1370 6630 1710 6716
rect 1370 6574 1444 6630
rect 1500 6574 1586 6630
rect 1642 6574 1710 6630
rect 1370 6488 1710 6574
rect 1370 6432 1444 6488
rect 1500 6432 1586 6488
rect 1642 6432 1710 6488
rect 1370 6346 1710 6432
rect 1370 6290 1444 6346
rect 1500 6290 1586 6346
rect 1642 6290 1710 6346
rect 1370 6204 1710 6290
rect 1370 6148 1444 6204
rect 1500 6148 1586 6204
rect 1642 6148 1710 6204
rect 1370 6062 1710 6148
rect 1370 6006 1444 6062
rect 1500 6006 1586 6062
rect 1642 6006 1710 6062
rect 1370 5920 1710 6006
rect 1370 5864 1444 5920
rect 1500 5864 1586 5920
rect 1642 5864 1710 5920
rect 1370 5778 1710 5864
rect 1370 5722 1444 5778
rect 1500 5722 1586 5778
rect 1642 5722 1710 5778
rect 1370 5636 1710 5722
rect 1370 5580 1444 5636
rect 1500 5580 1586 5636
rect 1642 5580 1710 5636
rect 1370 5494 1710 5580
rect 1370 5438 1444 5494
rect 1500 5438 1586 5494
rect 1642 5438 1710 5494
rect 1370 5352 1710 5438
rect 1370 5296 1444 5352
rect 1500 5296 1586 5352
rect 1642 5296 1710 5352
rect 1370 5210 1710 5296
rect 1370 5154 1444 5210
rect 1500 5154 1586 5210
rect 1642 5154 1710 5210
rect 1370 5068 1710 5154
rect 1370 5012 1444 5068
rect 1500 5012 1586 5068
rect 1642 5012 1710 5068
rect 1370 4926 1710 5012
rect 1370 4870 1444 4926
rect 1500 4870 1586 4926
rect 1642 4870 1710 4926
rect 1370 4784 1710 4870
rect 1370 4728 1444 4784
rect 1500 4728 1586 4784
rect 1642 4728 1710 4784
rect 1370 4642 1710 4728
rect 1370 4586 1444 4642
rect 1500 4586 1586 4642
rect 1642 4586 1710 4642
rect 1370 4500 1710 4586
rect 1370 4444 1444 4500
rect 1500 4444 1586 4500
rect 1642 4444 1710 4500
rect 1370 4358 1710 4444
rect 1370 4302 1444 4358
rect 1500 4302 1586 4358
rect 1642 4302 1710 4358
rect 1370 4216 1710 4302
rect 1370 4160 1444 4216
rect 1500 4160 1586 4216
rect 1642 4160 1710 4216
rect 1370 4074 1710 4160
rect 1370 4018 1444 4074
rect 1500 4018 1586 4074
rect 1642 4018 1710 4074
rect 1370 3932 1710 4018
rect 1370 3876 1444 3932
rect 1500 3876 1586 3932
rect 1642 3876 1710 3932
rect 1370 3790 1710 3876
rect 1370 3734 1444 3790
rect 1500 3734 1586 3790
rect 1642 3734 1710 3790
rect 1370 3648 1710 3734
rect 1370 3592 1444 3648
rect 1500 3592 1586 3648
rect 1642 3592 1710 3648
rect 1370 3506 1710 3592
rect 1370 3450 1444 3506
rect 1500 3450 1586 3506
rect 1642 3450 1710 3506
rect 1370 3364 1710 3450
rect 1370 3308 1444 3364
rect 1500 3308 1586 3364
rect 1642 3308 1710 3364
rect 1370 3222 1710 3308
rect 1370 3166 1444 3222
rect 1500 3166 1586 3222
rect 1642 3166 1710 3222
rect 1370 3080 1710 3166
rect 1370 3024 1444 3080
rect 1500 3024 1586 3080
rect 1642 3024 1710 3080
rect 1370 2938 1710 3024
rect 1370 2882 1444 2938
rect 1500 2882 1586 2938
rect 1642 2882 1710 2938
rect 1370 2796 1710 2882
rect 1370 2740 1444 2796
rect 1500 2740 1586 2796
rect 1642 2740 1710 2796
rect 1370 2654 1710 2740
rect 1370 2598 1444 2654
rect 1500 2598 1586 2654
rect 1642 2598 1710 2654
rect 1370 2512 1710 2598
rect 1370 2456 1444 2512
rect 1500 2456 1586 2512
rect 1642 2456 1710 2512
rect 1370 2370 1710 2456
rect 1370 2314 1444 2370
rect 1500 2314 1586 2370
rect 1642 2314 1710 2370
rect 1370 2228 1710 2314
rect 1370 2172 1444 2228
rect 1500 2172 1586 2228
rect 1642 2172 1710 2228
rect 1370 2086 1710 2172
rect 1370 2030 1444 2086
rect 1500 2030 1586 2086
rect 1642 2030 1710 2086
rect 1370 1944 1710 2030
rect 1370 1888 1444 1944
rect 1500 1888 1586 1944
rect 1642 1888 1710 1944
rect 1370 1802 1710 1888
rect 1370 1746 1444 1802
rect 1500 1746 1586 1802
rect 1642 1746 1710 1802
rect 1370 1660 1710 1746
rect 1370 1604 1444 1660
rect 1500 1604 1586 1660
rect 1642 1604 1710 1660
rect 1370 1518 1710 1604
rect 1370 1462 1444 1518
rect 1500 1462 1586 1518
rect 1642 1462 1710 1518
rect 1370 1376 1710 1462
rect 1370 1320 1444 1376
rect 1500 1320 1586 1376
rect 1642 1320 1710 1376
rect 1370 1234 1710 1320
rect 1370 1178 1444 1234
rect 1500 1178 1586 1234
rect 1642 1178 1710 1234
rect 1370 1092 1710 1178
rect 1370 1036 1444 1092
rect 1500 1036 1586 1092
rect 1642 1036 1710 1092
rect 1370 950 1710 1036
rect 1370 894 1444 950
rect 1500 894 1586 950
rect 1642 894 1710 950
rect 1370 808 1710 894
rect 1370 752 1444 808
rect 1500 752 1586 808
rect 1642 752 1710 808
rect 1370 666 1710 752
rect 1370 610 1444 666
rect 1500 610 1586 666
rect 1642 610 1710 666
rect 1370 524 1710 610
rect 1370 468 1444 524
rect 1500 468 1586 524
rect 1642 468 1710 524
rect 1370 458 1710 468
rect 1910 12310 2250 12320
rect 1910 12254 1984 12310
rect 2040 12254 2126 12310
rect 2182 12254 2250 12310
rect 1910 12168 2250 12254
rect 1910 12112 1984 12168
rect 2040 12112 2126 12168
rect 2182 12112 2250 12168
rect 1910 12026 2250 12112
rect 1910 11970 1984 12026
rect 2040 11970 2126 12026
rect 2182 11970 2250 12026
rect 1910 11884 2250 11970
rect 1910 11828 1984 11884
rect 2040 11828 2126 11884
rect 2182 11828 2250 11884
rect 1910 11742 2250 11828
rect 1910 11686 1984 11742
rect 2040 11686 2126 11742
rect 2182 11686 2250 11742
rect 1910 11600 2250 11686
rect 1910 11544 1984 11600
rect 2040 11544 2126 11600
rect 2182 11544 2250 11600
rect 1910 11458 2250 11544
rect 1910 11402 1984 11458
rect 2040 11402 2126 11458
rect 2182 11402 2250 11458
rect 1910 11316 2250 11402
rect 1910 11260 1984 11316
rect 2040 11260 2126 11316
rect 2182 11260 2250 11316
rect 1910 11174 2250 11260
rect 1910 11118 1984 11174
rect 2040 11118 2126 11174
rect 2182 11118 2250 11174
rect 1910 11032 2250 11118
rect 1910 10976 1984 11032
rect 2040 10976 2126 11032
rect 2182 10976 2250 11032
rect 1910 10890 2250 10976
rect 1910 10834 1984 10890
rect 2040 10834 2126 10890
rect 2182 10834 2250 10890
rect 1910 10748 2250 10834
rect 1910 10692 1984 10748
rect 2040 10692 2126 10748
rect 2182 10692 2250 10748
rect 1910 10606 2250 10692
rect 1910 10550 1984 10606
rect 2040 10550 2126 10606
rect 2182 10550 2250 10606
rect 1910 10464 2250 10550
rect 1910 10408 1984 10464
rect 2040 10408 2126 10464
rect 2182 10408 2250 10464
rect 1910 10322 2250 10408
rect 1910 10266 1984 10322
rect 2040 10266 2126 10322
rect 2182 10266 2250 10322
rect 1910 10180 2250 10266
rect 1910 10124 1984 10180
rect 2040 10124 2126 10180
rect 2182 10124 2250 10180
rect 1910 10038 2250 10124
rect 1910 9982 1984 10038
rect 2040 9982 2126 10038
rect 2182 9982 2250 10038
rect 1910 9896 2250 9982
rect 1910 9840 1984 9896
rect 2040 9840 2126 9896
rect 2182 9840 2250 9896
rect 1910 9754 2250 9840
rect 1910 9698 1984 9754
rect 2040 9698 2126 9754
rect 2182 9698 2250 9754
rect 1910 9612 2250 9698
rect 1910 9556 1984 9612
rect 2040 9556 2126 9612
rect 2182 9556 2250 9612
rect 1910 9470 2250 9556
rect 1910 9414 1984 9470
rect 2040 9414 2126 9470
rect 2182 9414 2250 9470
rect 1910 9328 2250 9414
rect 1910 9272 1984 9328
rect 2040 9272 2126 9328
rect 2182 9272 2250 9328
rect 1910 9186 2250 9272
rect 1910 9130 1984 9186
rect 2040 9130 2126 9186
rect 2182 9130 2250 9186
rect 1910 9044 2250 9130
rect 1910 8988 1984 9044
rect 2040 8988 2126 9044
rect 2182 8988 2250 9044
rect 1910 8902 2250 8988
rect 1910 8846 1984 8902
rect 2040 8846 2126 8902
rect 2182 8846 2250 8902
rect 1910 8760 2250 8846
rect 1910 8704 1984 8760
rect 2040 8704 2126 8760
rect 2182 8704 2250 8760
rect 1910 8618 2250 8704
rect 1910 8562 1984 8618
rect 2040 8562 2126 8618
rect 2182 8562 2250 8618
rect 1910 8476 2250 8562
rect 1910 8420 1984 8476
rect 2040 8420 2126 8476
rect 2182 8420 2250 8476
rect 1910 8334 2250 8420
rect 1910 8278 1984 8334
rect 2040 8278 2126 8334
rect 2182 8278 2250 8334
rect 1910 8192 2250 8278
rect 1910 8136 1984 8192
rect 2040 8136 2126 8192
rect 2182 8136 2250 8192
rect 1910 8050 2250 8136
rect 1910 7994 1984 8050
rect 2040 7994 2126 8050
rect 2182 7994 2250 8050
rect 1910 7908 2250 7994
rect 1910 7852 1984 7908
rect 2040 7852 2126 7908
rect 2182 7852 2250 7908
rect 1910 7766 2250 7852
rect 1910 7710 1984 7766
rect 2040 7710 2126 7766
rect 2182 7710 2250 7766
rect 1910 7624 2250 7710
rect 1910 7568 1984 7624
rect 2040 7568 2126 7624
rect 2182 7568 2250 7624
rect 1910 7482 2250 7568
rect 1910 7426 1984 7482
rect 2040 7426 2126 7482
rect 2182 7426 2250 7482
rect 1910 7340 2250 7426
rect 1910 7284 1984 7340
rect 2040 7284 2126 7340
rect 2182 7284 2250 7340
rect 1910 7198 2250 7284
rect 1910 7142 1984 7198
rect 2040 7142 2126 7198
rect 2182 7142 2250 7198
rect 1910 7056 2250 7142
rect 1910 7000 1984 7056
rect 2040 7000 2126 7056
rect 2182 7000 2250 7056
rect 1910 6914 2250 7000
rect 1910 6858 1984 6914
rect 2040 6858 2126 6914
rect 2182 6858 2250 6914
rect 1910 6772 2250 6858
rect 1910 6716 1984 6772
rect 2040 6716 2126 6772
rect 2182 6716 2250 6772
rect 1910 6630 2250 6716
rect 1910 6574 1984 6630
rect 2040 6574 2126 6630
rect 2182 6574 2250 6630
rect 1910 6488 2250 6574
rect 1910 6432 1984 6488
rect 2040 6432 2126 6488
rect 2182 6432 2250 6488
rect 1910 6346 2250 6432
rect 1910 6290 1984 6346
rect 2040 6290 2126 6346
rect 2182 6290 2250 6346
rect 1910 6204 2250 6290
rect 1910 6148 1984 6204
rect 2040 6148 2126 6204
rect 2182 6148 2250 6204
rect 1910 6062 2250 6148
rect 1910 6006 1984 6062
rect 2040 6006 2126 6062
rect 2182 6006 2250 6062
rect 1910 5920 2250 6006
rect 1910 5864 1984 5920
rect 2040 5864 2126 5920
rect 2182 5864 2250 5920
rect 1910 5778 2250 5864
rect 1910 5722 1984 5778
rect 2040 5722 2126 5778
rect 2182 5722 2250 5778
rect 1910 5636 2250 5722
rect 1910 5580 1984 5636
rect 2040 5580 2126 5636
rect 2182 5580 2250 5636
rect 1910 5494 2250 5580
rect 1910 5438 1984 5494
rect 2040 5438 2126 5494
rect 2182 5438 2250 5494
rect 1910 5352 2250 5438
rect 1910 5296 1984 5352
rect 2040 5296 2126 5352
rect 2182 5296 2250 5352
rect 1910 5210 2250 5296
rect 1910 5154 1984 5210
rect 2040 5154 2126 5210
rect 2182 5154 2250 5210
rect 1910 5068 2250 5154
rect 1910 5012 1984 5068
rect 2040 5012 2126 5068
rect 2182 5012 2250 5068
rect 1910 4926 2250 5012
rect 1910 4870 1984 4926
rect 2040 4870 2126 4926
rect 2182 4870 2250 4926
rect 1910 4784 2250 4870
rect 1910 4728 1984 4784
rect 2040 4728 2126 4784
rect 2182 4728 2250 4784
rect 1910 4642 2250 4728
rect 1910 4586 1984 4642
rect 2040 4586 2126 4642
rect 2182 4586 2250 4642
rect 1910 4500 2250 4586
rect 1910 4444 1984 4500
rect 2040 4444 2126 4500
rect 2182 4444 2250 4500
rect 1910 4358 2250 4444
rect 1910 4302 1984 4358
rect 2040 4302 2126 4358
rect 2182 4302 2250 4358
rect 1910 4216 2250 4302
rect 1910 4160 1984 4216
rect 2040 4160 2126 4216
rect 2182 4160 2250 4216
rect 1910 4074 2250 4160
rect 1910 4018 1984 4074
rect 2040 4018 2126 4074
rect 2182 4018 2250 4074
rect 1910 3932 2250 4018
rect 1910 3876 1984 3932
rect 2040 3876 2126 3932
rect 2182 3876 2250 3932
rect 1910 3790 2250 3876
rect 1910 3734 1984 3790
rect 2040 3734 2126 3790
rect 2182 3734 2250 3790
rect 1910 3648 2250 3734
rect 1910 3592 1984 3648
rect 2040 3592 2126 3648
rect 2182 3592 2250 3648
rect 1910 3506 2250 3592
rect 1910 3450 1984 3506
rect 2040 3450 2126 3506
rect 2182 3450 2250 3506
rect 1910 3364 2250 3450
rect 1910 3308 1984 3364
rect 2040 3308 2126 3364
rect 2182 3308 2250 3364
rect 1910 3222 2250 3308
rect 1910 3166 1984 3222
rect 2040 3166 2126 3222
rect 2182 3166 2250 3222
rect 1910 3080 2250 3166
rect 1910 3024 1984 3080
rect 2040 3024 2126 3080
rect 2182 3024 2250 3080
rect 1910 2938 2250 3024
rect 1910 2882 1984 2938
rect 2040 2882 2126 2938
rect 2182 2882 2250 2938
rect 1910 2796 2250 2882
rect 1910 2740 1984 2796
rect 2040 2740 2126 2796
rect 2182 2740 2250 2796
rect 1910 2654 2250 2740
rect 1910 2598 1984 2654
rect 2040 2598 2126 2654
rect 2182 2598 2250 2654
rect 1910 2512 2250 2598
rect 1910 2456 1984 2512
rect 2040 2456 2126 2512
rect 2182 2456 2250 2512
rect 1910 2370 2250 2456
rect 1910 2314 1984 2370
rect 2040 2314 2126 2370
rect 2182 2314 2250 2370
rect 1910 2228 2250 2314
rect 1910 2172 1984 2228
rect 2040 2172 2126 2228
rect 2182 2172 2250 2228
rect 1910 2086 2250 2172
rect 1910 2030 1984 2086
rect 2040 2030 2126 2086
rect 2182 2030 2250 2086
rect 1910 1944 2250 2030
rect 1910 1888 1984 1944
rect 2040 1888 2126 1944
rect 2182 1888 2250 1944
rect 1910 1802 2250 1888
rect 1910 1746 1984 1802
rect 2040 1746 2126 1802
rect 2182 1746 2250 1802
rect 1910 1660 2250 1746
rect 1910 1604 1984 1660
rect 2040 1604 2126 1660
rect 2182 1604 2250 1660
rect 1910 1518 2250 1604
rect 1910 1462 1984 1518
rect 2040 1462 2126 1518
rect 2182 1462 2250 1518
rect 1910 1376 2250 1462
rect 1910 1320 1984 1376
rect 2040 1320 2126 1376
rect 2182 1320 2250 1376
rect 1910 1234 2250 1320
rect 1910 1178 1984 1234
rect 2040 1178 2126 1234
rect 2182 1178 2250 1234
rect 1910 1092 2250 1178
rect 1910 1036 1984 1092
rect 2040 1036 2126 1092
rect 2182 1036 2250 1092
rect 1910 950 2250 1036
rect 1910 894 1984 950
rect 2040 894 2126 950
rect 2182 894 2250 950
rect 1910 808 2250 894
rect 1910 752 1984 808
rect 2040 752 2126 808
rect 2182 752 2250 808
rect 1910 666 2250 752
rect 1910 610 1984 666
rect 2040 610 2126 666
rect 2182 610 2250 666
rect 1910 524 2250 610
rect 1910 468 1984 524
rect 2040 468 2126 524
rect 2182 468 2250 524
rect 1910 458 2250 468
rect 2450 12310 2790 12320
rect 2450 12254 2521 12310
rect 2577 12254 2663 12310
rect 2719 12254 2790 12310
rect 2450 12168 2790 12254
rect 2450 12112 2521 12168
rect 2577 12112 2663 12168
rect 2719 12112 2790 12168
rect 2450 12026 2790 12112
rect 2450 11970 2521 12026
rect 2577 11970 2663 12026
rect 2719 11970 2790 12026
rect 2450 11884 2790 11970
rect 2450 11828 2521 11884
rect 2577 11828 2663 11884
rect 2719 11828 2790 11884
rect 2450 11742 2790 11828
rect 2450 11686 2521 11742
rect 2577 11686 2663 11742
rect 2719 11686 2790 11742
rect 2450 11600 2790 11686
rect 2450 11544 2521 11600
rect 2577 11544 2663 11600
rect 2719 11544 2790 11600
rect 2450 11458 2790 11544
rect 2450 11402 2521 11458
rect 2577 11402 2663 11458
rect 2719 11402 2790 11458
rect 2450 11316 2790 11402
rect 2450 11260 2521 11316
rect 2577 11260 2663 11316
rect 2719 11260 2790 11316
rect 2450 11174 2790 11260
rect 2450 11118 2521 11174
rect 2577 11118 2663 11174
rect 2719 11118 2790 11174
rect 2450 11032 2790 11118
rect 2450 10976 2521 11032
rect 2577 10976 2663 11032
rect 2719 10976 2790 11032
rect 2450 10890 2790 10976
rect 2450 10834 2521 10890
rect 2577 10834 2663 10890
rect 2719 10834 2790 10890
rect 2450 10748 2790 10834
rect 2450 10692 2521 10748
rect 2577 10692 2663 10748
rect 2719 10692 2790 10748
rect 2450 10606 2790 10692
rect 2450 10550 2521 10606
rect 2577 10550 2663 10606
rect 2719 10550 2790 10606
rect 2450 10464 2790 10550
rect 2450 10408 2521 10464
rect 2577 10408 2663 10464
rect 2719 10408 2790 10464
rect 2450 10322 2790 10408
rect 2450 10266 2521 10322
rect 2577 10266 2663 10322
rect 2719 10266 2790 10322
rect 2450 10180 2790 10266
rect 2450 10124 2521 10180
rect 2577 10124 2663 10180
rect 2719 10124 2790 10180
rect 2450 10038 2790 10124
rect 2450 9982 2521 10038
rect 2577 9982 2663 10038
rect 2719 9982 2790 10038
rect 2450 9896 2790 9982
rect 2450 9840 2521 9896
rect 2577 9840 2663 9896
rect 2719 9840 2790 9896
rect 2450 9754 2790 9840
rect 2450 9698 2521 9754
rect 2577 9698 2663 9754
rect 2719 9698 2790 9754
rect 2450 9612 2790 9698
rect 2450 9556 2521 9612
rect 2577 9556 2663 9612
rect 2719 9556 2790 9612
rect 2450 9470 2790 9556
rect 2450 9414 2521 9470
rect 2577 9414 2663 9470
rect 2719 9414 2790 9470
rect 2450 9328 2790 9414
rect 2450 9272 2521 9328
rect 2577 9272 2663 9328
rect 2719 9272 2790 9328
rect 2450 9186 2790 9272
rect 2450 9130 2521 9186
rect 2577 9130 2663 9186
rect 2719 9130 2790 9186
rect 2450 9044 2790 9130
rect 2450 8988 2521 9044
rect 2577 8988 2663 9044
rect 2719 8988 2790 9044
rect 2450 8902 2790 8988
rect 2450 8846 2521 8902
rect 2577 8846 2663 8902
rect 2719 8846 2790 8902
rect 2450 8760 2790 8846
rect 2450 8704 2521 8760
rect 2577 8704 2663 8760
rect 2719 8704 2790 8760
rect 2450 8618 2790 8704
rect 2450 8562 2521 8618
rect 2577 8562 2663 8618
rect 2719 8562 2790 8618
rect 2450 8476 2790 8562
rect 2450 8420 2521 8476
rect 2577 8420 2663 8476
rect 2719 8420 2790 8476
rect 2450 8334 2790 8420
rect 2450 8278 2521 8334
rect 2577 8278 2663 8334
rect 2719 8278 2790 8334
rect 2450 8192 2790 8278
rect 2450 8136 2521 8192
rect 2577 8136 2663 8192
rect 2719 8136 2790 8192
rect 2450 8050 2790 8136
rect 2450 7994 2521 8050
rect 2577 7994 2663 8050
rect 2719 7994 2790 8050
rect 2450 7908 2790 7994
rect 2450 7852 2521 7908
rect 2577 7852 2663 7908
rect 2719 7852 2790 7908
rect 2450 7766 2790 7852
rect 2450 7710 2521 7766
rect 2577 7710 2663 7766
rect 2719 7710 2790 7766
rect 2450 7624 2790 7710
rect 2450 7568 2521 7624
rect 2577 7568 2663 7624
rect 2719 7568 2790 7624
rect 2450 7482 2790 7568
rect 2450 7426 2521 7482
rect 2577 7426 2663 7482
rect 2719 7426 2790 7482
rect 2450 7340 2790 7426
rect 2450 7284 2521 7340
rect 2577 7284 2663 7340
rect 2719 7284 2790 7340
rect 2450 7198 2790 7284
rect 2450 7142 2521 7198
rect 2577 7142 2663 7198
rect 2719 7142 2790 7198
rect 2450 7056 2790 7142
rect 2450 7000 2521 7056
rect 2577 7000 2663 7056
rect 2719 7000 2790 7056
rect 2450 6914 2790 7000
rect 2450 6858 2521 6914
rect 2577 6858 2663 6914
rect 2719 6858 2790 6914
rect 2450 6772 2790 6858
rect 2450 6716 2521 6772
rect 2577 6716 2663 6772
rect 2719 6716 2790 6772
rect 2450 6630 2790 6716
rect 2450 6574 2521 6630
rect 2577 6574 2663 6630
rect 2719 6574 2790 6630
rect 2450 6488 2790 6574
rect 2450 6432 2521 6488
rect 2577 6432 2663 6488
rect 2719 6432 2790 6488
rect 2450 6346 2790 6432
rect 2450 6290 2521 6346
rect 2577 6290 2663 6346
rect 2719 6290 2790 6346
rect 2450 6204 2790 6290
rect 2450 6148 2521 6204
rect 2577 6148 2663 6204
rect 2719 6148 2790 6204
rect 2450 6062 2790 6148
rect 2450 6006 2521 6062
rect 2577 6006 2663 6062
rect 2719 6006 2790 6062
rect 2450 5920 2790 6006
rect 2450 5864 2521 5920
rect 2577 5864 2663 5920
rect 2719 5864 2790 5920
rect 2450 5778 2790 5864
rect 2450 5722 2521 5778
rect 2577 5722 2663 5778
rect 2719 5722 2790 5778
rect 2450 5636 2790 5722
rect 2450 5580 2521 5636
rect 2577 5580 2663 5636
rect 2719 5580 2790 5636
rect 2450 5494 2790 5580
rect 2450 5438 2521 5494
rect 2577 5438 2663 5494
rect 2719 5438 2790 5494
rect 2450 5352 2790 5438
rect 2450 5296 2521 5352
rect 2577 5296 2663 5352
rect 2719 5296 2790 5352
rect 2450 5210 2790 5296
rect 2450 5154 2521 5210
rect 2577 5154 2663 5210
rect 2719 5154 2790 5210
rect 2450 5068 2790 5154
rect 2450 5012 2521 5068
rect 2577 5012 2663 5068
rect 2719 5012 2790 5068
rect 2450 4926 2790 5012
rect 2450 4870 2521 4926
rect 2577 4870 2663 4926
rect 2719 4870 2790 4926
rect 2450 4784 2790 4870
rect 2450 4728 2521 4784
rect 2577 4728 2663 4784
rect 2719 4728 2790 4784
rect 2450 4642 2790 4728
rect 2450 4586 2521 4642
rect 2577 4586 2663 4642
rect 2719 4586 2790 4642
rect 2450 4500 2790 4586
rect 2450 4444 2521 4500
rect 2577 4444 2663 4500
rect 2719 4444 2790 4500
rect 2450 4358 2790 4444
rect 2450 4302 2521 4358
rect 2577 4302 2663 4358
rect 2719 4302 2790 4358
rect 2450 4216 2790 4302
rect 2450 4160 2521 4216
rect 2577 4160 2663 4216
rect 2719 4160 2790 4216
rect 2450 4074 2790 4160
rect 2450 4018 2521 4074
rect 2577 4018 2663 4074
rect 2719 4018 2790 4074
rect 2450 3932 2790 4018
rect 2450 3876 2521 3932
rect 2577 3876 2663 3932
rect 2719 3876 2790 3932
rect 2450 3790 2790 3876
rect 2450 3734 2521 3790
rect 2577 3734 2663 3790
rect 2719 3734 2790 3790
rect 2450 3648 2790 3734
rect 2450 3592 2521 3648
rect 2577 3592 2663 3648
rect 2719 3592 2790 3648
rect 2450 3506 2790 3592
rect 2450 3450 2521 3506
rect 2577 3450 2663 3506
rect 2719 3450 2790 3506
rect 2450 3364 2790 3450
rect 2450 3308 2521 3364
rect 2577 3308 2663 3364
rect 2719 3308 2790 3364
rect 2450 3222 2790 3308
rect 2450 3166 2521 3222
rect 2577 3166 2663 3222
rect 2719 3166 2790 3222
rect 2450 3080 2790 3166
rect 2450 3024 2521 3080
rect 2577 3024 2663 3080
rect 2719 3024 2790 3080
rect 2450 2938 2790 3024
rect 2450 2882 2521 2938
rect 2577 2882 2663 2938
rect 2719 2882 2790 2938
rect 2450 2796 2790 2882
rect 2450 2740 2521 2796
rect 2577 2740 2663 2796
rect 2719 2740 2790 2796
rect 2450 2654 2790 2740
rect 2450 2598 2521 2654
rect 2577 2598 2663 2654
rect 2719 2598 2790 2654
rect 2450 2512 2790 2598
rect 2450 2456 2521 2512
rect 2577 2456 2663 2512
rect 2719 2456 2790 2512
rect 2450 2370 2790 2456
rect 2450 2314 2521 2370
rect 2577 2314 2663 2370
rect 2719 2314 2790 2370
rect 2450 2228 2790 2314
rect 2450 2172 2521 2228
rect 2577 2172 2663 2228
rect 2719 2172 2790 2228
rect 2450 2086 2790 2172
rect 2450 2030 2521 2086
rect 2577 2030 2663 2086
rect 2719 2030 2790 2086
rect 2450 1944 2790 2030
rect 2450 1888 2521 1944
rect 2577 1888 2663 1944
rect 2719 1888 2790 1944
rect 2450 1802 2790 1888
rect 2450 1746 2521 1802
rect 2577 1746 2663 1802
rect 2719 1746 2790 1802
rect 2450 1660 2790 1746
rect 2450 1604 2521 1660
rect 2577 1604 2663 1660
rect 2719 1604 2790 1660
rect 2450 1518 2790 1604
rect 2450 1462 2521 1518
rect 2577 1462 2663 1518
rect 2719 1462 2790 1518
rect 2450 1376 2790 1462
rect 2450 1320 2521 1376
rect 2577 1320 2663 1376
rect 2719 1320 2790 1376
rect 2450 1234 2790 1320
rect 2450 1178 2521 1234
rect 2577 1178 2663 1234
rect 2719 1178 2790 1234
rect 2450 1092 2790 1178
rect 2450 1036 2521 1092
rect 2577 1036 2663 1092
rect 2719 1036 2790 1092
rect 2450 950 2790 1036
rect 2450 894 2521 950
rect 2577 894 2663 950
rect 2719 894 2790 950
rect 2450 808 2790 894
rect 2450 752 2521 808
rect 2577 752 2663 808
rect 2719 752 2790 808
rect 2450 666 2790 752
rect 2450 610 2521 666
rect 2577 610 2663 666
rect 2719 610 2790 666
rect 2450 524 2790 610
rect 2450 468 2521 524
rect 2577 468 2663 524
rect 2719 468 2790 524
rect 2450 458 2790 468
rect 2990 12310 3330 12320
rect 2990 12254 3058 12310
rect 3114 12254 3200 12310
rect 3256 12254 3330 12310
rect 2990 12168 3330 12254
rect 2990 12112 3058 12168
rect 3114 12112 3200 12168
rect 3256 12112 3330 12168
rect 2990 12026 3330 12112
rect 2990 11970 3058 12026
rect 3114 11970 3200 12026
rect 3256 11970 3330 12026
rect 2990 11884 3330 11970
rect 2990 11828 3058 11884
rect 3114 11828 3200 11884
rect 3256 11828 3330 11884
rect 2990 11742 3330 11828
rect 2990 11686 3058 11742
rect 3114 11686 3200 11742
rect 3256 11686 3330 11742
rect 2990 11600 3330 11686
rect 2990 11544 3058 11600
rect 3114 11544 3200 11600
rect 3256 11544 3330 11600
rect 2990 11458 3330 11544
rect 2990 11402 3058 11458
rect 3114 11402 3200 11458
rect 3256 11402 3330 11458
rect 2990 11316 3330 11402
rect 2990 11260 3058 11316
rect 3114 11260 3200 11316
rect 3256 11260 3330 11316
rect 2990 11174 3330 11260
rect 2990 11118 3058 11174
rect 3114 11118 3200 11174
rect 3256 11118 3330 11174
rect 2990 11032 3330 11118
rect 2990 10976 3058 11032
rect 3114 10976 3200 11032
rect 3256 10976 3330 11032
rect 2990 10890 3330 10976
rect 2990 10834 3058 10890
rect 3114 10834 3200 10890
rect 3256 10834 3330 10890
rect 2990 10748 3330 10834
rect 2990 10692 3058 10748
rect 3114 10692 3200 10748
rect 3256 10692 3330 10748
rect 2990 10606 3330 10692
rect 2990 10550 3058 10606
rect 3114 10550 3200 10606
rect 3256 10550 3330 10606
rect 2990 10464 3330 10550
rect 2990 10408 3058 10464
rect 3114 10408 3200 10464
rect 3256 10408 3330 10464
rect 2990 10322 3330 10408
rect 2990 10266 3058 10322
rect 3114 10266 3200 10322
rect 3256 10266 3330 10322
rect 2990 10180 3330 10266
rect 2990 10124 3058 10180
rect 3114 10124 3200 10180
rect 3256 10124 3330 10180
rect 2990 10038 3330 10124
rect 2990 9982 3058 10038
rect 3114 9982 3200 10038
rect 3256 9982 3330 10038
rect 2990 9896 3330 9982
rect 2990 9840 3058 9896
rect 3114 9840 3200 9896
rect 3256 9840 3330 9896
rect 2990 9754 3330 9840
rect 2990 9698 3058 9754
rect 3114 9698 3200 9754
rect 3256 9698 3330 9754
rect 2990 9612 3330 9698
rect 2990 9556 3058 9612
rect 3114 9556 3200 9612
rect 3256 9556 3330 9612
rect 2990 9470 3330 9556
rect 2990 9414 3058 9470
rect 3114 9414 3200 9470
rect 3256 9414 3330 9470
rect 2990 9328 3330 9414
rect 2990 9272 3058 9328
rect 3114 9272 3200 9328
rect 3256 9272 3330 9328
rect 2990 9186 3330 9272
rect 2990 9130 3058 9186
rect 3114 9130 3200 9186
rect 3256 9130 3330 9186
rect 2990 9044 3330 9130
rect 2990 8988 3058 9044
rect 3114 8988 3200 9044
rect 3256 8988 3330 9044
rect 2990 8902 3330 8988
rect 2990 8846 3058 8902
rect 3114 8846 3200 8902
rect 3256 8846 3330 8902
rect 2990 8760 3330 8846
rect 2990 8704 3058 8760
rect 3114 8704 3200 8760
rect 3256 8704 3330 8760
rect 2990 8618 3330 8704
rect 2990 8562 3058 8618
rect 3114 8562 3200 8618
rect 3256 8562 3330 8618
rect 2990 8476 3330 8562
rect 2990 8420 3058 8476
rect 3114 8420 3200 8476
rect 3256 8420 3330 8476
rect 2990 8334 3330 8420
rect 2990 8278 3058 8334
rect 3114 8278 3200 8334
rect 3256 8278 3330 8334
rect 2990 8192 3330 8278
rect 2990 8136 3058 8192
rect 3114 8136 3200 8192
rect 3256 8136 3330 8192
rect 2990 8050 3330 8136
rect 2990 7994 3058 8050
rect 3114 7994 3200 8050
rect 3256 7994 3330 8050
rect 2990 7908 3330 7994
rect 2990 7852 3058 7908
rect 3114 7852 3200 7908
rect 3256 7852 3330 7908
rect 2990 7766 3330 7852
rect 2990 7710 3058 7766
rect 3114 7710 3200 7766
rect 3256 7710 3330 7766
rect 2990 7624 3330 7710
rect 2990 7568 3058 7624
rect 3114 7568 3200 7624
rect 3256 7568 3330 7624
rect 2990 7482 3330 7568
rect 2990 7426 3058 7482
rect 3114 7426 3200 7482
rect 3256 7426 3330 7482
rect 2990 7340 3330 7426
rect 2990 7284 3058 7340
rect 3114 7284 3200 7340
rect 3256 7284 3330 7340
rect 2990 7198 3330 7284
rect 2990 7142 3058 7198
rect 3114 7142 3200 7198
rect 3256 7142 3330 7198
rect 2990 7056 3330 7142
rect 2990 7000 3058 7056
rect 3114 7000 3200 7056
rect 3256 7000 3330 7056
rect 2990 6914 3330 7000
rect 2990 6858 3058 6914
rect 3114 6858 3200 6914
rect 3256 6858 3330 6914
rect 2990 6772 3330 6858
rect 2990 6716 3058 6772
rect 3114 6716 3200 6772
rect 3256 6716 3330 6772
rect 2990 6630 3330 6716
rect 2990 6574 3058 6630
rect 3114 6574 3200 6630
rect 3256 6574 3330 6630
rect 2990 6488 3330 6574
rect 2990 6432 3058 6488
rect 3114 6432 3200 6488
rect 3256 6432 3330 6488
rect 2990 6346 3330 6432
rect 2990 6290 3058 6346
rect 3114 6290 3200 6346
rect 3256 6290 3330 6346
rect 2990 6204 3330 6290
rect 2990 6148 3058 6204
rect 3114 6148 3200 6204
rect 3256 6148 3330 6204
rect 2990 6062 3330 6148
rect 2990 6006 3058 6062
rect 3114 6006 3200 6062
rect 3256 6006 3330 6062
rect 2990 5920 3330 6006
rect 2990 5864 3058 5920
rect 3114 5864 3200 5920
rect 3256 5864 3330 5920
rect 2990 5778 3330 5864
rect 2990 5722 3058 5778
rect 3114 5722 3200 5778
rect 3256 5722 3330 5778
rect 2990 5636 3330 5722
rect 2990 5580 3058 5636
rect 3114 5580 3200 5636
rect 3256 5580 3330 5636
rect 2990 5494 3330 5580
rect 2990 5438 3058 5494
rect 3114 5438 3200 5494
rect 3256 5438 3330 5494
rect 2990 5352 3330 5438
rect 2990 5296 3058 5352
rect 3114 5296 3200 5352
rect 3256 5296 3330 5352
rect 2990 5210 3330 5296
rect 2990 5154 3058 5210
rect 3114 5154 3200 5210
rect 3256 5154 3330 5210
rect 2990 5068 3330 5154
rect 2990 5012 3058 5068
rect 3114 5012 3200 5068
rect 3256 5012 3330 5068
rect 2990 4926 3330 5012
rect 2990 4870 3058 4926
rect 3114 4870 3200 4926
rect 3256 4870 3330 4926
rect 2990 4784 3330 4870
rect 2990 4728 3058 4784
rect 3114 4728 3200 4784
rect 3256 4728 3330 4784
rect 2990 4642 3330 4728
rect 2990 4586 3058 4642
rect 3114 4586 3200 4642
rect 3256 4586 3330 4642
rect 2990 4500 3330 4586
rect 2990 4444 3058 4500
rect 3114 4444 3200 4500
rect 3256 4444 3330 4500
rect 2990 4358 3330 4444
rect 2990 4302 3058 4358
rect 3114 4302 3200 4358
rect 3256 4302 3330 4358
rect 2990 4216 3330 4302
rect 2990 4160 3058 4216
rect 3114 4160 3200 4216
rect 3256 4160 3330 4216
rect 2990 4074 3330 4160
rect 2990 4018 3058 4074
rect 3114 4018 3200 4074
rect 3256 4018 3330 4074
rect 2990 3932 3330 4018
rect 2990 3876 3058 3932
rect 3114 3876 3200 3932
rect 3256 3876 3330 3932
rect 2990 3790 3330 3876
rect 2990 3734 3058 3790
rect 3114 3734 3200 3790
rect 3256 3734 3330 3790
rect 2990 3648 3330 3734
rect 2990 3592 3058 3648
rect 3114 3592 3200 3648
rect 3256 3592 3330 3648
rect 2990 3506 3330 3592
rect 2990 3450 3058 3506
rect 3114 3450 3200 3506
rect 3256 3450 3330 3506
rect 2990 3364 3330 3450
rect 2990 3308 3058 3364
rect 3114 3308 3200 3364
rect 3256 3308 3330 3364
rect 2990 3222 3330 3308
rect 2990 3166 3058 3222
rect 3114 3166 3200 3222
rect 3256 3166 3330 3222
rect 2990 3080 3330 3166
rect 2990 3024 3058 3080
rect 3114 3024 3200 3080
rect 3256 3024 3330 3080
rect 2990 2938 3330 3024
rect 2990 2882 3058 2938
rect 3114 2882 3200 2938
rect 3256 2882 3330 2938
rect 2990 2796 3330 2882
rect 2990 2740 3058 2796
rect 3114 2740 3200 2796
rect 3256 2740 3330 2796
rect 2990 2654 3330 2740
rect 2990 2598 3058 2654
rect 3114 2598 3200 2654
rect 3256 2598 3330 2654
rect 2990 2512 3330 2598
rect 2990 2456 3058 2512
rect 3114 2456 3200 2512
rect 3256 2456 3330 2512
rect 2990 2370 3330 2456
rect 2990 2314 3058 2370
rect 3114 2314 3200 2370
rect 3256 2314 3330 2370
rect 2990 2228 3330 2314
rect 2990 2172 3058 2228
rect 3114 2172 3200 2228
rect 3256 2172 3330 2228
rect 2990 2086 3330 2172
rect 2990 2030 3058 2086
rect 3114 2030 3200 2086
rect 3256 2030 3330 2086
rect 2990 1944 3330 2030
rect 2990 1888 3058 1944
rect 3114 1888 3200 1944
rect 3256 1888 3330 1944
rect 2990 1802 3330 1888
rect 2990 1746 3058 1802
rect 3114 1746 3200 1802
rect 3256 1746 3330 1802
rect 2990 1660 3330 1746
rect 2990 1604 3058 1660
rect 3114 1604 3200 1660
rect 3256 1604 3330 1660
rect 2990 1518 3330 1604
rect 2990 1462 3058 1518
rect 3114 1462 3200 1518
rect 3256 1462 3330 1518
rect 2990 1376 3330 1462
rect 2990 1320 3058 1376
rect 3114 1320 3200 1376
rect 3256 1320 3330 1376
rect 2990 1234 3330 1320
rect 2990 1178 3058 1234
rect 3114 1178 3200 1234
rect 3256 1178 3330 1234
rect 2990 1092 3330 1178
rect 2990 1036 3058 1092
rect 3114 1036 3200 1092
rect 3256 1036 3330 1092
rect 2990 950 3330 1036
rect 2990 894 3058 950
rect 3114 894 3200 950
rect 3256 894 3330 950
rect 2990 808 3330 894
rect 2990 752 3058 808
rect 3114 752 3200 808
rect 3256 752 3330 808
rect 2990 666 3330 752
rect 2990 610 3058 666
rect 3114 610 3200 666
rect 3256 610 3330 666
rect 2990 524 3330 610
rect 2990 468 3058 524
rect 3114 468 3200 524
rect 3256 468 3330 524
rect 2990 458 3330 468
rect 3530 12310 3870 12320
rect 3530 12254 3602 12310
rect 3658 12254 3744 12310
rect 3800 12254 3870 12310
rect 3530 12168 3870 12254
rect 3530 12112 3602 12168
rect 3658 12112 3744 12168
rect 3800 12112 3870 12168
rect 3530 12026 3870 12112
rect 3530 11970 3602 12026
rect 3658 11970 3744 12026
rect 3800 11970 3870 12026
rect 3530 11884 3870 11970
rect 3530 11828 3602 11884
rect 3658 11828 3744 11884
rect 3800 11828 3870 11884
rect 3530 11742 3870 11828
rect 3530 11686 3602 11742
rect 3658 11686 3744 11742
rect 3800 11686 3870 11742
rect 3530 11600 3870 11686
rect 3530 11544 3602 11600
rect 3658 11544 3744 11600
rect 3800 11544 3870 11600
rect 3530 11458 3870 11544
rect 3530 11402 3602 11458
rect 3658 11402 3744 11458
rect 3800 11402 3870 11458
rect 3530 11316 3870 11402
rect 3530 11260 3602 11316
rect 3658 11260 3744 11316
rect 3800 11260 3870 11316
rect 3530 11174 3870 11260
rect 3530 11118 3602 11174
rect 3658 11118 3744 11174
rect 3800 11118 3870 11174
rect 3530 11032 3870 11118
rect 3530 10976 3602 11032
rect 3658 10976 3744 11032
rect 3800 10976 3870 11032
rect 3530 10890 3870 10976
rect 3530 10834 3602 10890
rect 3658 10834 3744 10890
rect 3800 10834 3870 10890
rect 3530 10748 3870 10834
rect 3530 10692 3602 10748
rect 3658 10692 3744 10748
rect 3800 10692 3870 10748
rect 3530 10606 3870 10692
rect 3530 10550 3602 10606
rect 3658 10550 3744 10606
rect 3800 10550 3870 10606
rect 3530 10464 3870 10550
rect 3530 10408 3602 10464
rect 3658 10408 3744 10464
rect 3800 10408 3870 10464
rect 3530 10322 3870 10408
rect 3530 10266 3602 10322
rect 3658 10266 3744 10322
rect 3800 10266 3870 10322
rect 3530 10180 3870 10266
rect 3530 10124 3602 10180
rect 3658 10124 3744 10180
rect 3800 10124 3870 10180
rect 3530 10038 3870 10124
rect 3530 9982 3602 10038
rect 3658 9982 3744 10038
rect 3800 9982 3870 10038
rect 3530 9896 3870 9982
rect 3530 9840 3602 9896
rect 3658 9840 3744 9896
rect 3800 9840 3870 9896
rect 3530 9754 3870 9840
rect 3530 9698 3602 9754
rect 3658 9698 3744 9754
rect 3800 9698 3870 9754
rect 3530 9612 3870 9698
rect 3530 9556 3602 9612
rect 3658 9556 3744 9612
rect 3800 9556 3870 9612
rect 3530 9470 3870 9556
rect 3530 9414 3602 9470
rect 3658 9414 3744 9470
rect 3800 9414 3870 9470
rect 3530 9328 3870 9414
rect 3530 9272 3602 9328
rect 3658 9272 3744 9328
rect 3800 9272 3870 9328
rect 3530 9186 3870 9272
rect 3530 9130 3602 9186
rect 3658 9130 3744 9186
rect 3800 9130 3870 9186
rect 3530 9044 3870 9130
rect 3530 8988 3602 9044
rect 3658 8988 3744 9044
rect 3800 8988 3870 9044
rect 3530 8902 3870 8988
rect 3530 8846 3602 8902
rect 3658 8846 3744 8902
rect 3800 8846 3870 8902
rect 3530 8760 3870 8846
rect 3530 8704 3602 8760
rect 3658 8704 3744 8760
rect 3800 8704 3870 8760
rect 3530 8618 3870 8704
rect 3530 8562 3602 8618
rect 3658 8562 3744 8618
rect 3800 8562 3870 8618
rect 3530 8476 3870 8562
rect 3530 8420 3602 8476
rect 3658 8420 3744 8476
rect 3800 8420 3870 8476
rect 3530 8334 3870 8420
rect 3530 8278 3602 8334
rect 3658 8278 3744 8334
rect 3800 8278 3870 8334
rect 3530 8192 3870 8278
rect 3530 8136 3602 8192
rect 3658 8136 3744 8192
rect 3800 8136 3870 8192
rect 3530 8050 3870 8136
rect 3530 7994 3602 8050
rect 3658 7994 3744 8050
rect 3800 7994 3870 8050
rect 3530 7908 3870 7994
rect 3530 7852 3602 7908
rect 3658 7852 3744 7908
rect 3800 7852 3870 7908
rect 3530 7766 3870 7852
rect 3530 7710 3602 7766
rect 3658 7710 3744 7766
rect 3800 7710 3870 7766
rect 3530 7624 3870 7710
rect 3530 7568 3602 7624
rect 3658 7568 3744 7624
rect 3800 7568 3870 7624
rect 3530 7482 3870 7568
rect 3530 7426 3602 7482
rect 3658 7426 3744 7482
rect 3800 7426 3870 7482
rect 3530 7340 3870 7426
rect 3530 7284 3602 7340
rect 3658 7284 3744 7340
rect 3800 7284 3870 7340
rect 3530 7198 3870 7284
rect 3530 7142 3602 7198
rect 3658 7142 3744 7198
rect 3800 7142 3870 7198
rect 3530 7056 3870 7142
rect 3530 7000 3602 7056
rect 3658 7000 3744 7056
rect 3800 7000 3870 7056
rect 3530 6914 3870 7000
rect 3530 6858 3602 6914
rect 3658 6858 3744 6914
rect 3800 6858 3870 6914
rect 3530 6772 3870 6858
rect 3530 6716 3602 6772
rect 3658 6716 3744 6772
rect 3800 6716 3870 6772
rect 3530 6630 3870 6716
rect 3530 6574 3602 6630
rect 3658 6574 3744 6630
rect 3800 6574 3870 6630
rect 3530 6488 3870 6574
rect 3530 6432 3602 6488
rect 3658 6432 3744 6488
rect 3800 6432 3870 6488
rect 3530 6346 3870 6432
rect 3530 6290 3602 6346
rect 3658 6290 3744 6346
rect 3800 6290 3870 6346
rect 3530 6204 3870 6290
rect 3530 6148 3602 6204
rect 3658 6148 3744 6204
rect 3800 6148 3870 6204
rect 3530 6062 3870 6148
rect 3530 6006 3602 6062
rect 3658 6006 3744 6062
rect 3800 6006 3870 6062
rect 3530 5920 3870 6006
rect 3530 5864 3602 5920
rect 3658 5864 3744 5920
rect 3800 5864 3870 5920
rect 3530 5778 3870 5864
rect 3530 5722 3602 5778
rect 3658 5722 3744 5778
rect 3800 5722 3870 5778
rect 3530 5636 3870 5722
rect 3530 5580 3602 5636
rect 3658 5580 3744 5636
rect 3800 5580 3870 5636
rect 3530 5494 3870 5580
rect 3530 5438 3602 5494
rect 3658 5438 3744 5494
rect 3800 5438 3870 5494
rect 3530 5352 3870 5438
rect 3530 5296 3602 5352
rect 3658 5296 3744 5352
rect 3800 5296 3870 5352
rect 3530 5210 3870 5296
rect 3530 5154 3602 5210
rect 3658 5154 3744 5210
rect 3800 5154 3870 5210
rect 3530 5068 3870 5154
rect 3530 5012 3602 5068
rect 3658 5012 3744 5068
rect 3800 5012 3870 5068
rect 3530 4926 3870 5012
rect 3530 4870 3602 4926
rect 3658 4870 3744 4926
rect 3800 4870 3870 4926
rect 3530 4784 3870 4870
rect 3530 4728 3602 4784
rect 3658 4728 3744 4784
rect 3800 4728 3870 4784
rect 3530 4642 3870 4728
rect 3530 4586 3602 4642
rect 3658 4586 3744 4642
rect 3800 4586 3870 4642
rect 3530 4500 3870 4586
rect 3530 4444 3602 4500
rect 3658 4444 3744 4500
rect 3800 4444 3870 4500
rect 3530 4358 3870 4444
rect 3530 4302 3602 4358
rect 3658 4302 3744 4358
rect 3800 4302 3870 4358
rect 3530 4216 3870 4302
rect 3530 4160 3602 4216
rect 3658 4160 3744 4216
rect 3800 4160 3870 4216
rect 3530 4074 3870 4160
rect 3530 4018 3602 4074
rect 3658 4018 3744 4074
rect 3800 4018 3870 4074
rect 3530 3932 3870 4018
rect 3530 3876 3602 3932
rect 3658 3876 3744 3932
rect 3800 3876 3870 3932
rect 3530 3790 3870 3876
rect 3530 3734 3602 3790
rect 3658 3734 3744 3790
rect 3800 3734 3870 3790
rect 3530 3648 3870 3734
rect 3530 3592 3602 3648
rect 3658 3592 3744 3648
rect 3800 3592 3870 3648
rect 3530 3506 3870 3592
rect 3530 3450 3602 3506
rect 3658 3450 3744 3506
rect 3800 3450 3870 3506
rect 3530 3364 3870 3450
rect 3530 3308 3602 3364
rect 3658 3308 3744 3364
rect 3800 3308 3870 3364
rect 3530 3222 3870 3308
rect 3530 3166 3602 3222
rect 3658 3166 3744 3222
rect 3800 3166 3870 3222
rect 3530 3080 3870 3166
rect 3530 3024 3602 3080
rect 3658 3024 3744 3080
rect 3800 3024 3870 3080
rect 3530 2938 3870 3024
rect 3530 2882 3602 2938
rect 3658 2882 3744 2938
rect 3800 2882 3870 2938
rect 3530 2796 3870 2882
rect 3530 2740 3602 2796
rect 3658 2740 3744 2796
rect 3800 2740 3870 2796
rect 3530 2654 3870 2740
rect 3530 2598 3602 2654
rect 3658 2598 3744 2654
rect 3800 2598 3870 2654
rect 3530 2512 3870 2598
rect 3530 2456 3602 2512
rect 3658 2456 3744 2512
rect 3800 2456 3870 2512
rect 3530 2370 3870 2456
rect 3530 2314 3602 2370
rect 3658 2314 3744 2370
rect 3800 2314 3870 2370
rect 3530 2228 3870 2314
rect 3530 2172 3602 2228
rect 3658 2172 3744 2228
rect 3800 2172 3870 2228
rect 3530 2086 3870 2172
rect 3530 2030 3602 2086
rect 3658 2030 3744 2086
rect 3800 2030 3870 2086
rect 3530 1944 3870 2030
rect 3530 1888 3602 1944
rect 3658 1888 3744 1944
rect 3800 1888 3870 1944
rect 3530 1802 3870 1888
rect 3530 1746 3602 1802
rect 3658 1746 3744 1802
rect 3800 1746 3870 1802
rect 3530 1660 3870 1746
rect 3530 1604 3602 1660
rect 3658 1604 3744 1660
rect 3800 1604 3870 1660
rect 3530 1518 3870 1604
rect 3530 1462 3602 1518
rect 3658 1462 3744 1518
rect 3800 1462 3870 1518
rect 3530 1376 3870 1462
rect 3530 1320 3602 1376
rect 3658 1320 3744 1376
rect 3800 1320 3870 1376
rect 3530 1234 3870 1320
rect 3530 1178 3602 1234
rect 3658 1178 3744 1234
rect 3800 1178 3870 1234
rect 3530 1092 3870 1178
rect 3530 1036 3602 1092
rect 3658 1036 3744 1092
rect 3800 1036 3870 1092
rect 3530 950 3870 1036
rect 3530 894 3602 950
rect 3658 894 3744 950
rect 3800 894 3870 950
rect 3530 808 3870 894
rect 3530 752 3602 808
rect 3658 752 3744 808
rect 3800 752 3870 808
rect 3530 666 3870 752
rect 3530 610 3602 666
rect 3658 610 3744 666
rect 3800 610 3870 666
rect 3530 524 3870 610
rect 3530 468 3602 524
rect 3658 468 3744 524
rect 3800 468 3870 524
rect 3530 458 3870 468
rect 4070 12310 4410 12320
rect 4070 12254 4138 12310
rect 4194 12254 4280 12310
rect 4336 12254 4410 12310
rect 4070 12168 4410 12254
rect 4070 12112 4138 12168
rect 4194 12112 4280 12168
rect 4336 12112 4410 12168
rect 4070 12026 4410 12112
rect 4070 11970 4138 12026
rect 4194 11970 4280 12026
rect 4336 11970 4410 12026
rect 4070 11884 4410 11970
rect 4070 11828 4138 11884
rect 4194 11828 4280 11884
rect 4336 11828 4410 11884
rect 4070 11742 4410 11828
rect 4070 11686 4138 11742
rect 4194 11686 4280 11742
rect 4336 11686 4410 11742
rect 4070 11600 4410 11686
rect 4070 11544 4138 11600
rect 4194 11544 4280 11600
rect 4336 11544 4410 11600
rect 4070 11458 4410 11544
rect 4070 11402 4138 11458
rect 4194 11402 4280 11458
rect 4336 11402 4410 11458
rect 4070 11316 4410 11402
rect 4070 11260 4138 11316
rect 4194 11260 4280 11316
rect 4336 11260 4410 11316
rect 4070 11174 4410 11260
rect 4070 11118 4138 11174
rect 4194 11118 4280 11174
rect 4336 11118 4410 11174
rect 4070 11032 4410 11118
rect 4070 10976 4138 11032
rect 4194 10976 4280 11032
rect 4336 10976 4410 11032
rect 4070 10890 4410 10976
rect 4070 10834 4138 10890
rect 4194 10834 4280 10890
rect 4336 10834 4410 10890
rect 4070 10748 4410 10834
rect 4070 10692 4138 10748
rect 4194 10692 4280 10748
rect 4336 10692 4410 10748
rect 4070 10606 4410 10692
rect 4070 10550 4138 10606
rect 4194 10550 4280 10606
rect 4336 10550 4410 10606
rect 4070 10464 4410 10550
rect 4070 10408 4138 10464
rect 4194 10408 4280 10464
rect 4336 10408 4410 10464
rect 4070 10322 4410 10408
rect 4070 10266 4138 10322
rect 4194 10266 4280 10322
rect 4336 10266 4410 10322
rect 4070 10180 4410 10266
rect 4070 10124 4138 10180
rect 4194 10124 4280 10180
rect 4336 10124 4410 10180
rect 4070 10038 4410 10124
rect 4070 9982 4138 10038
rect 4194 9982 4280 10038
rect 4336 9982 4410 10038
rect 4070 9896 4410 9982
rect 4070 9840 4138 9896
rect 4194 9840 4280 9896
rect 4336 9840 4410 9896
rect 4070 9754 4410 9840
rect 4070 9698 4138 9754
rect 4194 9698 4280 9754
rect 4336 9698 4410 9754
rect 4070 9612 4410 9698
rect 4070 9556 4138 9612
rect 4194 9556 4280 9612
rect 4336 9556 4410 9612
rect 4070 9470 4410 9556
rect 4070 9414 4138 9470
rect 4194 9414 4280 9470
rect 4336 9414 4410 9470
rect 4070 9328 4410 9414
rect 4070 9272 4138 9328
rect 4194 9272 4280 9328
rect 4336 9272 4410 9328
rect 4070 9186 4410 9272
rect 4070 9130 4138 9186
rect 4194 9130 4280 9186
rect 4336 9130 4410 9186
rect 4070 9044 4410 9130
rect 4070 8988 4138 9044
rect 4194 8988 4280 9044
rect 4336 8988 4410 9044
rect 4070 8902 4410 8988
rect 4070 8846 4138 8902
rect 4194 8846 4280 8902
rect 4336 8846 4410 8902
rect 4070 8760 4410 8846
rect 4070 8704 4138 8760
rect 4194 8704 4280 8760
rect 4336 8704 4410 8760
rect 4070 8618 4410 8704
rect 4070 8562 4138 8618
rect 4194 8562 4280 8618
rect 4336 8562 4410 8618
rect 4070 8476 4410 8562
rect 4070 8420 4138 8476
rect 4194 8420 4280 8476
rect 4336 8420 4410 8476
rect 4070 8334 4410 8420
rect 4070 8278 4138 8334
rect 4194 8278 4280 8334
rect 4336 8278 4410 8334
rect 4070 8192 4410 8278
rect 4070 8136 4138 8192
rect 4194 8136 4280 8192
rect 4336 8136 4410 8192
rect 4070 8050 4410 8136
rect 4070 7994 4138 8050
rect 4194 7994 4280 8050
rect 4336 7994 4410 8050
rect 4070 7908 4410 7994
rect 4070 7852 4138 7908
rect 4194 7852 4280 7908
rect 4336 7852 4410 7908
rect 4070 7766 4410 7852
rect 4070 7710 4138 7766
rect 4194 7710 4280 7766
rect 4336 7710 4410 7766
rect 4070 7624 4410 7710
rect 4070 7568 4138 7624
rect 4194 7568 4280 7624
rect 4336 7568 4410 7624
rect 4070 7482 4410 7568
rect 4070 7426 4138 7482
rect 4194 7426 4280 7482
rect 4336 7426 4410 7482
rect 4070 7340 4410 7426
rect 4070 7284 4138 7340
rect 4194 7284 4280 7340
rect 4336 7284 4410 7340
rect 4070 7198 4410 7284
rect 4070 7142 4138 7198
rect 4194 7142 4280 7198
rect 4336 7142 4410 7198
rect 4070 7056 4410 7142
rect 4070 7000 4138 7056
rect 4194 7000 4280 7056
rect 4336 7000 4410 7056
rect 4070 6914 4410 7000
rect 4070 6858 4138 6914
rect 4194 6858 4280 6914
rect 4336 6858 4410 6914
rect 4070 6772 4410 6858
rect 4070 6716 4138 6772
rect 4194 6716 4280 6772
rect 4336 6716 4410 6772
rect 4070 6630 4410 6716
rect 4070 6574 4138 6630
rect 4194 6574 4280 6630
rect 4336 6574 4410 6630
rect 4070 6488 4410 6574
rect 4070 6432 4138 6488
rect 4194 6432 4280 6488
rect 4336 6432 4410 6488
rect 4070 6346 4410 6432
rect 4070 6290 4138 6346
rect 4194 6290 4280 6346
rect 4336 6290 4410 6346
rect 4070 6204 4410 6290
rect 4070 6148 4138 6204
rect 4194 6148 4280 6204
rect 4336 6148 4410 6204
rect 4070 6062 4410 6148
rect 4070 6006 4138 6062
rect 4194 6006 4280 6062
rect 4336 6006 4410 6062
rect 4070 5920 4410 6006
rect 4070 5864 4138 5920
rect 4194 5864 4280 5920
rect 4336 5864 4410 5920
rect 4070 5778 4410 5864
rect 4070 5722 4138 5778
rect 4194 5722 4280 5778
rect 4336 5722 4410 5778
rect 4070 5636 4410 5722
rect 4070 5580 4138 5636
rect 4194 5580 4280 5636
rect 4336 5580 4410 5636
rect 4070 5494 4410 5580
rect 4070 5438 4138 5494
rect 4194 5438 4280 5494
rect 4336 5438 4410 5494
rect 4070 5352 4410 5438
rect 4070 5296 4138 5352
rect 4194 5296 4280 5352
rect 4336 5296 4410 5352
rect 4070 5210 4410 5296
rect 4070 5154 4138 5210
rect 4194 5154 4280 5210
rect 4336 5154 4410 5210
rect 4070 5068 4410 5154
rect 4070 5012 4138 5068
rect 4194 5012 4280 5068
rect 4336 5012 4410 5068
rect 4070 4926 4410 5012
rect 4070 4870 4138 4926
rect 4194 4870 4280 4926
rect 4336 4870 4410 4926
rect 4070 4784 4410 4870
rect 4070 4728 4138 4784
rect 4194 4728 4280 4784
rect 4336 4728 4410 4784
rect 4070 4642 4410 4728
rect 4070 4586 4138 4642
rect 4194 4586 4280 4642
rect 4336 4586 4410 4642
rect 4070 4500 4410 4586
rect 4070 4444 4138 4500
rect 4194 4444 4280 4500
rect 4336 4444 4410 4500
rect 4070 4358 4410 4444
rect 4070 4302 4138 4358
rect 4194 4302 4280 4358
rect 4336 4302 4410 4358
rect 4070 4216 4410 4302
rect 4070 4160 4138 4216
rect 4194 4160 4280 4216
rect 4336 4160 4410 4216
rect 4070 4074 4410 4160
rect 4070 4018 4138 4074
rect 4194 4018 4280 4074
rect 4336 4018 4410 4074
rect 4070 3932 4410 4018
rect 4070 3876 4138 3932
rect 4194 3876 4280 3932
rect 4336 3876 4410 3932
rect 4070 3790 4410 3876
rect 4070 3734 4138 3790
rect 4194 3734 4280 3790
rect 4336 3734 4410 3790
rect 4070 3648 4410 3734
rect 4070 3592 4138 3648
rect 4194 3592 4280 3648
rect 4336 3592 4410 3648
rect 4070 3506 4410 3592
rect 4070 3450 4138 3506
rect 4194 3450 4280 3506
rect 4336 3450 4410 3506
rect 4070 3364 4410 3450
rect 4070 3308 4138 3364
rect 4194 3308 4280 3364
rect 4336 3308 4410 3364
rect 4070 3222 4410 3308
rect 4070 3166 4138 3222
rect 4194 3166 4280 3222
rect 4336 3166 4410 3222
rect 4070 3080 4410 3166
rect 4070 3024 4138 3080
rect 4194 3024 4280 3080
rect 4336 3024 4410 3080
rect 4070 2938 4410 3024
rect 4070 2882 4138 2938
rect 4194 2882 4280 2938
rect 4336 2882 4410 2938
rect 4070 2796 4410 2882
rect 4070 2740 4138 2796
rect 4194 2740 4280 2796
rect 4336 2740 4410 2796
rect 4070 2654 4410 2740
rect 4070 2598 4138 2654
rect 4194 2598 4280 2654
rect 4336 2598 4410 2654
rect 4070 2512 4410 2598
rect 4070 2456 4138 2512
rect 4194 2456 4280 2512
rect 4336 2456 4410 2512
rect 4070 2370 4410 2456
rect 4070 2314 4138 2370
rect 4194 2314 4280 2370
rect 4336 2314 4410 2370
rect 4070 2228 4410 2314
rect 4070 2172 4138 2228
rect 4194 2172 4280 2228
rect 4336 2172 4410 2228
rect 4070 2086 4410 2172
rect 4070 2030 4138 2086
rect 4194 2030 4280 2086
rect 4336 2030 4410 2086
rect 4070 1944 4410 2030
rect 4070 1888 4138 1944
rect 4194 1888 4280 1944
rect 4336 1888 4410 1944
rect 4070 1802 4410 1888
rect 4070 1746 4138 1802
rect 4194 1746 4280 1802
rect 4336 1746 4410 1802
rect 4070 1660 4410 1746
rect 4070 1604 4138 1660
rect 4194 1604 4280 1660
rect 4336 1604 4410 1660
rect 4070 1518 4410 1604
rect 4070 1462 4138 1518
rect 4194 1462 4280 1518
rect 4336 1462 4410 1518
rect 4070 1376 4410 1462
rect 4070 1320 4138 1376
rect 4194 1320 4280 1376
rect 4336 1320 4410 1376
rect 4070 1234 4410 1320
rect 4070 1178 4138 1234
rect 4194 1178 4280 1234
rect 4336 1178 4410 1234
rect 4070 1092 4410 1178
rect 4070 1036 4138 1092
rect 4194 1036 4280 1092
rect 4336 1036 4410 1092
rect 4070 950 4410 1036
rect 4070 894 4138 950
rect 4194 894 4280 950
rect 4336 894 4410 950
rect 4070 808 4410 894
rect 4070 752 4138 808
rect 4194 752 4280 808
rect 4336 752 4410 808
rect 4070 666 4410 752
rect 4070 610 4138 666
rect 4194 610 4280 666
rect 4336 610 4410 666
rect 4070 524 4410 610
rect 4070 468 4138 524
rect 4194 468 4280 524
rect 4336 468 4410 524
rect 4070 458 4410 468
rect 4610 12310 4950 12320
rect 4610 12254 4678 12310
rect 4734 12254 4820 12310
rect 4876 12254 4950 12310
rect 4610 12168 4950 12254
rect 4610 12112 4678 12168
rect 4734 12112 4820 12168
rect 4876 12112 4950 12168
rect 4610 12026 4950 12112
rect 4610 11970 4678 12026
rect 4734 11970 4820 12026
rect 4876 11970 4950 12026
rect 4610 11884 4950 11970
rect 4610 11828 4678 11884
rect 4734 11828 4820 11884
rect 4876 11828 4950 11884
rect 4610 11742 4950 11828
rect 4610 11686 4678 11742
rect 4734 11686 4820 11742
rect 4876 11686 4950 11742
rect 4610 11600 4950 11686
rect 4610 11544 4678 11600
rect 4734 11544 4820 11600
rect 4876 11544 4950 11600
rect 4610 11458 4950 11544
rect 4610 11402 4678 11458
rect 4734 11402 4820 11458
rect 4876 11402 4950 11458
rect 4610 11316 4950 11402
rect 4610 11260 4678 11316
rect 4734 11260 4820 11316
rect 4876 11260 4950 11316
rect 4610 11174 4950 11260
rect 4610 11118 4678 11174
rect 4734 11118 4820 11174
rect 4876 11118 4950 11174
rect 4610 11032 4950 11118
rect 4610 10976 4678 11032
rect 4734 10976 4820 11032
rect 4876 10976 4950 11032
rect 4610 10890 4950 10976
rect 4610 10834 4678 10890
rect 4734 10834 4820 10890
rect 4876 10834 4950 10890
rect 4610 10748 4950 10834
rect 4610 10692 4678 10748
rect 4734 10692 4820 10748
rect 4876 10692 4950 10748
rect 4610 10606 4950 10692
rect 4610 10550 4678 10606
rect 4734 10550 4820 10606
rect 4876 10550 4950 10606
rect 4610 10464 4950 10550
rect 4610 10408 4678 10464
rect 4734 10408 4820 10464
rect 4876 10408 4950 10464
rect 4610 10322 4950 10408
rect 4610 10266 4678 10322
rect 4734 10266 4820 10322
rect 4876 10266 4950 10322
rect 4610 10180 4950 10266
rect 4610 10124 4678 10180
rect 4734 10124 4820 10180
rect 4876 10124 4950 10180
rect 4610 10038 4950 10124
rect 4610 9982 4678 10038
rect 4734 9982 4820 10038
rect 4876 9982 4950 10038
rect 4610 9896 4950 9982
rect 4610 9840 4678 9896
rect 4734 9840 4820 9896
rect 4876 9840 4950 9896
rect 4610 9754 4950 9840
rect 4610 9698 4678 9754
rect 4734 9698 4820 9754
rect 4876 9698 4950 9754
rect 4610 9612 4950 9698
rect 4610 9556 4678 9612
rect 4734 9556 4820 9612
rect 4876 9556 4950 9612
rect 4610 9470 4950 9556
rect 4610 9414 4678 9470
rect 4734 9414 4820 9470
rect 4876 9414 4950 9470
rect 4610 9328 4950 9414
rect 4610 9272 4678 9328
rect 4734 9272 4820 9328
rect 4876 9272 4950 9328
rect 4610 9186 4950 9272
rect 4610 9130 4678 9186
rect 4734 9130 4820 9186
rect 4876 9130 4950 9186
rect 4610 9044 4950 9130
rect 4610 8988 4678 9044
rect 4734 8988 4820 9044
rect 4876 8988 4950 9044
rect 4610 8902 4950 8988
rect 4610 8846 4678 8902
rect 4734 8846 4820 8902
rect 4876 8846 4950 8902
rect 4610 8760 4950 8846
rect 4610 8704 4678 8760
rect 4734 8704 4820 8760
rect 4876 8704 4950 8760
rect 4610 8618 4950 8704
rect 4610 8562 4678 8618
rect 4734 8562 4820 8618
rect 4876 8562 4950 8618
rect 4610 8476 4950 8562
rect 4610 8420 4678 8476
rect 4734 8420 4820 8476
rect 4876 8420 4950 8476
rect 4610 8334 4950 8420
rect 4610 8278 4678 8334
rect 4734 8278 4820 8334
rect 4876 8278 4950 8334
rect 4610 8192 4950 8278
rect 4610 8136 4678 8192
rect 4734 8136 4820 8192
rect 4876 8136 4950 8192
rect 4610 8050 4950 8136
rect 4610 7994 4678 8050
rect 4734 7994 4820 8050
rect 4876 7994 4950 8050
rect 4610 7908 4950 7994
rect 4610 7852 4678 7908
rect 4734 7852 4820 7908
rect 4876 7852 4950 7908
rect 4610 7766 4950 7852
rect 4610 7710 4678 7766
rect 4734 7710 4820 7766
rect 4876 7710 4950 7766
rect 4610 7624 4950 7710
rect 4610 7568 4678 7624
rect 4734 7568 4820 7624
rect 4876 7568 4950 7624
rect 4610 7482 4950 7568
rect 4610 7426 4678 7482
rect 4734 7426 4820 7482
rect 4876 7426 4950 7482
rect 4610 7340 4950 7426
rect 4610 7284 4678 7340
rect 4734 7284 4820 7340
rect 4876 7284 4950 7340
rect 4610 7198 4950 7284
rect 4610 7142 4678 7198
rect 4734 7142 4820 7198
rect 4876 7142 4950 7198
rect 4610 7056 4950 7142
rect 4610 7000 4678 7056
rect 4734 7000 4820 7056
rect 4876 7000 4950 7056
rect 4610 6914 4950 7000
rect 4610 6858 4678 6914
rect 4734 6858 4820 6914
rect 4876 6858 4950 6914
rect 4610 6772 4950 6858
rect 4610 6716 4678 6772
rect 4734 6716 4820 6772
rect 4876 6716 4950 6772
rect 4610 6630 4950 6716
rect 4610 6574 4678 6630
rect 4734 6574 4820 6630
rect 4876 6574 4950 6630
rect 4610 6488 4950 6574
rect 4610 6432 4678 6488
rect 4734 6432 4820 6488
rect 4876 6432 4950 6488
rect 4610 6346 4950 6432
rect 4610 6290 4678 6346
rect 4734 6290 4820 6346
rect 4876 6290 4950 6346
rect 4610 6204 4950 6290
rect 4610 6148 4678 6204
rect 4734 6148 4820 6204
rect 4876 6148 4950 6204
rect 4610 6062 4950 6148
rect 4610 6006 4678 6062
rect 4734 6006 4820 6062
rect 4876 6006 4950 6062
rect 4610 5920 4950 6006
rect 4610 5864 4678 5920
rect 4734 5864 4820 5920
rect 4876 5864 4950 5920
rect 4610 5778 4950 5864
rect 4610 5722 4678 5778
rect 4734 5722 4820 5778
rect 4876 5722 4950 5778
rect 4610 5636 4950 5722
rect 4610 5580 4678 5636
rect 4734 5580 4820 5636
rect 4876 5580 4950 5636
rect 4610 5494 4950 5580
rect 4610 5438 4678 5494
rect 4734 5438 4820 5494
rect 4876 5438 4950 5494
rect 4610 5352 4950 5438
rect 4610 5296 4678 5352
rect 4734 5296 4820 5352
rect 4876 5296 4950 5352
rect 4610 5210 4950 5296
rect 4610 5154 4678 5210
rect 4734 5154 4820 5210
rect 4876 5154 4950 5210
rect 4610 5068 4950 5154
rect 4610 5012 4678 5068
rect 4734 5012 4820 5068
rect 4876 5012 4950 5068
rect 4610 4926 4950 5012
rect 4610 4870 4678 4926
rect 4734 4870 4820 4926
rect 4876 4870 4950 4926
rect 4610 4784 4950 4870
rect 4610 4728 4678 4784
rect 4734 4728 4820 4784
rect 4876 4728 4950 4784
rect 4610 4642 4950 4728
rect 4610 4586 4678 4642
rect 4734 4586 4820 4642
rect 4876 4586 4950 4642
rect 4610 4500 4950 4586
rect 4610 4444 4678 4500
rect 4734 4444 4820 4500
rect 4876 4444 4950 4500
rect 4610 4358 4950 4444
rect 4610 4302 4678 4358
rect 4734 4302 4820 4358
rect 4876 4302 4950 4358
rect 4610 4216 4950 4302
rect 4610 4160 4678 4216
rect 4734 4160 4820 4216
rect 4876 4160 4950 4216
rect 4610 4074 4950 4160
rect 4610 4018 4678 4074
rect 4734 4018 4820 4074
rect 4876 4018 4950 4074
rect 4610 3932 4950 4018
rect 4610 3876 4678 3932
rect 4734 3876 4820 3932
rect 4876 3876 4950 3932
rect 4610 3790 4950 3876
rect 4610 3734 4678 3790
rect 4734 3734 4820 3790
rect 4876 3734 4950 3790
rect 4610 3648 4950 3734
rect 4610 3592 4678 3648
rect 4734 3592 4820 3648
rect 4876 3592 4950 3648
rect 4610 3506 4950 3592
rect 4610 3450 4678 3506
rect 4734 3450 4820 3506
rect 4876 3450 4950 3506
rect 4610 3364 4950 3450
rect 4610 3308 4678 3364
rect 4734 3308 4820 3364
rect 4876 3308 4950 3364
rect 4610 3222 4950 3308
rect 4610 3166 4678 3222
rect 4734 3166 4820 3222
rect 4876 3166 4950 3222
rect 4610 3080 4950 3166
rect 4610 3024 4678 3080
rect 4734 3024 4820 3080
rect 4876 3024 4950 3080
rect 4610 2938 4950 3024
rect 4610 2882 4678 2938
rect 4734 2882 4820 2938
rect 4876 2882 4950 2938
rect 4610 2796 4950 2882
rect 4610 2740 4678 2796
rect 4734 2740 4820 2796
rect 4876 2740 4950 2796
rect 4610 2654 4950 2740
rect 4610 2598 4678 2654
rect 4734 2598 4820 2654
rect 4876 2598 4950 2654
rect 4610 2512 4950 2598
rect 4610 2456 4678 2512
rect 4734 2456 4820 2512
rect 4876 2456 4950 2512
rect 4610 2370 4950 2456
rect 4610 2314 4678 2370
rect 4734 2314 4820 2370
rect 4876 2314 4950 2370
rect 4610 2228 4950 2314
rect 4610 2172 4678 2228
rect 4734 2172 4820 2228
rect 4876 2172 4950 2228
rect 4610 2086 4950 2172
rect 4610 2030 4678 2086
rect 4734 2030 4820 2086
rect 4876 2030 4950 2086
rect 4610 1944 4950 2030
rect 4610 1888 4678 1944
rect 4734 1888 4820 1944
rect 4876 1888 4950 1944
rect 4610 1802 4950 1888
rect 4610 1746 4678 1802
rect 4734 1746 4820 1802
rect 4876 1746 4950 1802
rect 4610 1660 4950 1746
rect 4610 1604 4678 1660
rect 4734 1604 4820 1660
rect 4876 1604 4950 1660
rect 4610 1518 4950 1604
rect 4610 1462 4678 1518
rect 4734 1462 4820 1518
rect 4876 1462 4950 1518
rect 4610 1376 4950 1462
rect 4610 1320 4678 1376
rect 4734 1320 4820 1376
rect 4876 1320 4950 1376
rect 4610 1234 4950 1320
rect 4610 1178 4678 1234
rect 4734 1178 4820 1234
rect 4876 1178 4950 1234
rect 4610 1092 4950 1178
rect 4610 1036 4678 1092
rect 4734 1036 4820 1092
rect 4876 1036 4950 1092
rect 4610 950 4950 1036
rect 4610 894 4678 950
rect 4734 894 4820 950
rect 4876 894 4950 950
rect 4610 808 4950 894
rect 4610 752 4678 808
rect 4734 752 4820 808
rect 4876 752 4950 808
rect 4610 666 4950 752
rect 4610 610 4678 666
rect 4734 610 4820 666
rect 4876 610 4950 666
rect 4610 524 4950 610
rect 4610 468 4678 524
rect 4734 468 4820 524
rect 4876 468 4950 524
rect 4610 458 4950 468
rect 5150 12310 5490 12320
rect 5150 12254 5215 12310
rect 5271 12254 5357 12310
rect 5413 12254 5490 12310
rect 5150 12168 5490 12254
rect 5150 12112 5215 12168
rect 5271 12112 5357 12168
rect 5413 12112 5490 12168
rect 5150 12026 5490 12112
rect 5150 11970 5215 12026
rect 5271 11970 5357 12026
rect 5413 11970 5490 12026
rect 5150 11884 5490 11970
rect 5150 11828 5215 11884
rect 5271 11828 5357 11884
rect 5413 11828 5490 11884
rect 5150 11742 5490 11828
rect 5150 11686 5215 11742
rect 5271 11686 5357 11742
rect 5413 11686 5490 11742
rect 5150 11600 5490 11686
rect 5150 11544 5215 11600
rect 5271 11544 5357 11600
rect 5413 11544 5490 11600
rect 5150 11458 5490 11544
rect 5150 11402 5215 11458
rect 5271 11402 5357 11458
rect 5413 11402 5490 11458
rect 5150 11316 5490 11402
rect 5150 11260 5215 11316
rect 5271 11260 5357 11316
rect 5413 11260 5490 11316
rect 5150 11174 5490 11260
rect 5150 11118 5215 11174
rect 5271 11118 5357 11174
rect 5413 11118 5490 11174
rect 5150 11032 5490 11118
rect 5150 10976 5215 11032
rect 5271 10976 5357 11032
rect 5413 10976 5490 11032
rect 5150 10890 5490 10976
rect 5150 10834 5215 10890
rect 5271 10834 5357 10890
rect 5413 10834 5490 10890
rect 5150 10748 5490 10834
rect 5150 10692 5215 10748
rect 5271 10692 5357 10748
rect 5413 10692 5490 10748
rect 5150 10606 5490 10692
rect 5150 10550 5215 10606
rect 5271 10550 5357 10606
rect 5413 10550 5490 10606
rect 5150 10464 5490 10550
rect 5150 10408 5215 10464
rect 5271 10408 5357 10464
rect 5413 10408 5490 10464
rect 5150 10322 5490 10408
rect 5150 10266 5215 10322
rect 5271 10266 5357 10322
rect 5413 10266 5490 10322
rect 5150 10180 5490 10266
rect 5150 10124 5215 10180
rect 5271 10124 5357 10180
rect 5413 10124 5490 10180
rect 5150 10038 5490 10124
rect 5150 9982 5215 10038
rect 5271 9982 5357 10038
rect 5413 9982 5490 10038
rect 5150 9896 5490 9982
rect 5150 9840 5215 9896
rect 5271 9840 5357 9896
rect 5413 9840 5490 9896
rect 5150 9754 5490 9840
rect 5150 9698 5215 9754
rect 5271 9698 5357 9754
rect 5413 9698 5490 9754
rect 5150 9612 5490 9698
rect 5150 9556 5215 9612
rect 5271 9556 5357 9612
rect 5413 9556 5490 9612
rect 5150 9470 5490 9556
rect 5150 9414 5215 9470
rect 5271 9414 5357 9470
rect 5413 9414 5490 9470
rect 5150 9328 5490 9414
rect 5150 9272 5215 9328
rect 5271 9272 5357 9328
rect 5413 9272 5490 9328
rect 5150 9186 5490 9272
rect 5150 9130 5215 9186
rect 5271 9130 5357 9186
rect 5413 9130 5490 9186
rect 5150 9044 5490 9130
rect 5150 8988 5215 9044
rect 5271 8988 5357 9044
rect 5413 8988 5490 9044
rect 5150 8902 5490 8988
rect 5150 8846 5215 8902
rect 5271 8846 5357 8902
rect 5413 8846 5490 8902
rect 5150 8760 5490 8846
rect 5150 8704 5215 8760
rect 5271 8704 5357 8760
rect 5413 8704 5490 8760
rect 5150 8618 5490 8704
rect 5150 8562 5215 8618
rect 5271 8562 5357 8618
rect 5413 8562 5490 8618
rect 5150 8476 5490 8562
rect 5150 8420 5215 8476
rect 5271 8420 5357 8476
rect 5413 8420 5490 8476
rect 5150 8334 5490 8420
rect 5150 8278 5215 8334
rect 5271 8278 5357 8334
rect 5413 8278 5490 8334
rect 5150 8192 5490 8278
rect 5150 8136 5215 8192
rect 5271 8136 5357 8192
rect 5413 8136 5490 8192
rect 5150 8050 5490 8136
rect 5150 7994 5215 8050
rect 5271 7994 5357 8050
rect 5413 7994 5490 8050
rect 5150 7908 5490 7994
rect 5150 7852 5215 7908
rect 5271 7852 5357 7908
rect 5413 7852 5490 7908
rect 5150 7766 5490 7852
rect 5150 7710 5215 7766
rect 5271 7710 5357 7766
rect 5413 7710 5490 7766
rect 5150 7624 5490 7710
rect 5150 7568 5215 7624
rect 5271 7568 5357 7624
rect 5413 7568 5490 7624
rect 5150 7482 5490 7568
rect 5150 7426 5215 7482
rect 5271 7426 5357 7482
rect 5413 7426 5490 7482
rect 5150 7340 5490 7426
rect 5150 7284 5215 7340
rect 5271 7284 5357 7340
rect 5413 7284 5490 7340
rect 5150 7198 5490 7284
rect 5150 7142 5215 7198
rect 5271 7142 5357 7198
rect 5413 7142 5490 7198
rect 5150 7056 5490 7142
rect 5150 7000 5215 7056
rect 5271 7000 5357 7056
rect 5413 7000 5490 7056
rect 5150 6914 5490 7000
rect 5150 6858 5215 6914
rect 5271 6858 5357 6914
rect 5413 6858 5490 6914
rect 5150 6772 5490 6858
rect 5150 6716 5215 6772
rect 5271 6716 5357 6772
rect 5413 6716 5490 6772
rect 5150 6630 5490 6716
rect 5150 6574 5215 6630
rect 5271 6574 5357 6630
rect 5413 6574 5490 6630
rect 5150 6488 5490 6574
rect 5150 6432 5215 6488
rect 5271 6432 5357 6488
rect 5413 6432 5490 6488
rect 5150 6346 5490 6432
rect 5150 6290 5215 6346
rect 5271 6290 5357 6346
rect 5413 6290 5490 6346
rect 5150 6204 5490 6290
rect 5150 6148 5215 6204
rect 5271 6148 5357 6204
rect 5413 6148 5490 6204
rect 5150 6062 5490 6148
rect 5150 6006 5215 6062
rect 5271 6006 5357 6062
rect 5413 6006 5490 6062
rect 5150 5920 5490 6006
rect 5150 5864 5215 5920
rect 5271 5864 5357 5920
rect 5413 5864 5490 5920
rect 5150 5778 5490 5864
rect 5150 5722 5215 5778
rect 5271 5722 5357 5778
rect 5413 5722 5490 5778
rect 5150 5636 5490 5722
rect 5150 5580 5215 5636
rect 5271 5580 5357 5636
rect 5413 5580 5490 5636
rect 5150 5494 5490 5580
rect 5150 5438 5215 5494
rect 5271 5438 5357 5494
rect 5413 5438 5490 5494
rect 5150 5352 5490 5438
rect 5150 5296 5215 5352
rect 5271 5296 5357 5352
rect 5413 5296 5490 5352
rect 5150 5210 5490 5296
rect 5150 5154 5215 5210
rect 5271 5154 5357 5210
rect 5413 5154 5490 5210
rect 5150 5068 5490 5154
rect 5150 5012 5215 5068
rect 5271 5012 5357 5068
rect 5413 5012 5490 5068
rect 5150 4926 5490 5012
rect 5150 4870 5215 4926
rect 5271 4870 5357 4926
rect 5413 4870 5490 4926
rect 5150 4784 5490 4870
rect 5150 4728 5215 4784
rect 5271 4728 5357 4784
rect 5413 4728 5490 4784
rect 5150 4642 5490 4728
rect 5150 4586 5215 4642
rect 5271 4586 5357 4642
rect 5413 4586 5490 4642
rect 5150 4500 5490 4586
rect 5150 4444 5215 4500
rect 5271 4444 5357 4500
rect 5413 4444 5490 4500
rect 5150 4358 5490 4444
rect 5150 4302 5215 4358
rect 5271 4302 5357 4358
rect 5413 4302 5490 4358
rect 5150 4216 5490 4302
rect 5150 4160 5215 4216
rect 5271 4160 5357 4216
rect 5413 4160 5490 4216
rect 5150 4074 5490 4160
rect 5150 4018 5215 4074
rect 5271 4018 5357 4074
rect 5413 4018 5490 4074
rect 5150 3932 5490 4018
rect 5150 3876 5215 3932
rect 5271 3876 5357 3932
rect 5413 3876 5490 3932
rect 5150 3790 5490 3876
rect 5150 3734 5215 3790
rect 5271 3734 5357 3790
rect 5413 3734 5490 3790
rect 5150 3648 5490 3734
rect 5150 3592 5215 3648
rect 5271 3592 5357 3648
rect 5413 3592 5490 3648
rect 5150 3506 5490 3592
rect 5150 3450 5215 3506
rect 5271 3450 5357 3506
rect 5413 3450 5490 3506
rect 5150 3364 5490 3450
rect 5150 3308 5215 3364
rect 5271 3308 5357 3364
rect 5413 3308 5490 3364
rect 5150 3222 5490 3308
rect 5150 3166 5215 3222
rect 5271 3166 5357 3222
rect 5413 3166 5490 3222
rect 5150 3080 5490 3166
rect 5150 3024 5215 3080
rect 5271 3024 5357 3080
rect 5413 3024 5490 3080
rect 5150 2938 5490 3024
rect 5150 2882 5215 2938
rect 5271 2882 5357 2938
rect 5413 2882 5490 2938
rect 5150 2796 5490 2882
rect 5150 2740 5215 2796
rect 5271 2740 5357 2796
rect 5413 2740 5490 2796
rect 5150 2654 5490 2740
rect 5150 2598 5215 2654
rect 5271 2598 5357 2654
rect 5413 2598 5490 2654
rect 5150 2512 5490 2598
rect 5150 2456 5215 2512
rect 5271 2456 5357 2512
rect 5413 2456 5490 2512
rect 5150 2370 5490 2456
rect 5150 2314 5215 2370
rect 5271 2314 5357 2370
rect 5413 2314 5490 2370
rect 5150 2228 5490 2314
rect 5150 2172 5215 2228
rect 5271 2172 5357 2228
rect 5413 2172 5490 2228
rect 5150 2086 5490 2172
rect 5150 2030 5215 2086
rect 5271 2030 5357 2086
rect 5413 2030 5490 2086
rect 5150 1944 5490 2030
rect 5150 1888 5215 1944
rect 5271 1888 5357 1944
rect 5413 1888 5490 1944
rect 5150 1802 5490 1888
rect 5150 1746 5215 1802
rect 5271 1746 5357 1802
rect 5413 1746 5490 1802
rect 5150 1660 5490 1746
rect 5150 1604 5215 1660
rect 5271 1604 5357 1660
rect 5413 1604 5490 1660
rect 5150 1518 5490 1604
rect 5150 1462 5215 1518
rect 5271 1462 5357 1518
rect 5413 1462 5490 1518
rect 5150 1376 5490 1462
rect 5150 1320 5215 1376
rect 5271 1320 5357 1376
rect 5413 1320 5490 1376
rect 5150 1234 5490 1320
rect 5150 1178 5215 1234
rect 5271 1178 5357 1234
rect 5413 1178 5490 1234
rect 5150 1092 5490 1178
rect 5150 1036 5215 1092
rect 5271 1036 5357 1092
rect 5413 1036 5490 1092
rect 5150 950 5490 1036
rect 5150 894 5215 950
rect 5271 894 5357 950
rect 5413 894 5490 950
rect 5150 808 5490 894
rect 5150 752 5215 808
rect 5271 752 5357 808
rect 5413 752 5490 808
rect 5150 666 5490 752
rect 5150 610 5215 666
rect 5271 610 5357 666
rect 5413 610 5490 666
rect 5150 524 5490 610
rect 5150 468 5215 524
rect 5271 468 5357 524
rect 5413 468 5490 524
rect 5150 458 5490 468
rect 5690 12310 6030 12320
rect 5690 12254 5760 12310
rect 5816 12254 5902 12310
rect 5958 12254 6030 12310
rect 5690 12168 6030 12254
rect 5690 12112 5760 12168
rect 5816 12112 5902 12168
rect 5958 12112 6030 12168
rect 5690 12026 6030 12112
rect 5690 11970 5760 12026
rect 5816 11970 5902 12026
rect 5958 11970 6030 12026
rect 5690 11884 6030 11970
rect 5690 11828 5760 11884
rect 5816 11828 5902 11884
rect 5958 11828 6030 11884
rect 5690 11742 6030 11828
rect 5690 11686 5760 11742
rect 5816 11686 5902 11742
rect 5958 11686 6030 11742
rect 5690 11600 6030 11686
rect 5690 11544 5760 11600
rect 5816 11544 5902 11600
rect 5958 11544 6030 11600
rect 5690 11458 6030 11544
rect 5690 11402 5760 11458
rect 5816 11402 5902 11458
rect 5958 11402 6030 11458
rect 5690 11316 6030 11402
rect 5690 11260 5760 11316
rect 5816 11260 5902 11316
rect 5958 11260 6030 11316
rect 5690 11174 6030 11260
rect 5690 11118 5760 11174
rect 5816 11118 5902 11174
rect 5958 11118 6030 11174
rect 5690 11032 6030 11118
rect 5690 10976 5760 11032
rect 5816 10976 5902 11032
rect 5958 10976 6030 11032
rect 5690 10890 6030 10976
rect 5690 10834 5760 10890
rect 5816 10834 5902 10890
rect 5958 10834 6030 10890
rect 5690 10748 6030 10834
rect 5690 10692 5760 10748
rect 5816 10692 5902 10748
rect 5958 10692 6030 10748
rect 5690 10606 6030 10692
rect 5690 10550 5760 10606
rect 5816 10550 5902 10606
rect 5958 10550 6030 10606
rect 5690 10464 6030 10550
rect 5690 10408 5760 10464
rect 5816 10408 5902 10464
rect 5958 10408 6030 10464
rect 5690 10322 6030 10408
rect 5690 10266 5760 10322
rect 5816 10266 5902 10322
rect 5958 10266 6030 10322
rect 5690 10180 6030 10266
rect 5690 10124 5760 10180
rect 5816 10124 5902 10180
rect 5958 10124 6030 10180
rect 5690 10038 6030 10124
rect 5690 9982 5760 10038
rect 5816 9982 5902 10038
rect 5958 9982 6030 10038
rect 5690 9896 6030 9982
rect 5690 9840 5760 9896
rect 5816 9840 5902 9896
rect 5958 9840 6030 9896
rect 5690 9754 6030 9840
rect 5690 9698 5760 9754
rect 5816 9698 5902 9754
rect 5958 9698 6030 9754
rect 5690 9612 6030 9698
rect 5690 9556 5760 9612
rect 5816 9556 5902 9612
rect 5958 9556 6030 9612
rect 5690 9470 6030 9556
rect 5690 9414 5760 9470
rect 5816 9414 5902 9470
rect 5958 9414 6030 9470
rect 5690 9328 6030 9414
rect 5690 9272 5760 9328
rect 5816 9272 5902 9328
rect 5958 9272 6030 9328
rect 5690 9186 6030 9272
rect 5690 9130 5760 9186
rect 5816 9130 5902 9186
rect 5958 9130 6030 9186
rect 5690 9044 6030 9130
rect 5690 8988 5760 9044
rect 5816 8988 5902 9044
rect 5958 8988 6030 9044
rect 5690 8902 6030 8988
rect 5690 8846 5760 8902
rect 5816 8846 5902 8902
rect 5958 8846 6030 8902
rect 5690 8760 6030 8846
rect 5690 8704 5760 8760
rect 5816 8704 5902 8760
rect 5958 8704 6030 8760
rect 5690 8618 6030 8704
rect 5690 8562 5760 8618
rect 5816 8562 5902 8618
rect 5958 8562 6030 8618
rect 5690 8476 6030 8562
rect 5690 8420 5760 8476
rect 5816 8420 5902 8476
rect 5958 8420 6030 8476
rect 5690 8334 6030 8420
rect 5690 8278 5760 8334
rect 5816 8278 5902 8334
rect 5958 8278 6030 8334
rect 5690 8192 6030 8278
rect 5690 8136 5760 8192
rect 5816 8136 5902 8192
rect 5958 8136 6030 8192
rect 5690 8050 6030 8136
rect 5690 7994 5760 8050
rect 5816 7994 5902 8050
rect 5958 7994 6030 8050
rect 5690 7908 6030 7994
rect 5690 7852 5760 7908
rect 5816 7852 5902 7908
rect 5958 7852 6030 7908
rect 5690 7766 6030 7852
rect 5690 7710 5760 7766
rect 5816 7710 5902 7766
rect 5958 7710 6030 7766
rect 5690 7624 6030 7710
rect 5690 7568 5760 7624
rect 5816 7568 5902 7624
rect 5958 7568 6030 7624
rect 5690 7482 6030 7568
rect 5690 7426 5760 7482
rect 5816 7426 5902 7482
rect 5958 7426 6030 7482
rect 5690 7340 6030 7426
rect 5690 7284 5760 7340
rect 5816 7284 5902 7340
rect 5958 7284 6030 7340
rect 5690 7198 6030 7284
rect 5690 7142 5760 7198
rect 5816 7142 5902 7198
rect 5958 7142 6030 7198
rect 5690 7056 6030 7142
rect 5690 7000 5760 7056
rect 5816 7000 5902 7056
rect 5958 7000 6030 7056
rect 5690 6914 6030 7000
rect 5690 6858 5760 6914
rect 5816 6858 5902 6914
rect 5958 6858 6030 6914
rect 5690 6772 6030 6858
rect 5690 6716 5760 6772
rect 5816 6716 5902 6772
rect 5958 6716 6030 6772
rect 5690 6630 6030 6716
rect 5690 6574 5760 6630
rect 5816 6574 5902 6630
rect 5958 6574 6030 6630
rect 5690 6488 6030 6574
rect 5690 6432 5760 6488
rect 5816 6432 5902 6488
rect 5958 6432 6030 6488
rect 5690 6346 6030 6432
rect 5690 6290 5760 6346
rect 5816 6290 5902 6346
rect 5958 6290 6030 6346
rect 5690 6204 6030 6290
rect 5690 6148 5760 6204
rect 5816 6148 5902 6204
rect 5958 6148 6030 6204
rect 5690 6062 6030 6148
rect 5690 6006 5760 6062
rect 5816 6006 5902 6062
rect 5958 6006 6030 6062
rect 5690 5920 6030 6006
rect 5690 5864 5760 5920
rect 5816 5864 5902 5920
rect 5958 5864 6030 5920
rect 5690 5778 6030 5864
rect 5690 5722 5760 5778
rect 5816 5722 5902 5778
rect 5958 5722 6030 5778
rect 5690 5636 6030 5722
rect 5690 5580 5760 5636
rect 5816 5580 5902 5636
rect 5958 5580 6030 5636
rect 5690 5494 6030 5580
rect 5690 5438 5760 5494
rect 5816 5438 5902 5494
rect 5958 5438 6030 5494
rect 5690 5352 6030 5438
rect 5690 5296 5760 5352
rect 5816 5296 5902 5352
rect 5958 5296 6030 5352
rect 5690 5210 6030 5296
rect 5690 5154 5760 5210
rect 5816 5154 5902 5210
rect 5958 5154 6030 5210
rect 5690 5068 6030 5154
rect 5690 5012 5760 5068
rect 5816 5012 5902 5068
rect 5958 5012 6030 5068
rect 5690 4926 6030 5012
rect 5690 4870 5760 4926
rect 5816 4870 5902 4926
rect 5958 4870 6030 4926
rect 5690 4784 6030 4870
rect 5690 4728 5760 4784
rect 5816 4728 5902 4784
rect 5958 4728 6030 4784
rect 5690 4642 6030 4728
rect 5690 4586 5760 4642
rect 5816 4586 5902 4642
rect 5958 4586 6030 4642
rect 5690 4500 6030 4586
rect 5690 4444 5760 4500
rect 5816 4444 5902 4500
rect 5958 4444 6030 4500
rect 5690 4358 6030 4444
rect 5690 4302 5760 4358
rect 5816 4302 5902 4358
rect 5958 4302 6030 4358
rect 5690 4216 6030 4302
rect 5690 4160 5760 4216
rect 5816 4160 5902 4216
rect 5958 4160 6030 4216
rect 5690 4074 6030 4160
rect 5690 4018 5760 4074
rect 5816 4018 5902 4074
rect 5958 4018 6030 4074
rect 5690 3932 6030 4018
rect 5690 3876 5760 3932
rect 5816 3876 5902 3932
rect 5958 3876 6030 3932
rect 5690 3790 6030 3876
rect 5690 3734 5760 3790
rect 5816 3734 5902 3790
rect 5958 3734 6030 3790
rect 5690 3648 6030 3734
rect 5690 3592 5760 3648
rect 5816 3592 5902 3648
rect 5958 3592 6030 3648
rect 5690 3506 6030 3592
rect 5690 3450 5760 3506
rect 5816 3450 5902 3506
rect 5958 3450 6030 3506
rect 5690 3364 6030 3450
rect 5690 3308 5760 3364
rect 5816 3308 5902 3364
rect 5958 3308 6030 3364
rect 5690 3222 6030 3308
rect 5690 3166 5760 3222
rect 5816 3166 5902 3222
rect 5958 3166 6030 3222
rect 5690 3080 6030 3166
rect 5690 3024 5760 3080
rect 5816 3024 5902 3080
rect 5958 3024 6030 3080
rect 5690 2938 6030 3024
rect 5690 2882 5760 2938
rect 5816 2882 5902 2938
rect 5958 2882 6030 2938
rect 5690 2796 6030 2882
rect 5690 2740 5760 2796
rect 5816 2740 5902 2796
rect 5958 2740 6030 2796
rect 5690 2654 6030 2740
rect 5690 2598 5760 2654
rect 5816 2598 5902 2654
rect 5958 2598 6030 2654
rect 5690 2512 6030 2598
rect 5690 2456 5760 2512
rect 5816 2456 5902 2512
rect 5958 2456 6030 2512
rect 5690 2370 6030 2456
rect 5690 2314 5760 2370
rect 5816 2314 5902 2370
rect 5958 2314 6030 2370
rect 5690 2228 6030 2314
rect 5690 2172 5760 2228
rect 5816 2172 5902 2228
rect 5958 2172 6030 2228
rect 5690 2086 6030 2172
rect 5690 2030 5760 2086
rect 5816 2030 5902 2086
rect 5958 2030 6030 2086
rect 5690 1944 6030 2030
rect 5690 1888 5760 1944
rect 5816 1888 5902 1944
rect 5958 1888 6030 1944
rect 5690 1802 6030 1888
rect 5690 1746 5760 1802
rect 5816 1746 5902 1802
rect 5958 1746 6030 1802
rect 5690 1660 6030 1746
rect 5690 1604 5760 1660
rect 5816 1604 5902 1660
rect 5958 1604 6030 1660
rect 5690 1518 6030 1604
rect 5690 1462 5760 1518
rect 5816 1462 5902 1518
rect 5958 1462 6030 1518
rect 5690 1376 6030 1462
rect 5690 1320 5760 1376
rect 5816 1320 5902 1376
rect 5958 1320 6030 1376
rect 5690 1234 6030 1320
rect 5690 1178 5760 1234
rect 5816 1178 5902 1234
rect 5958 1178 6030 1234
rect 5690 1092 6030 1178
rect 5690 1036 5760 1092
rect 5816 1036 5902 1092
rect 5958 1036 6030 1092
rect 5690 950 6030 1036
rect 5690 894 5760 950
rect 5816 894 5902 950
rect 5958 894 6030 950
rect 5690 808 6030 894
rect 5690 752 5760 808
rect 5816 752 5902 808
rect 5958 752 6030 808
rect 5690 666 6030 752
rect 5690 610 5760 666
rect 5816 610 5902 666
rect 5958 610 6030 666
rect 5690 524 6030 610
rect 5690 468 5760 524
rect 5816 468 5902 524
rect 5958 468 6030 524
rect 5690 458 6030 468
rect 6230 12310 6570 12320
rect 6230 12254 6300 12310
rect 6356 12254 6442 12310
rect 6498 12254 6570 12310
rect 6230 12168 6570 12254
rect 6230 12112 6300 12168
rect 6356 12112 6442 12168
rect 6498 12112 6570 12168
rect 6230 12026 6570 12112
rect 6230 11970 6300 12026
rect 6356 11970 6442 12026
rect 6498 11970 6570 12026
rect 6230 11884 6570 11970
rect 6230 11828 6300 11884
rect 6356 11828 6442 11884
rect 6498 11828 6570 11884
rect 6230 11742 6570 11828
rect 6230 11686 6300 11742
rect 6356 11686 6442 11742
rect 6498 11686 6570 11742
rect 6230 11600 6570 11686
rect 6230 11544 6300 11600
rect 6356 11544 6442 11600
rect 6498 11544 6570 11600
rect 6230 11458 6570 11544
rect 6230 11402 6300 11458
rect 6356 11402 6442 11458
rect 6498 11402 6570 11458
rect 6230 11316 6570 11402
rect 6230 11260 6300 11316
rect 6356 11260 6442 11316
rect 6498 11260 6570 11316
rect 6230 11174 6570 11260
rect 6230 11118 6300 11174
rect 6356 11118 6442 11174
rect 6498 11118 6570 11174
rect 6230 11032 6570 11118
rect 6230 10976 6300 11032
rect 6356 10976 6442 11032
rect 6498 10976 6570 11032
rect 6230 10890 6570 10976
rect 6230 10834 6300 10890
rect 6356 10834 6442 10890
rect 6498 10834 6570 10890
rect 6230 10748 6570 10834
rect 6230 10692 6300 10748
rect 6356 10692 6442 10748
rect 6498 10692 6570 10748
rect 6230 10606 6570 10692
rect 6230 10550 6300 10606
rect 6356 10550 6442 10606
rect 6498 10550 6570 10606
rect 6230 10464 6570 10550
rect 6230 10408 6300 10464
rect 6356 10408 6442 10464
rect 6498 10408 6570 10464
rect 6230 10322 6570 10408
rect 6230 10266 6300 10322
rect 6356 10266 6442 10322
rect 6498 10266 6570 10322
rect 6230 10180 6570 10266
rect 6230 10124 6300 10180
rect 6356 10124 6442 10180
rect 6498 10124 6570 10180
rect 6230 10038 6570 10124
rect 6230 9982 6300 10038
rect 6356 9982 6442 10038
rect 6498 9982 6570 10038
rect 6230 9896 6570 9982
rect 6230 9840 6300 9896
rect 6356 9840 6442 9896
rect 6498 9840 6570 9896
rect 6230 9754 6570 9840
rect 6230 9698 6300 9754
rect 6356 9698 6442 9754
rect 6498 9698 6570 9754
rect 6230 9612 6570 9698
rect 6230 9556 6300 9612
rect 6356 9556 6442 9612
rect 6498 9556 6570 9612
rect 6230 9470 6570 9556
rect 6230 9414 6300 9470
rect 6356 9414 6442 9470
rect 6498 9414 6570 9470
rect 6230 9328 6570 9414
rect 6230 9272 6300 9328
rect 6356 9272 6442 9328
rect 6498 9272 6570 9328
rect 6230 9186 6570 9272
rect 6230 9130 6300 9186
rect 6356 9130 6442 9186
rect 6498 9130 6570 9186
rect 6230 9044 6570 9130
rect 6230 8988 6300 9044
rect 6356 8988 6442 9044
rect 6498 8988 6570 9044
rect 6230 8902 6570 8988
rect 6230 8846 6300 8902
rect 6356 8846 6442 8902
rect 6498 8846 6570 8902
rect 6230 8760 6570 8846
rect 6230 8704 6300 8760
rect 6356 8704 6442 8760
rect 6498 8704 6570 8760
rect 6230 8618 6570 8704
rect 6230 8562 6300 8618
rect 6356 8562 6442 8618
rect 6498 8562 6570 8618
rect 6230 8476 6570 8562
rect 6230 8420 6300 8476
rect 6356 8420 6442 8476
rect 6498 8420 6570 8476
rect 6230 8334 6570 8420
rect 6230 8278 6300 8334
rect 6356 8278 6442 8334
rect 6498 8278 6570 8334
rect 6230 8192 6570 8278
rect 6230 8136 6300 8192
rect 6356 8136 6442 8192
rect 6498 8136 6570 8192
rect 6230 8050 6570 8136
rect 6230 7994 6300 8050
rect 6356 7994 6442 8050
rect 6498 7994 6570 8050
rect 6230 7908 6570 7994
rect 6230 7852 6300 7908
rect 6356 7852 6442 7908
rect 6498 7852 6570 7908
rect 6230 7766 6570 7852
rect 6230 7710 6300 7766
rect 6356 7710 6442 7766
rect 6498 7710 6570 7766
rect 6230 7624 6570 7710
rect 6230 7568 6300 7624
rect 6356 7568 6442 7624
rect 6498 7568 6570 7624
rect 6230 7482 6570 7568
rect 6230 7426 6300 7482
rect 6356 7426 6442 7482
rect 6498 7426 6570 7482
rect 6230 7340 6570 7426
rect 6230 7284 6300 7340
rect 6356 7284 6442 7340
rect 6498 7284 6570 7340
rect 6230 7198 6570 7284
rect 6230 7142 6300 7198
rect 6356 7142 6442 7198
rect 6498 7142 6570 7198
rect 6230 7056 6570 7142
rect 6230 7000 6300 7056
rect 6356 7000 6442 7056
rect 6498 7000 6570 7056
rect 6230 6914 6570 7000
rect 6230 6858 6300 6914
rect 6356 6858 6442 6914
rect 6498 6858 6570 6914
rect 6230 6772 6570 6858
rect 6230 6716 6300 6772
rect 6356 6716 6442 6772
rect 6498 6716 6570 6772
rect 6230 6630 6570 6716
rect 6230 6574 6300 6630
rect 6356 6574 6442 6630
rect 6498 6574 6570 6630
rect 6230 6488 6570 6574
rect 6230 6432 6300 6488
rect 6356 6432 6442 6488
rect 6498 6432 6570 6488
rect 6230 6346 6570 6432
rect 6230 6290 6300 6346
rect 6356 6290 6442 6346
rect 6498 6290 6570 6346
rect 6230 6204 6570 6290
rect 6230 6148 6300 6204
rect 6356 6148 6442 6204
rect 6498 6148 6570 6204
rect 6230 6062 6570 6148
rect 6230 6006 6300 6062
rect 6356 6006 6442 6062
rect 6498 6006 6570 6062
rect 6230 5920 6570 6006
rect 6230 5864 6300 5920
rect 6356 5864 6442 5920
rect 6498 5864 6570 5920
rect 6230 5778 6570 5864
rect 6230 5722 6300 5778
rect 6356 5722 6442 5778
rect 6498 5722 6570 5778
rect 6230 5636 6570 5722
rect 6230 5580 6300 5636
rect 6356 5580 6442 5636
rect 6498 5580 6570 5636
rect 6230 5494 6570 5580
rect 6230 5438 6300 5494
rect 6356 5438 6442 5494
rect 6498 5438 6570 5494
rect 6230 5352 6570 5438
rect 6230 5296 6300 5352
rect 6356 5296 6442 5352
rect 6498 5296 6570 5352
rect 6230 5210 6570 5296
rect 6230 5154 6300 5210
rect 6356 5154 6442 5210
rect 6498 5154 6570 5210
rect 6230 5068 6570 5154
rect 6230 5012 6300 5068
rect 6356 5012 6442 5068
rect 6498 5012 6570 5068
rect 6230 4926 6570 5012
rect 6230 4870 6300 4926
rect 6356 4870 6442 4926
rect 6498 4870 6570 4926
rect 6230 4784 6570 4870
rect 6230 4728 6300 4784
rect 6356 4728 6442 4784
rect 6498 4728 6570 4784
rect 6230 4642 6570 4728
rect 6230 4586 6300 4642
rect 6356 4586 6442 4642
rect 6498 4586 6570 4642
rect 6230 4500 6570 4586
rect 6230 4444 6300 4500
rect 6356 4444 6442 4500
rect 6498 4444 6570 4500
rect 6230 4358 6570 4444
rect 6230 4302 6300 4358
rect 6356 4302 6442 4358
rect 6498 4302 6570 4358
rect 6230 4216 6570 4302
rect 6230 4160 6300 4216
rect 6356 4160 6442 4216
rect 6498 4160 6570 4216
rect 6230 4074 6570 4160
rect 6230 4018 6300 4074
rect 6356 4018 6442 4074
rect 6498 4018 6570 4074
rect 6230 3932 6570 4018
rect 6230 3876 6300 3932
rect 6356 3876 6442 3932
rect 6498 3876 6570 3932
rect 6230 3790 6570 3876
rect 6230 3734 6300 3790
rect 6356 3734 6442 3790
rect 6498 3734 6570 3790
rect 6230 3648 6570 3734
rect 6230 3592 6300 3648
rect 6356 3592 6442 3648
rect 6498 3592 6570 3648
rect 6230 3506 6570 3592
rect 6230 3450 6300 3506
rect 6356 3450 6442 3506
rect 6498 3450 6570 3506
rect 6230 3364 6570 3450
rect 6230 3308 6300 3364
rect 6356 3308 6442 3364
rect 6498 3308 6570 3364
rect 6230 3222 6570 3308
rect 6230 3166 6300 3222
rect 6356 3166 6442 3222
rect 6498 3166 6570 3222
rect 6230 3080 6570 3166
rect 6230 3024 6300 3080
rect 6356 3024 6442 3080
rect 6498 3024 6570 3080
rect 6230 2938 6570 3024
rect 6230 2882 6300 2938
rect 6356 2882 6442 2938
rect 6498 2882 6570 2938
rect 6230 2796 6570 2882
rect 6230 2740 6300 2796
rect 6356 2740 6442 2796
rect 6498 2740 6570 2796
rect 6230 2654 6570 2740
rect 6230 2598 6300 2654
rect 6356 2598 6442 2654
rect 6498 2598 6570 2654
rect 6230 2512 6570 2598
rect 6230 2456 6300 2512
rect 6356 2456 6442 2512
rect 6498 2456 6570 2512
rect 6230 2370 6570 2456
rect 6230 2314 6300 2370
rect 6356 2314 6442 2370
rect 6498 2314 6570 2370
rect 6230 2228 6570 2314
rect 6230 2172 6300 2228
rect 6356 2172 6442 2228
rect 6498 2172 6570 2228
rect 6230 2086 6570 2172
rect 6230 2030 6300 2086
rect 6356 2030 6442 2086
rect 6498 2030 6570 2086
rect 6230 1944 6570 2030
rect 6230 1888 6300 1944
rect 6356 1888 6442 1944
rect 6498 1888 6570 1944
rect 6230 1802 6570 1888
rect 6230 1746 6300 1802
rect 6356 1746 6442 1802
rect 6498 1746 6570 1802
rect 6230 1660 6570 1746
rect 6230 1604 6300 1660
rect 6356 1604 6442 1660
rect 6498 1604 6570 1660
rect 6230 1518 6570 1604
rect 6230 1462 6300 1518
rect 6356 1462 6442 1518
rect 6498 1462 6570 1518
rect 6230 1376 6570 1462
rect 6230 1320 6300 1376
rect 6356 1320 6442 1376
rect 6498 1320 6570 1376
rect 6230 1234 6570 1320
rect 6230 1178 6300 1234
rect 6356 1178 6442 1234
rect 6498 1178 6570 1234
rect 6230 1092 6570 1178
rect 6230 1036 6300 1092
rect 6356 1036 6442 1092
rect 6498 1036 6570 1092
rect 6230 950 6570 1036
rect 6230 894 6300 950
rect 6356 894 6442 950
rect 6498 894 6570 950
rect 6230 808 6570 894
rect 6230 752 6300 808
rect 6356 752 6442 808
rect 6498 752 6570 808
rect 6230 666 6570 752
rect 6230 610 6300 666
rect 6356 610 6442 666
rect 6498 610 6570 666
rect 6230 524 6570 610
rect 6230 468 6300 524
rect 6356 468 6442 524
rect 6498 468 6570 524
rect 6230 458 6570 468
rect 6770 12310 7110 12320
rect 6770 12254 6845 12310
rect 6901 12254 6987 12310
rect 7043 12254 7110 12310
rect 6770 12168 7110 12254
rect 6770 12112 6845 12168
rect 6901 12112 6987 12168
rect 7043 12112 7110 12168
rect 6770 12026 7110 12112
rect 6770 11970 6845 12026
rect 6901 11970 6987 12026
rect 7043 11970 7110 12026
rect 6770 11884 7110 11970
rect 6770 11828 6845 11884
rect 6901 11828 6987 11884
rect 7043 11828 7110 11884
rect 6770 11742 7110 11828
rect 6770 11686 6845 11742
rect 6901 11686 6987 11742
rect 7043 11686 7110 11742
rect 6770 11600 7110 11686
rect 6770 11544 6845 11600
rect 6901 11544 6987 11600
rect 7043 11544 7110 11600
rect 6770 11458 7110 11544
rect 6770 11402 6845 11458
rect 6901 11402 6987 11458
rect 7043 11402 7110 11458
rect 6770 11316 7110 11402
rect 6770 11260 6845 11316
rect 6901 11260 6987 11316
rect 7043 11260 7110 11316
rect 6770 11174 7110 11260
rect 6770 11118 6845 11174
rect 6901 11118 6987 11174
rect 7043 11118 7110 11174
rect 6770 11032 7110 11118
rect 6770 10976 6845 11032
rect 6901 10976 6987 11032
rect 7043 10976 7110 11032
rect 6770 10890 7110 10976
rect 6770 10834 6845 10890
rect 6901 10834 6987 10890
rect 7043 10834 7110 10890
rect 6770 10748 7110 10834
rect 6770 10692 6845 10748
rect 6901 10692 6987 10748
rect 7043 10692 7110 10748
rect 6770 10606 7110 10692
rect 6770 10550 6845 10606
rect 6901 10550 6987 10606
rect 7043 10550 7110 10606
rect 6770 10464 7110 10550
rect 6770 10408 6845 10464
rect 6901 10408 6987 10464
rect 7043 10408 7110 10464
rect 6770 10322 7110 10408
rect 6770 10266 6845 10322
rect 6901 10266 6987 10322
rect 7043 10266 7110 10322
rect 6770 10180 7110 10266
rect 6770 10124 6845 10180
rect 6901 10124 6987 10180
rect 7043 10124 7110 10180
rect 6770 10038 7110 10124
rect 6770 9982 6845 10038
rect 6901 9982 6987 10038
rect 7043 9982 7110 10038
rect 6770 9896 7110 9982
rect 6770 9840 6845 9896
rect 6901 9840 6987 9896
rect 7043 9840 7110 9896
rect 6770 9754 7110 9840
rect 6770 9698 6845 9754
rect 6901 9698 6987 9754
rect 7043 9698 7110 9754
rect 6770 9612 7110 9698
rect 6770 9556 6845 9612
rect 6901 9556 6987 9612
rect 7043 9556 7110 9612
rect 6770 9470 7110 9556
rect 6770 9414 6845 9470
rect 6901 9414 6987 9470
rect 7043 9414 7110 9470
rect 6770 9328 7110 9414
rect 6770 9272 6845 9328
rect 6901 9272 6987 9328
rect 7043 9272 7110 9328
rect 6770 9186 7110 9272
rect 6770 9130 6845 9186
rect 6901 9130 6987 9186
rect 7043 9130 7110 9186
rect 6770 9044 7110 9130
rect 6770 8988 6845 9044
rect 6901 8988 6987 9044
rect 7043 8988 7110 9044
rect 6770 8902 7110 8988
rect 6770 8846 6845 8902
rect 6901 8846 6987 8902
rect 7043 8846 7110 8902
rect 6770 8760 7110 8846
rect 6770 8704 6845 8760
rect 6901 8704 6987 8760
rect 7043 8704 7110 8760
rect 6770 8618 7110 8704
rect 6770 8562 6845 8618
rect 6901 8562 6987 8618
rect 7043 8562 7110 8618
rect 6770 8476 7110 8562
rect 6770 8420 6845 8476
rect 6901 8420 6987 8476
rect 7043 8420 7110 8476
rect 6770 8334 7110 8420
rect 6770 8278 6845 8334
rect 6901 8278 6987 8334
rect 7043 8278 7110 8334
rect 6770 8192 7110 8278
rect 6770 8136 6845 8192
rect 6901 8136 6987 8192
rect 7043 8136 7110 8192
rect 6770 8050 7110 8136
rect 6770 7994 6845 8050
rect 6901 7994 6987 8050
rect 7043 7994 7110 8050
rect 6770 7908 7110 7994
rect 6770 7852 6845 7908
rect 6901 7852 6987 7908
rect 7043 7852 7110 7908
rect 6770 7766 7110 7852
rect 6770 7710 6845 7766
rect 6901 7710 6987 7766
rect 7043 7710 7110 7766
rect 6770 7624 7110 7710
rect 6770 7568 6845 7624
rect 6901 7568 6987 7624
rect 7043 7568 7110 7624
rect 6770 7482 7110 7568
rect 6770 7426 6845 7482
rect 6901 7426 6987 7482
rect 7043 7426 7110 7482
rect 6770 7340 7110 7426
rect 6770 7284 6845 7340
rect 6901 7284 6987 7340
rect 7043 7284 7110 7340
rect 6770 7198 7110 7284
rect 6770 7142 6845 7198
rect 6901 7142 6987 7198
rect 7043 7142 7110 7198
rect 6770 7056 7110 7142
rect 6770 7000 6845 7056
rect 6901 7000 6987 7056
rect 7043 7000 7110 7056
rect 6770 6914 7110 7000
rect 6770 6858 6845 6914
rect 6901 6858 6987 6914
rect 7043 6858 7110 6914
rect 6770 6772 7110 6858
rect 6770 6716 6845 6772
rect 6901 6716 6987 6772
rect 7043 6716 7110 6772
rect 6770 6630 7110 6716
rect 6770 6574 6845 6630
rect 6901 6574 6987 6630
rect 7043 6574 7110 6630
rect 6770 6488 7110 6574
rect 6770 6432 6845 6488
rect 6901 6432 6987 6488
rect 7043 6432 7110 6488
rect 6770 6346 7110 6432
rect 6770 6290 6845 6346
rect 6901 6290 6987 6346
rect 7043 6290 7110 6346
rect 6770 6204 7110 6290
rect 6770 6148 6845 6204
rect 6901 6148 6987 6204
rect 7043 6148 7110 6204
rect 6770 6062 7110 6148
rect 6770 6006 6845 6062
rect 6901 6006 6987 6062
rect 7043 6006 7110 6062
rect 6770 5920 7110 6006
rect 6770 5864 6845 5920
rect 6901 5864 6987 5920
rect 7043 5864 7110 5920
rect 6770 5778 7110 5864
rect 6770 5722 6845 5778
rect 6901 5722 6987 5778
rect 7043 5722 7110 5778
rect 6770 5636 7110 5722
rect 6770 5580 6845 5636
rect 6901 5580 6987 5636
rect 7043 5580 7110 5636
rect 6770 5494 7110 5580
rect 6770 5438 6845 5494
rect 6901 5438 6987 5494
rect 7043 5438 7110 5494
rect 6770 5352 7110 5438
rect 6770 5296 6845 5352
rect 6901 5296 6987 5352
rect 7043 5296 7110 5352
rect 6770 5210 7110 5296
rect 6770 5154 6845 5210
rect 6901 5154 6987 5210
rect 7043 5154 7110 5210
rect 6770 5068 7110 5154
rect 6770 5012 6845 5068
rect 6901 5012 6987 5068
rect 7043 5012 7110 5068
rect 6770 4926 7110 5012
rect 6770 4870 6845 4926
rect 6901 4870 6987 4926
rect 7043 4870 7110 4926
rect 6770 4784 7110 4870
rect 6770 4728 6845 4784
rect 6901 4728 6987 4784
rect 7043 4728 7110 4784
rect 6770 4642 7110 4728
rect 6770 4586 6845 4642
rect 6901 4586 6987 4642
rect 7043 4586 7110 4642
rect 6770 4500 7110 4586
rect 6770 4444 6845 4500
rect 6901 4444 6987 4500
rect 7043 4444 7110 4500
rect 6770 4358 7110 4444
rect 6770 4302 6845 4358
rect 6901 4302 6987 4358
rect 7043 4302 7110 4358
rect 6770 4216 7110 4302
rect 6770 4160 6845 4216
rect 6901 4160 6987 4216
rect 7043 4160 7110 4216
rect 6770 4074 7110 4160
rect 6770 4018 6845 4074
rect 6901 4018 6987 4074
rect 7043 4018 7110 4074
rect 6770 3932 7110 4018
rect 6770 3876 6845 3932
rect 6901 3876 6987 3932
rect 7043 3876 7110 3932
rect 6770 3790 7110 3876
rect 6770 3734 6845 3790
rect 6901 3734 6987 3790
rect 7043 3734 7110 3790
rect 6770 3648 7110 3734
rect 6770 3592 6845 3648
rect 6901 3592 6987 3648
rect 7043 3592 7110 3648
rect 6770 3506 7110 3592
rect 6770 3450 6845 3506
rect 6901 3450 6987 3506
rect 7043 3450 7110 3506
rect 6770 3364 7110 3450
rect 6770 3308 6845 3364
rect 6901 3308 6987 3364
rect 7043 3308 7110 3364
rect 6770 3222 7110 3308
rect 6770 3166 6845 3222
rect 6901 3166 6987 3222
rect 7043 3166 7110 3222
rect 6770 3080 7110 3166
rect 6770 3024 6845 3080
rect 6901 3024 6987 3080
rect 7043 3024 7110 3080
rect 6770 2938 7110 3024
rect 6770 2882 6845 2938
rect 6901 2882 6987 2938
rect 7043 2882 7110 2938
rect 6770 2796 7110 2882
rect 6770 2740 6845 2796
rect 6901 2740 6987 2796
rect 7043 2740 7110 2796
rect 6770 2654 7110 2740
rect 6770 2598 6845 2654
rect 6901 2598 6987 2654
rect 7043 2598 7110 2654
rect 6770 2512 7110 2598
rect 6770 2456 6845 2512
rect 6901 2456 6987 2512
rect 7043 2456 7110 2512
rect 6770 2370 7110 2456
rect 6770 2314 6845 2370
rect 6901 2314 6987 2370
rect 7043 2314 7110 2370
rect 6770 2228 7110 2314
rect 6770 2172 6845 2228
rect 6901 2172 6987 2228
rect 7043 2172 7110 2228
rect 6770 2086 7110 2172
rect 6770 2030 6845 2086
rect 6901 2030 6987 2086
rect 7043 2030 7110 2086
rect 6770 1944 7110 2030
rect 6770 1888 6845 1944
rect 6901 1888 6987 1944
rect 7043 1888 7110 1944
rect 6770 1802 7110 1888
rect 6770 1746 6845 1802
rect 6901 1746 6987 1802
rect 7043 1746 7110 1802
rect 6770 1660 7110 1746
rect 6770 1604 6845 1660
rect 6901 1604 6987 1660
rect 7043 1604 7110 1660
rect 6770 1518 7110 1604
rect 6770 1462 6845 1518
rect 6901 1462 6987 1518
rect 7043 1462 7110 1518
rect 6770 1376 7110 1462
rect 6770 1320 6845 1376
rect 6901 1320 6987 1376
rect 7043 1320 7110 1376
rect 6770 1234 7110 1320
rect 6770 1178 6845 1234
rect 6901 1178 6987 1234
rect 7043 1178 7110 1234
rect 6770 1092 7110 1178
rect 6770 1036 6845 1092
rect 6901 1036 6987 1092
rect 7043 1036 7110 1092
rect 6770 950 7110 1036
rect 6770 894 6845 950
rect 6901 894 6987 950
rect 7043 894 7110 950
rect 6770 808 7110 894
rect 6770 752 6845 808
rect 6901 752 6987 808
rect 7043 752 7110 808
rect 6770 666 7110 752
rect 6770 610 6845 666
rect 6901 610 6987 666
rect 7043 610 7110 666
rect 6770 524 7110 610
rect 6770 468 6845 524
rect 6901 468 6987 524
rect 7043 468 7110 524
rect 6770 458 7110 468
rect 7310 12310 7650 12320
rect 7310 12254 7382 12310
rect 7438 12254 7524 12310
rect 7580 12254 7650 12310
rect 7310 12168 7650 12254
rect 7310 12112 7382 12168
rect 7438 12112 7524 12168
rect 7580 12112 7650 12168
rect 7310 12026 7650 12112
rect 7310 11970 7382 12026
rect 7438 11970 7524 12026
rect 7580 11970 7650 12026
rect 7310 11884 7650 11970
rect 7310 11828 7382 11884
rect 7438 11828 7524 11884
rect 7580 11828 7650 11884
rect 7310 11742 7650 11828
rect 7310 11686 7382 11742
rect 7438 11686 7524 11742
rect 7580 11686 7650 11742
rect 7310 11600 7650 11686
rect 7310 11544 7382 11600
rect 7438 11544 7524 11600
rect 7580 11544 7650 11600
rect 7310 11458 7650 11544
rect 7310 11402 7382 11458
rect 7438 11402 7524 11458
rect 7580 11402 7650 11458
rect 7310 11316 7650 11402
rect 7310 11260 7382 11316
rect 7438 11260 7524 11316
rect 7580 11260 7650 11316
rect 7310 11174 7650 11260
rect 7310 11118 7382 11174
rect 7438 11118 7524 11174
rect 7580 11118 7650 11174
rect 7310 11032 7650 11118
rect 7310 10976 7382 11032
rect 7438 10976 7524 11032
rect 7580 10976 7650 11032
rect 7310 10890 7650 10976
rect 7310 10834 7382 10890
rect 7438 10834 7524 10890
rect 7580 10834 7650 10890
rect 7310 10748 7650 10834
rect 7310 10692 7382 10748
rect 7438 10692 7524 10748
rect 7580 10692 7650 10748
rect 7310 10606 7650 10692
rect 7310 10550 7382 10606
rect 7438 10550 7524 10606
rect 7580 10550 7650 10606
rect 7310 10464 7650 10550
rect 7310 10408 7382 10464
rect 7438 10408 7524 10464
rect 7580 10408 7650 10464
rect 7310 10322 7650 10408
rect 7310 10266 7382 10322
rect 7438 10266 7524 10322
rect 7580 10266 7650 10322
rect 7310 10180 7650 10266
rect 7310 10124 7382 10180
rect 7438 10124 7524 10180
rect 7580 10124 7650 10180
rect 7310 10038 7650 10124
rect 7310 9982 7382 10038
rect 7438 9982 7524 10038
rect 7580 9982 7650 10038
rect 7310 9896 7650 9982
rect 7310 9840 7382 9896
rect 7438 9840 7524 9896
rect 7580 9840 7650 9896
rect 7310 9754 7650 9840
rect 7310 9698 7382 9754
rect 7438 9698 7524 9754
rect 7580 9698 7650 9754
rect 7310 9612 7650 9698
rect 7310 9556 7382 9612
rect 7438 9556 7524 9612
rect 7580 9556 7650 9612
rect 7310 9470 7650 9556
rect 7310 9414 7382 9470
rect 7438 9414 7524 9470
rect 7580 9414 7650 9470
rect 7310 9328 7650 9414
rect 7310 9272 7382 9328
rect 7438 9272 7524 9328
rect 7580 9272 7650 9328
rect 7310 9186 7650 9272
rect 7310 9130 7382 9186
rect 7438 9130 7524 9186
rect 7580 9130 7650 9186
rect 7310 9044 7650 9130
rect 7310 8988 7382 9044
rect 7438 8988 7524 9044
rect 7580 8988 7650 9044
rect 7310 8902 7650 8988
rect 7310 8846 7382 8902
rect 7438 8846 7524 8902
rect 7580 8846 7650 8902
rect 7310 8760 7650 8846
rect 7310 8704 7382 8760
rect 7438 8704 7524 8760
rect 7580 8704 7650 8760
rect 7310 8618 7650 8704
rect 7310 8562 7382 8618
rect 7438 8562 7524 8618
rect 7580 8562 7650 8618
rect 7310 8476 7650 8562
rect 7310 8420 7382 8476
rect 7438 8420 7524 8476
rect 7580 8420 7650 8476
rect 7310 8334 7650 8420
rect 7310 8278 7382 8334
rect 7438 8278 7524 8334
rect 7580 8278 7650 8334
rect 7310 8192 7650 8278
rect 7310 8136 7382 8192
rect 7438 8136 7524 8192
rect 7580 8136 7650 8192
rect 7310 8050 7650 8136
rect 7310 7994 7382 8050
rect 7438 7994 7524 8050
rect 7580 7994 7650 8050
rect 7310 7908 7650 7994
rect 7310 7852 7382 7908
rect 7438 7852 7524 7908
rect 7580 7852 7650 7908
rect 7310 7766 7650 7852
rect 7310 7710 7382 7766
rect 7438 7710 7524 7766
rect 7580 7710 7650 7766
rect 7310 7624 7650 7710
rect 7310 7568 7382 7624
rect 7438 7568 7524 7624
rect 7580 7568 7650 7624
rect 7310 7482 7650 7568
rect 7310 7426 7382 7482
rect 7438 7426 7524 7482
rect 7580 7426 7650 7482
rect 7310 7340 7650 7426
rect 7310 7284 7382 7340
rect 7438 7284 7524 7340
rect 7580 7284 7650 7340
rect 7310 7198 7650 7284
rect 7310 7142 7382 7198
rect 7438 7142 7524 7198
rect 7580 7142 7650 7198
rect 7310 7056 7650 7142
rect 7310 7000 7382 7056
rect 7438 7000 7524 7056
rect 7580 7000 7650 7056
rect 7310 6914 7650 7000
rect 7310 6858 7382 6914
rect 7438 6858 7524 6914
rect 7580 6858 7650 6914
rect 7310 6772 7650 6858
rect 7310 6716 7382 6772
rect 7438 6716 7524 6772
rect 7580 6716 7650 6772
rect 7310 6630 7650 6716
rect 7310 6574 7382 6630
rect 7438 6574 7524 6630
rect 7580 6574 7650 6630
rect 7310 6488 7650 6574
rect 7310 6432 7382 6488
rect 7438 6432 7524 6488
rect 7580 6432 7650 6488
rect 7310 6346 7650 6432
rect 7310 6290 7382 6346
rect 7438 6290 7524 6346
rect 7580 6290 7650 6346
rect 7310 6204 7650 6290
rect 7310 6148 7382 6204
rect 7438 6148 7524 6204
rect 7580 6148 7650 6204
rect 7310 6062 7650 6148
rect 7310 6006 7382 6062
rect 7438 6006 7524 6062
rect 7580 6006 7650 6062
rect 7310 5920 7650 6006
rect 7310 5864 7382 5920
rect 7438 5864 7524 5920
rect 7580 5864 7650 5920
rect 7310 5778 7650 5864
rect 7310 5722 7382 5778
rect 7438 5722 7524 5778
rect 7580 5722 7650 5778
rect 7310 5636 7650 5722
rect 7310 5580 7382 5636
rect 7438 5580 7524 5636
rect 7580 5580 7650 5636
rect 7310 5494 7650 5580
rect 7310 5438 7382 5494
rect 7438 5438 7524 5494
rect 7580 5438 7650 5494
rect 7310 5352 7650 5438
rect 7310 5296 7382 5352
rect 7438 5296 7524 5352
rect 7580 5296 7650 5352
rect 7310 5210 7650 5296
rect 7310 5154 7382 5210
rect 7438 5154 7524 5210
rect 7580 5154 7650 5210
rect 7310 5068 7650 5154
rect 7310 5012 7382 5068
rect 7438 5012 7524 5068
rect 7580 5012 7650 5068
rect 7310 4926 7650 5012
rect 7310 4870 7382 4926
rect 7438 4870 7524 4926
rect 7580 4870 7650 4926
rect 7310 4784 7650 4870
rect 7310 4728 7382 4784
rect 7438 4728 7524 4784
rect 7580 4728 7650 4784
rect 7310 4642 7650 4728
rect 7310 4586 7382 4642
rect 7438 4586 7524 4642
rect 7580 4586 7650 4642
rect 7310 4500 7650 4586
rect 7310 4444 7382 4500
rect 7438 4444 7524 4500
rect 7580 4444 7650 4500
rect 7310 4358 7650 4444
rect 7310 4302 7382 4358
rect 7438 4302 7524 4358
rect 7580 4302 7650 4358
rect 7310 4216 7650 4302
rect 7310 4160 7382 4216
rect 7438 4160 7524 4216
rect 7580 4160 7650 4216
rect 7310 4074 7650 4160
rect 7310 4018 7382 4074
rect 7438 4018 7524 4074
rect 7580 4018 7650 4074
rect 7310 3932 7650 4018
rect 7310 3876 7382 3932
rect 7438 3876 7524 3932
rect 7580 3876 7650 3932
rect 7310 3790 7650 3876
rect 7310 3734 7382 3790
rect 7438 3734 7524 3790
rect 7580 3734 7650 3790
rect 7310 3648 7650 3734
rect 7310 3592 7382 3648
rect 7438 3592 7524 3648
rect 7580 3592 7650 3648
rect 7310 3506 7650 3592
rect 7310 3450 7382 3506
rect 7438 3450 7524 3506
rect 7580 3450 7650 3506
rect 7310 3364 7650 3450
rect 7310 3308 7382 3364
rect 7438 3308 7524 3364
rect 7580 3308 7650 3364
rect 7310 3222 7650 3308
rect 7310 3166 7382 3222
rect 7438 3166 7524 3222
rect 7580 3166 7650 3222
rect 7310 3080 7650 3166
rect 7310 3024 7382 3080
rect 7438 3024 7524 3080
rect 7580 3024 7650 3080
rect 7310 2938 7650 3024
rect 7310 2882 7382 2938
rect 7438 2882 7524 2938
rect 7580 2882 7650 2938
rect 7310 2796 7650 2882
rect 7310 2740 7382 2796
rect 7438 2740 7524 2796
rect 7580 2740 7650 2796
rect 7310 2654 7650 2740
rect 7310 2598 7382 2654
rect 7438 2598 7524 2654
rect 7580 2598 7650 2654
rect 7310 2512 7650 2598
rect 7310 2456 7382 2512
rect 7438 2456 7524 2512
rect 7580 2456 7650 2512
rect 7310 2370 7650 2456
rect 7310 2314 7382 2370
rect 7438 2314 7524 2370
rect 7580 2314 7650 2370
rect 7310 2228 7650 2314
rect 7310 2172 7382 2228
rect 7438 2172 7524 2228
rect 7580 2172 7650 2228
rect 7310 2086 7650 2172
rect 7310 2030 7382 2086
rect 7438 2030 7524 2086
rect 7580 2030 7650 2086
rect 7310 1944 7650 2030
rect 7310 1888 7382 1944
rect 7438 1888 7524 1944
rect 7580 1888 7650 1944
rect 7310 1802 7650 1888
rect 7310 1746 7382 1802
rect 7438 1746 7524 1802
rect 7580 1746 7650 1802
rect 7310 1660 7650 1746
rect 7310 1604 7382 1660
rect 7438 1604 7524 1660
rect 7580 1604 7650 1660
rect 7310 1518 7650 1604
rect 7310 1462 7382 1518
rect 7438 1462 7524 1518
rect 7580 1462 7650 1518
rect 7310 1376 7650 1462
rect 7310 1320 7382 1376
rect 7438 1320 7524 1376
rect 7580 1320 7650 1376
rect 7310 1234 7650 1320
rect 7310 1178 7382 1234
rect 7438 1178 7524 1234
rect 7580 1178 7650 1234
rect 7310 1092 7650 1178
rect 7310 1036 7382 1092
rect 7438 1036 7524 1092
rect 7580 1036 7650 1092
rect 7310 950 7650 1036
rect 7310 894 7382 950
rect 7438 894 7524 950
rect 7580 894 7650 950
rect 7310 808 7650 894
rect 7310 752 7382 808
rect 7438 752 7524 808
rect 7580 752 7650 808
rect 7310 666 7650 752
rect 7310 610 7382 666
rect 7438 610 7524 666
rect 7580 610 7650 666
rect 7310 524 7650 610
rect 7310 468 7382 524
rect 7438 468 7524 524
rect 7580 468 7650 524
rect 7310 458 7650 468
rect 7850 12310 8190 12320
rect 7850 12254 7919 12310
rect 7975 12254 8061 12310
rect 8117 12254 8190 12310
rect 7850 12168 8190 12254
rect 7850 12112 7919 12168
rect 7975 12112 8061 12168
rect 8117 12112 8190 12168
rect 7850 12026 8190 12112
rect 7850 11970 7919 12026
rect 7975 11970 8061 12026
rect 8117 11970 8190 12026
rect 7850 11884 8190 11970
rect 7850 11828 7919 11884
rect 7975 11828 8061 11884
rect 8117 11828 8190 11884
rect 7850 11742 8190 11828
rect 7850 11686 7919 11742
rect 7975 11686 8061 11742
rect 8117 11686 8190 11742
rect 7850 11600 8190 11686
rect 7850 11544 7919 11600
rect 7975 11544 8061 11600
rect 8117 11544 8190 11600
rect 7850 11458 8190 11544
rect 7850 11402 7919 11458
rect 7975 11402 8061 11458
rect 8117 11402 8190 11458
rect 7850 11316 8190 11402
rect 7850 11260 7919 11316
rect 7975 11260 8061 11316
rect 8117 11260 8190 11316
rect 7850 11174 8190 11260
rect 7850 11118 7919 11174
rect 7975 11118 8061 11174
rect 8117 11118 8190 11174
rect 7850 11032 8190 11118
rect 7850 10976 7919 11032
rect 7975 10976 8061 11032
rect 8117 10976 8190 11032
rect 7850 10890 8190 10976
rect 7850 10834 7919 10890
rect 7975 10834 8061 10890
rect 8117 10834 8190 10890
rect 7850 10748 8190 10834
rect 7850 10692 7919 10748
rect 7975 10692 8061 10748
rect 8117 10692 8190 10748
rect 7850 10606 8190 10692
rect 7850 10550 7919 10606
rect 7975 10550 8061 10606
rect 8117 10550 8190 10606
rect 7850 10464 8190 10550
rect 7850 10408 7919 10464
rect 7975 10408 8061 10464
rect 8117 10408 8190 10464
rect 7850 10322 8190 10408
rect 7850 10266 7919 10322
rect 7975 10266 8061 10322
rect 8117 10266 8190 10322
rect 7850 10180 8190 10266
rect 7850 10124 7919 10180
rect 7975 10124 8061 10180
rect 8117 10124 8190 10180
rect 7850 10038 8190 10124
rect 7850 9982 7919 10038
rect 7975 9982 8061 10038
rect 8117 9982 8190 10038
rect 7850 9896 8190 9982
rect 7850 9840 7919 9896
rect 7975 9840 8061 9896
rect 8117 9840 8190 9896
rect 7850 9754 8190 9840
rect 7850 9698 7919 9754
rect 7975 9698 8061 9754
rect 8117 9698 8190 9754
rect 7850 9612 8190 9698
rect 7850 9556 7919 9612
rect 7975 9556 8061 9612
rect 8117 9556 8190 9612
rect 7850 9470 8190 9556
rect 7850 9414 7919 9470
rect 7975 9414 8061 9470
rect 8117 9414 8190 9470
rect 7850 9328 8190 9414
rect 7850 9272 7919 9328
rect 7975 9272 8061 9328
rect 8117 9272 8190 9328
rect 7850 9186 8190 9272
rect 7850 9130 7919 9186
rect 7975 9130 8061 9186
rect 8117 9130 8190 9186
rect 7850 9044 8190 9130
rect 7850 8988 7919 9044
rect 7975 8988 8061 9044
rect 8117 8988 8190 9044
rect 7850 8902 8190 8988
rect 7850 8846 7919 8902
rect 7975 8846 8061 8902
rect 8117 8846 8190 8902
rect 7850 8760 8190 8846
rect 7850 8704 7919 8760
rect 7975 8704 8061 8760
rect 8117 8704 8190 8760
rect 7850 8618 8190 8704
rect 7850 8562 7919 8618
rect 7975 8562 8061 8618
rect 8117 8562 8190 8618
rect 7850 8476 8190 8562
rect 7850 8420 7919 8476
rect 7975 8420 8061 8476
rect 8117 8420 8190 8476
rect 7850 8334 8190 8420
rect 7850 8278 7919 8334
rect 7975 8278 8061 8334
rect 8117 8278 8190 8334
rect 7850 8192 8190 8278
rect 7850 8136 7919 8192
rect 7975 8136 8061 8192
rect 8117 8136 8190 8192
rect 7850 8050 8190 8136
rect 7850 7994 7919 8050
rect 7975 7994 8061 8050
rect 8117 7994 8190 8050
rect 7850 7908 8190 7994
rect 7850 7852 7919 7908
rect 7975 7852 8061 7908
rect 8117 7852 8190 7908
rect 7850 7766 8190 7852
rect 7850 7710 7919 7766
rect 7975 7710 8061 7766
rect 8117 7710 8190 7766
rect 7850 7624 8190 7710
rect 7850 7568 7919 7624
rect 7975 7568 8061 7624
rect 8117 7568 8190 7624
rect 7850 7482 8190 7568
rect 7850 7426 7919 7482
rect 7975 7426 8061 7482
rect 8117 7426 8190 7482
rect 7850 7340 8190 7426
rect 7850 7284 7919 7340
rect 7975 7284 8061 7340
rect 8117 7284 8190 7340
rect 7850 7198 8190 7284
rect 7850 7142 7919 7198
rect 7975 7142 8061 7198
rect 8117 7142 8190 7198
rect 7850 7056 8190 7142
rect 7850 7000 7919 7056
rect 7975 7000 8061 7056
rect 8117 7000 8190 7056
rect 7850 6914 8190 7000
rect 7850 6858 7919 6914
rect 7975 6858 8061 6914
rect 8117 6858 8190 6914
rect 7850 6772 8190 6858
rect 7850 6716 7919 6772
rect 7975 6716 8061 6772
rect 8117 6716 8190 6772
rect 7850 6630 8190 6716
rect 7850 6574 7919 6630
rect 7975 6574 8061 6630
rect 8117 6574 8190 6630
rect 7850 6488 8190 6574
rect 7850 6432 7919 6488
rect 7975 6432 8061 6488
rect 8117 6432 8190 6488
rect 7850 6346 8190 6432
rect 7850 6290 7919 6346
rect 7975 6290 8061 6346
rect 8117 6290 8190 6346
rect 7850 6204 8190 6290
rect 7850 6148 7919 6204
rect 7975 6148 8061 6204
rect 8117 6148 8190 6204
rect 7850 6062 8190 6148
rect 7850 6006 7919 6062
rect 7975 6006 8061 6062
rect 8117 6006 8190 6062
rect 7850 5920 8190 6006
rect 7850 5864 7919 5920
rect 7975 5864 8061 5920
rect 8117 5864 8190 5920
rect 7850 5778 8190 5864
rect 7850 5722 7919 5778
rect 7975 5722 8061 5778
rect 8117 5722 8190 5778
rect 7850 5636 8190 5722
rect 7850 5580 7919 5636
rect 7975 5580 8061 5636
rect 8117 5580 8190 5636
rect 7850 5494 8190 5580
rect 7850 5438 7919 5494
rect 7975 5438 8061 5494
rect 8117 5438 8190 5494
rect 7850 5352 8190 5438
rect 7850 5296 7919 5352
rect 7975 5296 8061 5352
rect 8117 5296 8190 5352
rect 7850 5210 8190 5296
rect 7850 5154 7919 5210
rect 7975 5154 8061 5210
rect 8117 5154 8190 5210
rect 7850 5068 8190 5154
rect 7850 5012 7919 5068
rect 7975 5012 8061 5068
rect 8117 5012 8190 5068
rect 7850 4926 8190 5012
rect 7850 4870 7919 4926
rect 7975 4870 8061 4926
rect 8117 4870 8190 4926
rect 7850 4784 8190 4870
rect 7850 4728 7919 4784
rect 7975 4728 8061 4784
rect 8117 4728 8190 4784
rect 7850 4642 8190 4728
rect 7850 4586 7919 4642
rect 7975 4586 8061 4642
rect 8117 4586 8190 4642
rect 7850 4500 8190 4586
rect 7850 4444 7919 4500
rect 7975 4444 8061 4500
rect 8117 4444 8190 4500
rect 7850 4358 8190 4444
rect 7850 4302 7919 4358
rect 7975 4302 8061 4358
rect 8117 4302 8190 4358
rect 7850 4216 8190 4302
rect 7850 4160 7919 4216
rect 7975 4160 8061 4216
rect 8117 4160 8190 4216
rect 7850 4074 8190 4160
rect 7850 4018 7919 4074
rect 7975 4018 8061 4074
rect 8117 4018 8190 4074
rect 7850 3932 8190 4018
rect 7850 3876 7919 3932
rect 7975 3876 8061 3932
rect 8117 3876 8190 3932
rect 7850 3790 8190 3876
rect 7850 3734 7919 3790
rect 7975 3734 8061 3790
rect 8117 3734 8190 3790
rect 7850 3648 8190 3734
rect 7850 3592 7919 3648
rect 7975 3592 8061 3648
rect 8117 3592 8190 3648
rect 7850 3506 8190 3592
rect 7850 3450 7919 3506
rect 7975 3450 8061 3506
rect 8117 3450 8190 3506
rect 7850 3364 8190 3450
rect 7850 3308 7919 3364
rect 7975 3308 8061 3364
rect 8117 3308 8190 3364
rect 7850 3222 8190 3308
rect 7850 3166 7919 3222
rect 7975 3166 8061 3222
rect 8117 3166 8190 3222
rect 7850 3080 8190 3166
rect 7850 3024 7919 3080
rect 7975 3024 8061 3080
rect 8117 3024 8190 3080
rect 7850 2938 8190 3024
rect 7850 2882 7919 2938
rect 7975 2882 8061 2938
rect 8117 2882 8190 2938
rect 7850 2796 8190 2882
rect 7850 2740 7919 2796
rect 7975 2740 8061 2796
rect 8117 2740 8190 2796
rect 7850 2654 8190 2740
rect 7850 2598 7919 2654
rect 7975 2598 8061 2654
rect 8117 2598 8190 2654
rect 7850 2512 8190 2598
rect 7850 2456 7919 2512
rect 7975 2456 8061 2512
rect 8117 2456 8190 2512
rect 7850 2370 8190 2456
rect 7850 2314 7919 2370
rect 7975 2314 8061 2370
rect 8117 2314 8190 2370
rect 7850 2228 8190 2314
rect 7850 2172 7919 2228
rect 7975 2172 8061 2228
rect 8117 2172 8190 2228
rect 7850 2086 8190 2172
rect 7850 2030 7919 2086
rect 7975 2030 8061 2086
rect 8117 2030 8190 2086
rect 7850 1944 8190 2030
rect 7850 1888 7919 1944
rect 7975 1888 8061 1944
rect 8117 1888 8190 1944
rect 7850 1802 8190 1888
rect 7850 1746 7919 1802
rect 7975 1746 8061 1802
rect 8117 1746 8190 1802
rect 7850 1660 8190 1746
rect 7850 1604 7919 1660
rect 7975 1604 8061 1660
rect 8117 1604 8190 1660
rect 7850 1518 8190 1604
rect 7850 1462 7919 1518
rect 7975 1462 8061 1518
rect 8117 1462 8190 1518
rect 7850 1376 8190 1462
rect 7850 1320 7919 1376
rect 7975 1320 8061 1376
rect 8117 1320 8190 1376
rect 7850 1234 8190 1320
rect 7850 1178 7919 1234
rect 7975 1178 8061 1234
rect 8117 1178 8190 1234
rect 7850 1092 8190 1178
rect 7850 1036 7919 1092
rect 7975 1036 8061 1092
rect 8117 1036 8190 1092
rect 7850 950 8190 1036
rect 7850 894 7919 950
rect 7975 894 8061 950
rect 8117 894 8190 950
rect 7850 808 8190 894
rect 7850 752 7919 808
rect 7975 752 8061 808
rect 8117 752 8190 808
rect 7850 666 8190 752
rect 7850 610 7919 666
rect 7975 610 8061 666
rect 8117 610 8190 666
rect 7850 524 8190 610
rect 7850 468 7919 524
rect 7975 468 8061 524
rect 8117 468 8190 524
rect 7850 458 8190 468
rect 8390 12310 8730 12320
rect 8390 12254 8462 12310
rect 8518 12254 8604 12310
rect 8660 12254 8730 12310
rect 8390 12168 8730 12254
rect 8390 12112 8462 12168
rect 8518 12112 8604 12168
rect 8660 12112 8730 12168
rect 8390 12026 8730 12112
rect 8390 11970 8462 12026
rect 8518 11970 8604 12026
rect 8660 11970 8730 12026
rect 8390 11884 8730 11970
rect 8390 11828 8462 11884
rect 8518 11828 8604 11884
rect 8660 11828 8730 11884
rect 8390 11742 8730 11828
rect 8390 11686 8462 11742
rect 8518 11686 8604 11742
rect 8660 11686 8730 11742
rect 8390 11600 8730 11686
rect 8390 11544 8462 11600
rect 8518 11544 8604 11600
rect 8660 11544 8730 11600
rect 8390 11458 8730 11544
rect 8390 11402 8462 11458
rect 8518 11402 8604 11458
rect 8660 11402 8730 11458
rect 8390 11316 8730 11402
rect 8390 11260 8462 11316
rect 8518 11260 8604 11316
rect 8660 11260 8730 11316
rect 8390 11174 8730 11260
rect 8390 11118 8462 11174
rect 8518 11118 8604 11174
rect 8660 11118 8730 11174
rect 8390 11032 8730 11118
rect 8390 10976 8462 11032
rect 8518 10976 8604 11032
rect 8660 10976 8730 11032
rect 8390 10890 8730 10976
rect 8390 10834 8462 10890
rect 8518 10834 8604 10890
rect 8660 10834 8730 10890
rect 8390 10748 8730 10834
rect 8390 10692 8462 10748
rect 8518 10692 8604 10748
rect 8660 10692 8730 10748
rect 8390 10606 8730 10692
rect 8390 10550 8462 10606
rect 8518 10550 8604 10606
rect 8660 10550 8730 10606
rect 8390 10464 8730 10550
rect 8390 10408 8462 10464
rect 8518 10408 8604 10464
rect 8660 10408 8730 10464
rect 8390 10322 8730 10408
rect 8390 10266 8462 10322
rect 8518 10266 8604 10322
rect 8660 10266 8730 10322
rect 8390 10180 8730 10266
rect 8390 10124 8462 10180
rect 8518 10124 8604 10180
rect 8660 10124 8730 10180
rect 8390 10038 8730 10124
rect 8390 9982 8462 10038
rect 8518 9982 8604 10038
rect 8660 9982 8730 10038
rect 8390 9896 8730 9982
rect 8390 9840 8462 9896
rect 8518 9840 8604 9896
rect 8660 9840 8730 9896
rect 8390 9754 8730 9840
rect 8390 9698 8462 9754
rect 8518 9698 8604 9754
rect 8660 9698 8730 9754
rect 8390 9612 8730 9698
rect 8390 9556 8462 9612
rect 8518 9556 8604 9612
rect 8660 9556 8730 9612
rect 8390 9470 8730 9556
rect 8390 9414 8462 9470
rect 8518 9414 8604 9470
rect 8660 9414 8730 9470
rect 8390 9328 8730 9414
rect 8390 9272 8462 9328
rect 8518 9272 8604 9328
rect 8660 9272 8730 9328
rect 8390 9186 8730 9272
rect 8390 9130 8462 9186
rect 8518 9130 8604 9186
rect 8660 9130 8730 9186
rect 8390 9044 8730 9130
rect 8390 8988 8462 9044
rect 8518 8988 8604 9044
rect 8660 8988 8730 9044
rect 8390 8902 8730 8988
rect 8390 8846 8462 8902
rect 8518 8846 8604 8902
rect 8660 8846 8730 8902
rect 8390 8760 8730 8846
rect 8390 8704 8462 8760
rect 8518 8704 8604 8760
rect 8660 8704 8730 8760
rect 8390 8618 8730 8704
rect 8390 8562 8462 8618
rect 8518 8562 8604 8618
rect 8660 8562 8730 8618
rect 8390 8476 8730 8562
rect 8390 8420 8462 8476
rect 8518 8420 8604 8476
rect 8660 8420 8730 8476
rect 8390 8334 8730 8420
rect 8390 8278 8462 8334
rect 8518 8278 8604 8334
rect 8660 8278 8730 8334
rect 8390 8192 8730 8278
rect 8390 8136 8462 8192
rect 8518 8136 8604 8192
rect 8660 8136 8730 8192
rect 8390 8050 8730 8136
rect 8390 7994 8462 8050
rect 8518 7994 8604 8050
rect 8660 7994 8730 8050
rect 8390 7908 8730 7994
rect 8390 7852 8462 7908
rect 8518 7852 8604 7908
rect 8660 7852 8730 7908
rect 8390 7766 8730 7852
rect 8390 7710 8462 7766
rect 8518 7710 8604 7766
rect 8660 7710 8730 7766
rect 8390 7624 8730 7710
rect 8390 7568 8462 7624
rect 8518 7568 8604 7624
rect 8660 7568 8730 7624
rect 8390 7482 8730 7568
rect 8390 7426 8462 7482
rect 8518 7426 8604 7482
rect 8660 7426 8730 7482
rect 8390 7340 8730 7426
rect 8390 7284 8462 7340
rect 8518 7284 8604 7340
rect 8660 7284 8730 7340
rect 8390 7198 8730 7284
rect 8390 7142 8462 7198
rect 8518 7142 8604 7198
rect 8660 7142 8730 7198
rect 8390 7056 8730 7142
rect 8390 7000 8462 7056
rect 8518 7000 8604 7056
rect 8660 7000 8730 7056
rect 8390 6914 8730 7000
rect 8390 6858 8462 6914
rect 8518 6858 8604 6914
rect 8660 6858 8730 6914
rect 8390 6772 8730 6858
rect 8390 6716 8462 6772
rect 8518 6716 8604 6772
rect 8660 6716 8730 6772
rect 8390 6630 8730 6716
rect 8390 6574 8462 6630
rect 8518 6574 8604 6630
rect 8660 6574 8730 6630
rect 8390 6488 8730 6574
rect 8390 6432 8462 6488
rect 8518 6432 8604 6488
rect 8660 6432 8730 6488
rect 8390 6346 8730 6432
rect 8390 6290 8462 6346
rect 8518 6290 8604 6346
rect 8660 6290 8730 6346
rect 8390 6204 8730 6290
rect 8390 6148 8462 6204
rect 8518 6148 8604 6204
rect 8660 6148 8730 6204
rect 8390 6062 8730 6148
rect 8390 6006 8462 6062
rect 8518 6006 8604 6062
rect 8660 6006 8730 6062
rect 8390 5920 8730 6006
rect 8390 5864 8462 5920
rect 8518 5864 8604 5920
rect 8660 5864 8730 5920
rect 8390 5778 8730 5864
rect 8390 5722 8462 5778
rect 8518 5722 8604 5778
rect 8660 5722 8730 5778
rect 8390 5636 8730 5722
rect 8390 5580 8462 5636
rect 8518 5580 8604 5636
rect 8660 5580 8730 5636
rect 8390 5494 8730 5580
rect 8390 5438 8462 5494
rect 8518 5438 8604 5494
rect 8660 5438 8730 5494
rect 8390 5352 8730 5438
rect 8390 5296 8462 5352
rect 8518 5296 8604 5352
rect 8660 5296 8730 5352
rect 8390 5210 8730 5296
rect 8390 5154 8462 5210
rect 8518 5154 8604 5210
rect 8660 5154 8730 5210
rect 8390 5068 8730 5154
rect 8390 5012 8462 5068
rect 8518 5012 8604 5068
rect 8660 5012 8730 5068
rect 8390 4926 8730 5012
rect 8390 4870 8462 4926
rect 8518 4870 8604 4926
rect 8660 4870 8730 4926
rect 8390 4784 8730 4870
rect 8390 4728 8462 4784
rect 8518 4728 8604 4784
rect 8660 4728 8730 4784
rect 8390 4642 8730 4728
rect 8390 4586 8462 4642
rect 8518 4586 8604 4642
rect 8660 4586 8730 4642
rect 8390 4500 8730 4586
rect 8390 4444 8462 4500
rect 8518 4444 8604 4500
rect 8660 4444 8730 4500
rect 8390 4358 8730 4444
rect 8390 4302 8462 4358
rect 8518 4302 8604 4358
rect 8660 4302 8730 4358
rect 8390 4216 8730 4302
rect 8390 4160 8462 4216
rect 8518 4160 8604 4216
rect 8660 4160 8730 4216
rect 8390 4074 8730 4160
rect 8390 4018 8462 4074
rect 8518 4018 8604 4074
rect 8660 4018 8730 4074
rect 8390 3932 8730 4018
rect 8390 3876 8462 3932
rect 8518 3876 8604 3932
rect 8660 3876 8730 3932
rect 8390 3790 8730 3876
rect 8390 3734 8462 3790
rect 8518 3734 8604 3790
rect 8660 3734 8730 3790
rect 8390 3648 8730 3734
rect 8390 3592 8462 3648
rect 8518 3592 8604 3648
rect 8660 3592 8730 3648
rect 8390 3506 8730 3592
rect 8390 3450 8462 3506
rect 8518 3450 8604 3506
rect 8660 3450 8730 3506
rect 8390 3364 8730 3450
rect 8390 3308 8462 3364
rect 8518 3308 8604 3364
rect 8660 3308 8730 3364
rect 8390 3222 8730 3308
rect 8390 3166 8462 3222
rect 8518 3166 8604 3222
rect 8660 3166 8730 3222
rect 8390 3080 8730 3166
rect 8390 3024 8462 3080
rect 8518 3024 8604 3080
rect 8660 3024 8730 3080
rect 8390 2938 8730 3024
rect 8390 2882 8462 2938
rect 8518 2882 8604 2938
rect 8660 2882 8730 2938
rect 8390 2796 8730 2882
rect 8390 2740 8462 2796
rect 8518 2740 8604 2796
rect 8660 2740 8730 2796
rect 8390 2654 8730 2740
rect 8390 2598 8462 2654
rect 8518 2598 8604 2654
rect 8660 2598 8730 2654
rect 8390 2512 8730 2598
rect 8390 2456 8462 2512
rect 8518 2456 8604 2512
rect 8660 2456 8730 2512
rect 8390 2370 8730 2456
rect 8390 2314 8462 2370
rect 8518 2314 8604 2370
rect 8660 2314 8730 2370
rect 8390 2228 8730 2314
rect 8390 2172 8462 2228
rect 8518 2172 8604 2228
rect 8660 2172 8730 2228
rect 8390 2086 8730 2172
rect 8390 2030 8462 2086
rect 8518 2030 8604 2086
rect 8660 2030 8730 2086
rect 8390 1944 8730 2030
rect 8390 1888 8462 1944
rect 8518 1888 8604 1944
rect 8660 1888 8730 1944
rect 8390 1802 8730 1888
rect 8390 1746 8462 1802
rect 8518 1746 8604 1802
rect 8660 1746 8730 1802
rect 8390 1660 8730 1746
rect 8390 1604 8462 1660
rect 8518 1604 8604 1660
rect 8660 1604 8730 1660
rect 8390 1518 8730 1604
rect 8390 1462 8462 1518
rect 8518 1462 8604 1518
rect 8660 1462 8730 1518
rect 8390 1376 8730 1462
rect 8390 1320 8462 1376
rect 8518 1320 8604 1376
rect 8660 1320 8730 1376
rect 8390 1234 8730 1320
rect 8390 1178 8462 1234
rect 8518 1178 8604 1234
rect 8660 1178 8730 1234
rect 8390 1092 8730 1178
rect 8390 1036 8462 1092
rect 8518 1036 8604 1092
rect 8660 1036 8730 1092
rect 8390 950 8730 1036
rect 8390 894 8462 950
rect 8518 894 8604 950
rect 8660 894 8730 950
rect 8390 808 8730 894
rect 8390 752 8462 808
rect 8518 752 8604 808
rect 8660 752 8730 808
rect 8390 666 8730 752
rect 8390 610 8462 666
rect 8518 610 8604 666
rect 8660 610 8730 666
rect 8390 524 8730 610
rect 8390 468 8462 524
rect 8518 468 8604 524
rect 8660 468 8730 524
rect 8390 458 8730 468
rect 8930 12310 9270 12320
rect 8930 12254 9004 12310
rect 9060 12254 9146 12310
rect 9202 12254 9270 12310
rect 8930 12168 9270 12254
rect 8930 12112 9004 12168
rect 9060 12112 9146 12168
rect 9202 12112 9270 12168
rect 8930 12026 9270 12112
rect 8930 11970 9004 12026
rect 9060 11970 9146 12026
rect 9202 11970 9270 12026
rect 8930 11884 9270 11970
rect 8930 11828 9004 11884
rect 9060 11828 9146 11884
rect 9202 11828 9270 11884
rect 8930 11742 9270 11828
rect 8930 11686 9004 11742
rect 9060 11686 9146 11742
rect 9202 11686 9270 11742
rect 8930 11600 9270 11686
rect 8930 11544 9004 11600
rect 9060 11544 9146 11600
rect 9202 11544 9270 11600
rect 8930 11458 9270 11544
rect 8930 11402 9004 11458
rect 9060 11402 9146 11458
rect 9202 11402 9270 11458
rect 8930 11316 9270 11402
rect 8930 11260 9004 11316
rect 9060 11260 9146 11316
rect 9202 11260 9270 11316
rect 8930 11174 9270 11260
rect 8930 11118 9004 11174
rect 9060 11118 9146 11174
rect 9202 11118 9270 11174
rect 8930 11032 9270 11118
rect 8930 10976 9004 11032
rect 9060 10976 9146 11032
rect 9202 10976 9270 11032
rect 8930 10890 9270 10976
rect 8930 10834 9004 10890
rect 9060 10834 9146 10890
rect 9202 10834 9270 10890
rect 8930 10748 9270 10834
rect 8930 10692 9004 10748
rect 9060 10692 9146 10748
rect 9202 10692 9270 10748
rect 8930 10606 9270 10692
rect 8930 10550 9004 10606
rect 9060 10550 9146 10606
rect 9202 10550 9270 10606
rect 8930 10464 9270 10550
rect 8930 10408 9004 10464
rect 9060 10408 9146 10464
rect 9202 10408 9270 10464
rect 8930 10322 9270 10408
rect 8930 10266 9004 10322
rect 9060 10266 9146 10322
rect 9202 10266 9270 10322
rect 8930 10180 9270 10266
rect 8930 10124 9004 10180
rect 9060 10124 9146 10180
rect 9202 10124 9270 10180
rect 8930 10038 9270 10124
rect 8930 9982 9004 10038
rect 9060 9982 9146 10038
rect 9202 9982 9270 10038
rect 8930 9896 9270 9982
rect 8930 9840 9004 9896
rect 9060 9840 9146 9896
rect 9202 9840 9270 9896
rect 8930 9754 9270 9840
rect 8930 9698 9004 9754
rect 9060 9698 9146 9754
rect 9202 9698 9270 9754
rect 8930 9612 9270 9698
rect 8930 9556 9004 9612
rect 9060 9556 9146 9612
rect 9202 9556 9270 9612
rect 8930 9470 9270 9556
rect 8930 9414 9004 9470
rect 9060 9414 9146 9470
rect 9202 9414 9270 9470
rect 8930 9328 9270 9414
rect 8930 9272 9004 9328
rect 9060 9272 9146 9328
rect 9202 9272 9270 9328
rect 8930 9186 9270 9272
rect 8930 9130 9004 9186
rect 9060 9130 9146 9186
rect 9202 9130 9270 9186
rect 8930 9044 9270 9130
rect 8930 8988 9004 9044
rect 9060 8988 9146 9044
rect 9202 8988 9270 9044
rect 8930 8902 9270 8988
rect 8930 8846 9004 8902
rect 9060 8846 9146 8902
rect 9202 8846 9270 8902
rect 8930 8760 9270 8846
rect 8930 8704 9004 8760
rect 9060 8704 9146 8760
rect 9202 8704 9270 8760
rect 8930 8618 9270 8704
rect 8930 8562 9004 8618
rect 9060 8562 9146 8618
rect 9202 8562 9270 8618
rect 8930 8476 9270 8562
rect 8930 8420 9004 8476
rect 9060 8420 9146 8476
rect 9202 8420 9270 8476
rect 8930 8334 9270 8420
rect 8930 8278 9004 8334
rect 9060 8278 9146 8334
rect 9202 8278 9270 8334
rect 8930 8192 9270 8278
rect 8930 8136 9004 8192
rect 9060 8136 9146 8192
rect 9202 8136 9270 8192
rect 8930 8050 9270 8136
rect 8930 7994 9004 8050
rect 9060 7994 9146 8050
rect 9202 7994 9270 8050
rect 8930 7908 9270 7994
rect 8930 7852 9004 7908
rect 9060 7852 9146 7908
rect 9202 7852 9270 7908
rect 8930 7766 9270 7852
rect 8930 7710 9004 7766
rect 9060 7710 9146 7766
rect 9202 7710 9270 7766
rect 8930 7624 9270 7710
rect 8930 7568 9004 7624
rect 9060 7568 9146 7624
rect 9202 7568 9270 7624
rect 8930 7482 9270 7568
rect 8930 7426 9004 7482
rect 9060 7426 9146 7482
rect 9202 7426 9270 7482
rect 8930 7340 9270 7426
rect 8930 7284 9004 7340
rect 9060 7284 9146 7340
rect 9202 7284 9270 7340
rect 8930 7198 9270 7284
rect 8930 7142 9004 7198
rect 9060 7142 9146 7198
rect 9202 7142 9270 7198
rect 8930 7056 9270 7142
rect 8930 7000 9004 7056
rect 9060 7000 9146 7056
rect 9202 7000 9270 7056
rect 8930 6914 9270 7000
rect 8930 6858 9004 6914
rect 9060 6858 9146 6914
rect 9202 6858 9270 6914
rect 8930 6772 9270 6858
rect 8930 6716 9004 6772
rect 9060 6716 9146 6772
rect 9202 6716 9270 6772
rect 8930 6630 9270 6716
rect 8930 6574 9004 6630
rect 9060 6574 9146 6630
rect 9202 6574 9270 6630
rect 8930 6488 9270 6574
rect 8930 6432 9004 6488
rect 9060 6432 9146 6488
rect 9202 6432 9270 6488
rect 8930 6346 9270 6432
rect 8930 6290 9004 6346
rect 9060 6290 9146 6346
rect 9202 6290 9270 6346
rect 8930 6204 9270 6290
rect 8930 6148 9004 6204
rect 9060 6148 9146 6204
rect 9202 6148 9270 6204
rect 8930 6062 9270 6148
rect 8930 6006 9004 6062
rect 9060 6006 9146 6062
rect 9202 6006 9270 6062
rect 8930 5920 9270 6006
rect 8930 5864 9004 5920
rect 9060 5864 9146 5920
rect 9202 5864 9270 5920
rect 8930 5778 9270 5864
rect 8930 5722 9004 5778
rect 9060 5722 9146 5778
rect 9202 5722 9270 5778
rect 8930 5636 9270 5722
rect 8930 5580 9004 5636
rect 9060 5580 9146 5636
rect 9202 5580 9270 5636
rect 8930 5494 9270 5580
rect 8930 5438 9004 5494
rect 9060 5438 9146 5494
rect 9202 5438 9270 5494
rect 8930 5352 9270 5438
rect 8930 5296 9004 5352
rect 9060 5296 9146 5352
rect 9202 5296 9270 5352
rect 8930 5210 9270 5296
rect 8930 5154 9004 5210
rect 9060 5154 9146 5210
rect 9202 5154 9270 5210
rect 8930 5068 9270 5154
rect 8930 5012 9004 5068
rect 9060 5012 9146 5068
rect 9202 5012 9270 5068
rect 8930 4926 9270 5012
rect 8930 4870 9004 4926
rect 9060 4870 9146 4926
rect 9202 4870 9270 4926
rect 8930 4784 9270 4870
rect 8930 4728 9004 4784
rect 9060 4728 9146 4784
rect 9202 4728 9270 4784
rect 8930 4642 9270 4728
rect 8930 4586 9004 4642
rect 9060 4586 9146 4642
rect 9202 4586 9270 4642
rect 8930 4500 9270 4586
rect 8930 4444 9004 4500
rect 9060 4444 9146 4500
rect 9202 4444 9270 4500
rect 8930 4358 9270 4444
rect 8930 4302 9004 4358
rect 9060 4302 9146 4358
rect 9202 4302 9270 4358
rect 8930 4216 9270 4302
rect 8930 4160 9004 4216
rect 9060 4160 9146 4216
rect 9202 4160 9270 4216
rect 8930 4074 9270 4160
rect 8930 4018 9004 4074
rect 9060 4018 9146 4074
rect 9202 4018 9270 4074
rect 8930 3932 9270 4018
rect 8930 3876 9004 3932
rect 9060 3876 9146 3932
rect 9202 3876 9270 3932
rect 8930 3790 9270 3876
rect 8930 3734 9004 3790
rect 9060 3734 9146 3790
rect 9202 3734 9270 3790
rect 8930 3648 9270 3734
rect 8930 3592 9004 3648
rect 9060 3592 9146 3648
rect 9202 3592 9270 3648
rect 8930 3506 9270 3592
rect 8930 3450 9004 3506
rect 9060 3450 9146 3506
rect 9202 3450 9270 3506
rect 8930 3364 9270 3450
rect 8930 3308 9004 3364
rect 9060 3308 9146 3364
rect 9202 3308 9270 3364
rect 8930 3222 9270 3308
rect 8930 3166 9004 3222
rect 9060 3166 9146 3222
rect 9202 3166 9270 3222
rect 8930 3080 9270 3166
rect 8930 3024 9004 3080
rect 9060 3024 9146 3080
rect 9202 3024 9270 3080
rect 8930 2938 9270 3024
rect 8930 2882 9004 2938
rect 9060 2882 9146 2938
rect 9202 2882 9270 2938
rect 8930 2796 9270 2882
rect 8930 2740 9004 2796
rect 9060 2740 9146 2796
rect 9202 2740 9270 2796
rect 8930 2654 9270 2740
rect 8930 2598 9004 2654
rect 9060 2598 9146 2654
rect 9202 2598 9270 2654
rect 8930 2512 9270 2598
rect 8930 2456 9004 2512
rect 9060 2456 9146 2512
rect 9202 2456 9270 2512
rect 8930 2370 9270 2456
rect 8930 2314 9004 2370
rect 9060 2314 9146 2370
rect 9202 2314 9270 2370
rect 8930 2228 9270 2314
rect 8930 2172 9004 2228
rect 9060 2172 9146 2228
rect 9202 2172 9270 2228
rect 8930 2086 9270 2172
rect 8930 2030 9004 2086
rect 9060 2030 9146 2086
rect 9202 2030 9270 2086
rect 8930 1944 9270 2030
rect 8930 1888 9004 1944
rect 9060 1888 9146 1944
rect 9202 1888 9270 1944
rect 8930 1802 9270 1888
rect 8930 1746 9004 1802
rect 9060 1746 9146 1802
rect 9202 1746 9270 1802
rect 8930 1660 9270 1746
rect 8930 1604 9004 1660
rect 9060 1604 9146 1660
rect 9202 1604 9270 1660
rect 8930 1518 9270 1604
rect 8930 1462 9004 1518
rect 9060 1462 9146 1518
rect 9202 1462 9270 1518
rect 8930 1376 9270 1462
rect 8930 1320 9004 1376
rect 9060 1320 9146 1376
rect 9202 1320 9270 1376
rect 8930 1234 9270 1320
rect 8930 1178 9004 1234
rect 9060 1178 9146 1234
rect 9202 1178 9270 1234
rect 8930 1092 9270 1178
rect 8930 1036 9004 1092
rect 9060 1036 9146 1092
rect 9202 1036 9270 1092
rect 8930 950 9270 1036
rect 8930 894 9004 950
rect 9060 894 9146 950
rect 9202 894 9270 950
rect 8930 808 9270 894
rect 8930 752 9004 808
rect 9060 752 9146 808
rect 9202 752 9270 808
rect 8930 666 9270 752
rect 8930 610 9004 666
rect 9060 610 9146 666
rect 9202 610 9270 666
rect 8930 524 9270 610
rect 8930 468 9004 524
rect 9060 468 9146 524
rect 9202 468 9270 524
rect 8930 458 9270 468
rect 9470 12310 9810 12320
rect 9470 12254 9547 12310
rect 9603 12254 9689 12310
rect 9745 12254 9810 12310
rect 9470 12168 9810 12254
rect 9470 12112 9547 12168
rect 9603 12112 9689 12168
rect 9745 12112 9810 12168
rect 9470 12026 9810 12112
rect 9470 11970 9547 12026
rect 9603 11970 9689 12026
rect 9745 11970 9810 12026
rect 9470 11884 9810 11970
rect 9470 11828 9547 11884
rect 9603 11828 9689 11884
rect 9745 11828 9810 11884
rect 9470 11742 9810 11828
rect 9470 11686 9547 11742
rect 9603 11686 9689 11742
rect 9745 11686 9810 11742
rect 9470 11600 9810 11686
rect 9470 11544 9547 11600
rect 9603 11544 9689 11600
rect 9745 11544 9810 11600
rect 9470 11458 9810 11544
rect 9470 11402 9547 11458
rect 9603 11402 9689 11458
rect 9745 11402 9810 11458
rect 9470 11316 9810 11402
rect 9470 11260 9547 11316
rect 9603 11260 9689 11316
rect 9745 11260 9810 11316
rect 9470 11174 9810 11260
rect 9470 11118 9547 11174
rect 9603 11118 9689 11174
rect 9745 11118 9810 11174
rect 9470 11032 9810 11118
rect 9470 10976 9547 11032
rect 9603 10976 9689 11032
rect 9745 10976 9810 11032
rect 9470 10890 9810 10976
rect 9470 10834 9547 10890
rect 9603 10834 9689 10890
rect 9745 10834 9810 10890
rect 9470 10748 9810 10834
rect 9470 10692 9547 10748
rect 9603 10692 9689 10748
rect 9745 10692 9810 10748
rect 9470 10606 9810 10692
rect 9470 10550 9547 10606
rect 9603 10550 9689 10606
rect 9745 10550 9810 10606
rect 9470 10464 9810 10550
rect 9470 10408 9547 10464
rect 9603 10408 9689 10464
rect 9745 10408 9810 10464
rect 9470 10322 9810 10408
rect 9470 10266 9547 10322
rect 9603 10266 9689 10322
rect 9745 10266 9810 10322
rect 9470 10180 9810 10266
rect 9470 10124 9547 10180
rect 9603 10124 9689 10180
rect 9745 10124 9810 10180
rect 9470 10038 9810 10124
rect 9470 9982 9547 10038
rect 9603 9982 9689 10038
rect 9745 9982 9810 10038
rect 9470 9896 9810 9982
rect 9470 9840 9547 9896
rect 9603 9840 9689 9896
rect 9745 9840 9810 9896
rect 9470 9754 9810 9840
rect 9470 9698 9547 9754
rect 9603 9698 9689 9754
rect 9745 9698 9810 9754
rect 9470 9612 9810 9698
rect 9470 9556 9547 9612
rect 9603 9556 9689 9612
rect 9745 9556 9810 9612
rect 9470 9470 9810 9556
rect 9470 9414 9547 9470
rect 9603 9414 9689 9470
rect 9745 9414 9810 9470
rect 9470 9328 9810 9414
rect 9470 9272 9547 9328
rect 9603 9272 9689 9328
rect 9745 9272 9810 9328
rect 9470 9186 9810 9272
rect 9470 9130 9547 9186
rect 9603 9130 9689 9186
rect 9745 9130 9810 9186
rect 9470 9044 9810 9130
rect 9470 8988 9547 9044
rect 9603 8988 9689 9044
rect 9745 8988 9810 9044
rect 9470 8902 9810 8988
rect 9470 8846 9547 8902
rect 9603 8846 9689 8902
rect 9745 8846 9810 8902
rect 9470 8760 9810 8846
rect 9470 8704 9547 8760
rect 9603 8704 9689 8760
rect 9745 8704 9810 8760
rect 9470 8618 9810 8704
rect 9470 8562 9547 8618
rect 9603 8562 9689 8618
rect 9745 8562 9810 8618
rect 9470 8476 9810 8562
rect 9470 8420 9547 8476
rect 9603 8420 9689 8476
rect 9745 8420 9810 8476
rect 9470 8334 9810 8420
rect 9470 8278 9547 8334
rect 9603 8278 9689 8334
rect 9745 8278 9810 8334
rect 9470 8192 9810 8278
rect 9470 8136 9547 8192
rect 9603 8136 9689 8192
rect 9745 8136 9810 8192
rect 9470 8050 9810 8136
rect 9470 7994 9547 8050
rect 9603 7994 9689 8050
rect 9745 7994 9810 8050
rect 9470 7908 9810 7994
rect 9470 7852 9547 7908
rect 9603 7852 9689 7908
rect 9745 7852 9810 7908
rect 9470 7766 9810 7852
rect 9470 7710 9547 7766
rect 9603 7710 9689 7766
rect 9745 7710 9810 7766
rect 9470 7624 9810 7710
rect 9470 7568 9547 7624
rect 9603 7568 9689 7624
rect 9745 7568 9810 7624
rect 9470 7482 9810 7568
rect 9470 7426 9547 7482
rect 9603 7426 9689 7482
rect 9745 7426 9810 7482
rect 9470 7340 9810 7426
rect 9470 7284 9547 7340
rect 9603 7284 9689 7340
rect 9745 7284 9810 7340
rect 9470 7198 9810 7284
rect 9470 7142 9547 7198
rect 9603 7142 9689 7198
rect 9745 7142 9810 7198
rect 9470 7056 9810 7142
rect 9470 7000 9547 7056
rect 9603 7000 9689 7056
rect 9745 7000 9810 7056
rect 9470 6914 9810 7000
rect 9470 6858 9547 6914
rect 9603 6858 9689 6914
rect 9745 6858 9810 6914
rect 9470 6772 9810 6858
rect 9470 6716 9547 6772
rect 9603 6716 9689 6772
rect 9745 6716 9810 6772
rect 9470 6630 9810 6716
rect 9470 6574 9547 6630
rect 9603 6574 9689 6630
rect 9745 6574 9810 6630
rect 9470 6488 9810 6574
rect 9470 6432 9547 6488
rect 9603 6432 9689 6488
rect 9745 6432 9810 6488
rect 9470 6346 9810 6432
rect 9470 6290 9547 6346
rect 9603 6290 9689 6346
rect 9745 6290 9810 6346
rect 9470 6204 9810 6290
rect 9470 6148 9547 6204
rect 9603 6148 9689 6204
rect 9745 6148 9810 6204
rect 9470 6062 9810 6148
rect 9470 6006 9547 6062
rect 9603 6006 9689 6062
rect 9745 6006 9810 6062
rect 9470 5920 9810 6006
rect 9470 5864 9547 5920
rect 9603 5864 9689 5920
rect 9745 5864 9810 5920
rect 9470 5778 9810 5864
rect 9470 5722 9547 5778
rect 9603 5722 9689 5778
rect 9745 5722 9810 5778
rect 9470 5636 9810 5722
rect 9470 5580 9547 5636
rect 9603 5580 9689 5636
rect 9745 5580 9810 5636
rect 9470 5494 9810 5580
rect 9470 5438 9547 5494
rect 9603 5438 9689 5494
rect 9745 5438 9810 5494
rect 9470 5352 9810 5438
rect 9470 5296 9547 5352
rect 9603 5296 9689 5352
rect 9745 5296 9810 5352
rect 9470 5210 9810 5296
rect 9470 5154 9547 5210
rect 9603 5154 9689 5210
rect 9745 5154 9810 5210
rect 9470 5068 9810 5154
rect 9470 5012 9547 5068
rect 9603 5012 9689 5068
rect 9745 5012 9810 5068
rect 9470 4926 9810 5012
rect 9470 4870 9547 4926
rect 9603 4870 9689 4926
rect 9745 4870 9810 4926
rect 9470 4784 9810 4870
rect 9470 4728 9547 4784
rect 9603 4728 9689 4784
rect 9745 4728 9810 4784
rect 9470 4642 9810 4728
rect 9470 4586 9547 4642
rect 9603 4586 9689 4642
rect 9745 4586 9810 4642
rect 9470 4500 9810 4586
rect 9470 4444 9547 4500
rect 9603 4444 9689 4500
rect 9745 4444 9810 4500
rect 9470 4358 9810 4444
rect 9470 4302 9547 4358
rect 9603 4302 9689 4358
rect 9745 4302 9810 4358
rect 9470 4216 9810 4302
rect 9470 4160 9547 4216
rect 9603 4160 9689 4216
rect 9745 4160 9810 4216
rect 9470 4074 9810 4160
rect 9470 4018 9547 4074
rect 9603 4018 9689 4074
rect 9745 4018 9810 4074
rect 9470 3932 9810 4018
rect 9470 3876 9547 3932
rect 9603 3876 9689 3932
rect 9745 3876 9810 3932
rect 9470 3790 9810 3876
rect 9470 3734 9547 3790
rect 9603 3734 9689 3790
rect 9745 3734 9810 3790
rect 9470 3648 9810 3734
rect 9470 3592 9547 3648
rect 9603 3592 9689 3648
rect 9745 3592 9810 3648
rect 9470 3506 9810 3592
rect 9470 3450 9547 3506
rect 9603 3450 9689 3506
rect 9745 3450 9810 3506
rect 9470 3364 9810 3450
rect 9470 3308 9547 3364
rect 9603 3308 9689 3364
rect 9745 3308 9810 3364
rect 9470 3222 9810 3308
rect 9470 3166 9547 3222
rect 9603 3166 9689 3222
rect 9745 3166 9810 3222
rect 9470 3080 9810 3166
rect 9470 3024 9547 3080
rect 9603 3024 9689 3080
rect 9745 3024 9810 3080
rect 9470 2938 9810 3024
rect 9470 2882 9547 2938
rect 9603 2882 9689 2938
rect 9745 2882 9810 2938
rect 9470 2796 9810 2882
rect 9470 2740 9547 2796
rect 9603 2740 9689 2796
rect 9745 2740 9810 2796
rect 9470 2654 9810 2740
rect 9470 2598 9547 2654
rect 9603 2598 9689 2654
rect 9745 2598 9810 2654
rect 9470 2512 9810 2598
rect 9470 2456 9547 2512
rect 9603 2456 9689 2512
rect 9745 2456 9810 2512
rect 9470 2370 9810 2456
rect 9470 2314 9547 2370
rect 9603 2314 9689 2370
rect 9745 2314 9810 2370
rect 9470 2228 9810 2314
rect 9470 2172 9547 2228
rect 9603 2172 9689 2228
rect 9745 2172 9810 2228
rect 9470 2086 9810 2172
rect 9470 2030 9547 2086
rect 9603 2030 9689 2086
rect 9745 2030 9810 2086
rect 9470 1944 9810 2030
rect 9470 1888 9547 1944
rect 9603 1888 9689 1944
rect 9745 1888 9810 1944
rect 9470 1802 9810 1888
rect 9470 1746 9547 1802
rect 9603 1746 9689 1802
rect 9745 1746 9810 1802
rect 9470 1660 9810 1746
rect 9470 1604 9547 1660
rect 9603 1604 9689 1660
rect 9745 1604 9810 1660
rect 9470 1518 9810 1604
rect 9470 1462 9547 1518
rect 9603 1462 9689 1518
rect 9745 1462 9810 1518
rect 9470 1376 9810 1462
rect 9470 1320 9547 1376
rect 9603 1320 9689 1376
rect 9745 1320 9810 1376
rect 9470 1234 9810 1320
rect 9470 1178 9547 1234
rect 9603 1178 9689 1234
rect 9745 1178 9810 1234
rect 9470 1092 9810 1178
rect 9470 1036 9547 1092
rect 9603 1036 9689 1092
rect 9745 1036 9810 1092
rect 9470 950 9810 1036
rect 9470 894 9547 950
rect 9603 894 9689 950
rect 9745 894 9810 950
rect 9470 808 9810 894
rect 9470 752 9547 808
rect 9603 752 9689 808
rect 9745 752 9810 808
rect 9470 666 9810 752
rect 9470 610 9547 666
rect 9603 610 9689 666
rect 9745 610 9810 666
rect 9470 524 9810 610
rect 9470 468 9547 524
rect 9603 468 9689 524
rect 9745 468 9810 524
rect 9470 458 9810 468
rect 10010 12310 10350 12320
rect 10010 12254 10081 12310
rect 10137 12254 10223 12310
rect 10279 12254 10350 12310
rect 10010 12168 10350 12254
rect 10010 12112 10081 12168
rect 10137 12112 10223 12168
rect 10279 12112 10350 12168
rect 10010 12026 10350 12112
rect 10010 11970 10081 12026
rect 10137 11970 10223 12026
rect 10279 11970 10350 12026
rect 10010 11884 10350 11970
rect 10010 11828 10081 11884
rect 10137 11828 10223 11884
rect 10279 11828 10350 11884
rect 10010 11742 10350 11828
rect 10010 11686 10081 11742
rect 10137 11686 10223 11742
rect 10279 11686 10350 11742
rect 10010 11600 10350 11686
rect 10010 11544 10081 11600
rect 10137 11544 10223 11600
rect 10279 11544 10350 11600
rect 10010 11458 10350 11544
rect 10010 11402 10081 11458
rect 10137 11402 10223 11458
rect 10279 11402 10350 11458
rect 10010 11316 10350 11402
rect 10010 11260 10081 11316
rect 10137 11260 10223 11316
rect 10279 11260 10350 11316
rect 10010 11174 10350 11260
rect 10010 11118 10081 11174
rect 10137 11118 10223 11174
rect 10279 11118 10350 11174
rect 10010 11032 10350 11118
rect 10010 10976 10081 11032
rect 10137 10976 10223 11032
rect 10279 10976 10350 11032
rect 10010 10890 10350 10976
rect 10010 10834 10081 10890
rect 10137 10834 10223 10890
rect 10279 10834 10350 10890
rect 10010 10748 10350 10834
rect 10010 10692 10081 10748
rect 10137 10692 10223 10748
rect 10279 10692 10350 10748
rect 10010 10606 10350 10692
rect 10010 10550 10081 10606
rect 10137 10550 10223 10606
rect 10279 10550 10350 10606
rect 10010 10464 10350 10550
rect 10010 10408 10081 10464
rect 10137 10408 10223 10464
rect 10279 10408 10350 10464
rect 10010 10322 10350 10408
rect 10010 10266 10081 10322
rect 10137 10266 10223 10322
rect 10279 10266 10350 10322
rect 10010 10180 10350 10266
rect 10010 10124 10081 10180
rect 10137 10124 10223 10180
rect 10279 10124 10350 10180
rect 10010 10038 10350 10124
rect 10010 9982 10081 10038
rect 10137 9982 10223 10038
rect 10279 9982 10350 10038
rect 10010 9896 10350 9982
rect 10010 9840 10081 9896
rect 10137 9840 10223 9896
rect 10279 9840 10350 9896
rect 10010 9754 10350 9840
rect 10010 9698 10081 9754
rect 10137 9698 10223 9754
rect 10279 9698 10350 9754
rect 10010 9612 10350 9698
rect 10010 9556 10081 9612
rect 10137 9556 10223 9612
rect 10279 9556 10350 9612
rect 10010 9470 10350 9556
rect 10010 9414 10081 9470
rect 10137 9414 10223 9470
rect 10279 9414 10350 9470
rect 10010 9328 10350 9414
rect 10010 9272 10081 9328
rect 10137 9272 10223 9328
rect 10279 9272 10350 9328
rect 10010 9186 10350 9272
rect 10010 9130 10081 9186
rect 10137 9130 10223 9186
rect 10279 9130 10350 9186
rect 10010 9044 10350 9130
rect 10010 8988 10081 9044
rect 10137 8988 10223 9044
rect 10279 8988 10350 9044
rect 10010 8902 10350 8988
rect 10010 8846 10081 8902
rect 10137 8846 10223 8902
rect 10279 8846 10350 8902
rect 10010 8760 10350 8846
rect 10010 8704 10081 8760
rect 10137 8704 10223 8760
rect 10279 8704 10350 8760
rect 10010 8618 10350 8704
rect 10010 8562 10081 8618
rect 10137 8562 10223 8618
rect 10279 8562 10350 8618
rect 10010 8476 10350 8562
rect 10010 8420 10081 8476
rect 10137 8420 10223 8476
rect 10279 8420 10350 8476
rect 10010 8334 10350 8420
rect 10010 8278 10081 8334
rect 10137 8278 10223 8334
rect 10279 8278 10350 8334
rect 10010 8192 10350 8278
rect 10010 8136 10081 8192
rect 10137 8136 10223 8192
rect 10279 8136 10350 8192
rect 10010 8050 10350 8136
rect 10010 7994 10081 8050
rect 10137 7994 10223 8050
rect 10279 7994 10350 8050
rect 10010 7908 10350 7994
rect 10010 7852 10081 7908
rect 10137 7852 10223 7908
rect 10279 7852 10350 7908
rect 10010 7766 10350 7852
rect 10010 7710 10081 7766
rect 10137 7710 10223 7766
rect 10279 7710 10350 7766
rect 10010 7624 10350 7710
rect 10010 7568 10081 7624
rect 10137 7568 10223 7624
rect 10279 7568 10350 7624
rect 10010 7482 10350 7568
rect 10010 7426 10081 7482
rect 10137 7426 10223 7482
rect 10279 7426 10350 7482
rect 10010 7340 10350 7426
rect 10010 7284 10081 7340
rect 10137 7284 10223 7340
rect 10279 7284 10350 7340
rect 10010 7198 10350 7284
rect 10010 7142 10081 7198
rect 10137 7142 10223 7198
rect 10279 7142 10350 7198
rect 10010 7056 10350 7142
rect 10010 7000 10081 7056
rect 10137 7000 10223 7056
rect 10279 7000 10350 7056
rect 10010 6914 10350 7000
rect 10010 6858 10081 6914
rect 10137 6858 10223 6914
rect 10279 6858 10350 6914
rect 10010 6772 10350 6858
rect 10010 6716 10081 6772
rect 10137 6716 10223 6772
rect 10279 6716 10350 6772
rect 10010 6630 10350 6716
rect 10010 6574 10081 6630
rect 10137 6574 10223 6630
rect 10279 6574 10350 6630
rect 10010 6488 10350 6574
rect 10010 6432 10081 6488
rect 10137 6432 10223 6488
rect 10279 6432 10350 6488
rect 10010 6346 10350 6432
rect 10010 6290 10081 6346
rect 10137 6290 10223 6346
rect 10279 6290 10350 6346
rect 10010 6204 10350 6290
rect 10010 6148 10081 6204
rect 10137 6148 10223 6204
rect 10279 6148 10350 6204
rect 10010 6062 10350 6148
rect 10010 6006 10081 6062
rect 10137 6006 10223 6062
rect 10279 6006 10350 6062
rect 10010 5920 10350 6006
rect 10010 5864 10081 5920
rect 10137 5864 10223 5920
rect 10279 5864 10350 5920
rect 10010 5778 10350 5864
rect 10010 5722 10081 5778
rect 10137 5722 10223 5778
rect 10279 5722 10350 5778
rect 10010 5636 10350 5722
rect 10010 5580 10081 5636
rect 10137 5580 10223 5636
rect 10279 5580 10350 5636
rect 10010 5494 10350 5580
rect 10010 5438 10081 5494
rect 10137 5438 10223 5494
rect 10279 5438 10350 5494
rect 10010 5352 10350 5438
rect 10010 5296 10081 5352
rect 10137 5296 10223 5352
rect 10279 5296 10350 5352
rect 10010 5210 10350 5296
rect 10010 5154 10081 5210
rect 10137 5154 10223 5210
rect 10279 5154 10350 5210
rect 10010 5068 10350 5154
rect 10010 5012 10081 5068
rect 10137 5012 10223 5068
rect 10279 5012 10350 5068
rect 10010 4926 10350 5012
rect 10010 4870 10081 4926
rect 10137 4870 10223 4926
rect 10279 4870 10350 4926
rect 10010 4784 10350 4870
rect 10010 4728 10081 4784
rect 10137 4728 10223 4784
rect 10279 4728 10350 4784
rect 10010 4642 10350 4728
rect 10010 4586 10081 4642
rect 10137 4586 10223 4642
rect 10279 4586 10350 4642
rect 10010 4500 10350 4586
rect 10010 4444 10081 4500
rect 10137 4444 10223 4500
rect 10279 4444 10350 4500
rect 10010 4358 10350 4444
rect 10010 4302 10081 4358
rect 10137 4302 10223 4358
rect 10279 4302 10350 4358
rect 10010 4216 10350 4302
rect 10010 4160 10081 4216
rect 10137 4160 10223 4216
rect 10279 4160 10350 4216
rect 10010 4074 10350 4160
rect 10010 4018 10081 4074
rect 10137 4018 10223 4074
rect 10279 4018 10350 4074
rect 10010 3932 10350 4018
rect 10010 3876 10081 3932
rect 10137 3876 10223 3932
rect 10279 3876 10350 3932
rect 10010 3790 10350 3876
rect 10010 3734 10081 3790
rect 10137 3734 10223 3790
rect 10279 3734 10350 3790
rect 10010 3648 10350 3734
rect 10010 3592 10081 3648
rect 10137 3592 10223 3648
rect 10279 3592 10350 3648
rect 10010 3506 10350 3592
rect 10010 3450 10081 3506
rect 10137 3450 10223 3506
rect 10279 3450 10350 3506
rect 10010 3364 10350 3450
rect 10010 3308 10081 3364
rect 10137 3308 10223 3364
rect 10279 3308 10350 3364
rect 10010 3222 10350 3308
rect 10010 3166 10081 3222
rect 10137 3166 10223 3222
rect 10279 3166 10350 3222
rect 10010 3080 10350 3166
rect 10010 3024 10081 3080
rect 10137 3024 10223 3080
rect 10279 3024 10350 3080
rect 10010 2938 10350 3024
rect 10010 2882 10081 2938
rect 10137 2882 10223 2938
rect 10279 2882 10350 2938
rect 10010 2796 10350 2882
rect 10010 2740 10081 2796
rect 10137 2740 10223 2796
rect 10279 2740 10350 2796
rect 10010 2654 10350 2740
rect 10010 2598 10081 2654
rect 10137 2598 10223 2654
rect 10279 2598 10350 2654
rect 10010 2512 10350 2598
rect 10010 2456 10081 2512
rect 10137 2456 10223 2512
rect 10279 2456 10350 2512
rect 10010 2370 10350 2456
rect 10010 2314 10081 2370
rect 10137 2314 10223 2370
rect 10279 2314 10350 2370
rect 10010 2228 10350 2314
rect 10010 2172 10081 2228
rect 10137 2172 10223 2228
rect 10279 2172 10350 2228
rect 10010 2086 10350 2172
rect 10010 2030 10081 2086
rect 10137 2030 10223 2086
rect 10279 2030 10350 2086
rect 10010 1944 10350 2030
rect 10010 1888 10081 1944
rect 10137 1888 10223 1944
rect 10279 1888 10350 1944
rect 10010 1802 10350 1888
rect 10010 1746 10081 1802
rect 10137 1746 10223 1802
rect 10279 1746 10350 1802
rect 10010 1660 10350 1746
rect 10010 1604 10081 1660
rect 10137 1604 10223 1660
rect 10279 1604 10350 1660
rect 10010 1518 10350 1604
rect 10010 1462 10081 1518
rect 10137 1462 10223 1518
rect 10279 1462 10350 1518
rect 10010 1376 10350 1462
rect 10010 1320 10081 1376
rect 10137 1320 10223 1376
rect 10279 1320 10350 1376
rect 10010 1234 10350 1320
rect 10010 1178 10081 1234
rect 10137 1178 10223 1234
rect 10279 1178 10350 1234
rect 10010 1092 10350 1178
rect 10010 1036 10081 1092
rect 10137 1036 10223 1092
rect 10279 1036 10350 1092
rect 10010 950 10350 1036
rect 10010 894 10081 950
rect 10137 894 10223 950
rect 10279 894 10350 950
rect 10010 808 10350 894
rect 10010 752 10081 808
rect 10137 752 10223 808
rect 10279 752 10350 808
rect 10010 666 10350 752
rect 10010 610 10081 666
rect 10137 610 10223 666
rect 10279 610 10350 666
rect 10010 524 10350 610
rect 10010 468 10081 524
rect 10137 468 10223 524
rect 10279 468 10350 524
rect 10010 458 10350 468
rect 10550 12310 10890 12320
rect 10550 12254 10622 12310
rect 10678 12254 10764 12310
rect 10820 12254 10890 12310
rect 10550 12168 10890 12254
rect 10550 12112 10622 12168
rect 10678 12112 10764 12168
rect 10820 12112 10890 12168
rect 10550 12026 10890 12112
rect 10550 11970 10622 12026
rect 10678 11970 10764 12026
rect 10820 11970 10890 12026
rect 10550 11884 10890 11970
rect 10550 11828 10622 11884
rect 10678 11828 10764 11884
rect 10820 11828 10890 11884
rect 10550 11742 10890 11828
rect 10550 11686 10622 11742
rect 10678 11686 10764 11742
rect 10820 11686 10890 11742
rect 10550 11600 10890 11686
rect 10550 11544 10622 11600
rect 10678 11544 10764 11600
rect 10820 11544 10890 11600
rect 10550 11458 10890 11544
rect 10550 11402 10622 11458
rect 10678 11402 10764 11458
rect 10820 11402 10890 11458
rect 10550 11316 10890 11402
rect 10550 11260 10622 11316
rect 10678 11260 10764 11316
rect 10820 11260 10890 11316
rect 10550 11174 10890 11260
rect 10550 11118 10622 11174
rect 10678 11118 10764 11174
rect 10820 11118 10890 11174
rect 10550 11032 10890 11118
rect 10550 10976 10622 11032
rect 10678 10976 10764 11032
rect 10820 10976 10890 11032
rect 10550 10890 10890 10976
rect 10550 10834 10622 10890
rect 10678 10834 10764 10890
rect 10820 10834 10890 10890
rect 10550 10748 10890 10834
rect 10550 10692 10622 10748
rect 10678 10692 10764 10748
rect 10820 10692 10890 10748
rect 10550 10606 10890 10692
rect 10550 10550 10622 10606
rect 10678 10550 10764 10606
rect 10820 10550 10890 10606
rect 10550 10464 10890 10550
rect 10550 10408 10622 10464
rect 10678 10408 10764 10464
rect 10820 10408 10890 10464
rect 10550 10322 10890 10408
rect 10550 10266 10622 10322
rect 10678 10266 10764 10322
rect 10820 10266 10890 10322
rect 10550 10180 10890 10266
rect 10550 10124 10622 10180
rect 10678 10124 10764 10180
rect 10820 10124 10890 10180
rect 10550 10038 10890 10124
rect 10550 9982 10622 10038
rect 10678 9982 10764 10038
rect 10820 9982 10890 10038
rect 10550 9896 10890 9982
rect 10550 9840 10622 9896
rect 10678 9840 10764 9896
rect 10820 9840 10890 9896
rect 10550 9754 10890 9840
rect 10550 9698 10622 9754
rect 10678 9698 10764 9754
rect 10820 9698 10890 9754
rect 10550 9612 10890 9698
rect 10550 9556 10622 9612
rect 10678 9556 10764 9612
rect 10820 9556 10890 9612
rect 10550 9470 10890 9556
rect 10550 9414 10622 9470
rect 10678 9414 10764 9470
rect 10820 9414 10890 9470
rect 10550 9328 10890 9414
rect 10550 9272 10622 9328
rect 10678 9272 10764 9328
rect 10820 9272 10890 9328
rect 10550 9186 10890 9272
rect 10550 9130 10622 9186
rect 10678 9130 10764 9186
rect 10820 9130 10890 9186
rect 10550 9044 10890 9130
rect 10550 8988 10622 9044
rect 10678 8988 10764 9044
rect 10820 8988 10890 9044
rect 10550 8902 10890 8988
rect 10550 8846 10622 8902
rect 10678 8846 10764 8902
rect 10820 8846 10890 8902
rect 10550 8760 10890 8846
rect 10550 8704 10622 8760
rect 10678 8704 10764 8760
rect 10820 8704 10890 8760
rect 10550 8618 10890 8704
rect 10550 8562 10622 8618
rect 10678 8562 10764 8618
rect 10820 8562 10890 8618
rect 10550 8476 10890 8562
rect 10550 8420 10622 8476
rect 10678 8420 10764 8476
rect 10820 8420 10890 8476
rect 10550 8334 10890 8420
rect 10550 8278 10622 8334
rect 10678 8278 10764 8334
rect 10820 8278 10890 8334
rect 10550 8192 10890 8278
rect 10550 8136 10622 8192
rect 10678 8136 10764 8192
rect 10820 8136 10890 8192
rect 10550 8050 10890 8136
rect 10550 7994 10622 8050
rect 10678 7994 10764 8050
rect 10820 7994 10890 8050
rect 10550 7908 10890 7994
rect 10550 7852 10622 7908
rect 10678 7852 10764 7908
rect 10820 7852 10890 7908
rect 10550 7766 10890 7852
rect 10550 7710 10622 7766
rect 10678 7710 10764 7766
rect 10820 7710 10890 7766
rect 10550 7624 10890 7710
rect 10550 7568 10622 7624
rect 10678 7568 10764 7624
rect 10820 7568 10890 7624
rect 10550 7482 10890 7568
rect 10550 7426 10622 7482
rect 10678 7426 10764 7482
rect 10820 7426 10890 7482
rect 10550 7340 10890 7426
rect 10550 7284 10622 7340
rect 10678 7284 10764 7340
rect 10820 7284 10890 7340
rect 10550 7198 10890 7284
rect 10550 7142 10622 7198
rect 10678 7142 10764 7198
rect 10820 7142 10890 7198
rect 10550 7056 10890 7142
rect 10550 7000 10622 7056
rect 10678 7000 10764 7056
rect 10820 7000 10890 7056
rect 10550 6914 10890 7000
rect 10550 6858 10622 6914
rect 10678 6858 10764 6914
rect 10820 6858 10890 6914
rect 10550 6772 10890 6858
rect 10550 6716 10622 6772
rect 10678 6716 10764 6772
rect 10820 6716 10890 6772
rect 10550 6630 10890 6716
rect 10550 6574 10622 6630
rect 10678 6574 10764 6630
rect 10820 6574 10890 6630
rect 10550 6488 10890 6574
rect 10550 6432 10622 6488
rect 10678 6432 10764 6488
rect 10820 6432 10890 6488
rect 10550 6346 10890 6432
rect 10550 6290 10622 6346
rect 10678 6290 10764 6346
rect 10820 6290 10890 6346
rect 10550 6204 10890 6290
rect 10550 6148 10622 6204
rect 10678 6148 10764 6204
rect 10820 6148 10890 6204
rect 10550 6062 10890 6148
rect 10550 6006 10622 6062
rect 10678 6006 10764 6062
rect 10820 6006 10890 6062
rect 10550 5920 10890 6006
rect 10550 5864 10622 5920
rect 10678 5864 10764 5920
rect 10820 5864 10890 5920
rect 10550 5778 10890 5864
rect 10550 5722 10622 5778
rect 10678 5722 10764 5778
rect 10820 5722 10890 5778
rect 10550 5636 10890 5722
rect 10550 5580 10622 5636
rect 10678 5580 10764 5636
rect 10820 5580 10890 5636
rect 10550 5494 10890 5580
rect 10550 5438 10622 5494
rect 10678 5438 10764 5494
rect 10820 5438 10890 5494
rect 10550 5352 10890 5438
rect 10550 5296 10622 5352
rect 10678 5296 10764 5352
rect 10820 5296 10890 5352
rect 10550 5210 10890 5296
rect 10550 5154 10622 5210
rect 10678 5154 10764 5210
rect 10820 5154 10890 5210
rect 10550 5068 10890 5154
rect 10550 5012 10622 5068
rect 10678 5012 10764 5068
rect 10820 5012 10890 5068
rect 10550 4926 10890 5012
rect 10550 4870 10622 4926
rect 10678 4870 10764 4926
rect 10820 4870 10890 4926
rect 10550 4784 10890 4870
rect 10550 4728 10622 4784
rect 10678 4728 10764 4784
rect 10820 4728 10890 4784
rect 10550 4642 10890 4728
rect 10550 4586 10622 4642
rect 10678 4586 10764 4642
rect 10820 4586 10890 4642
rect 10550 4500 10890 4586
rect 10550 4444 10622 4500
rect 10678 4444 10764 4500
rect 10820 4444 10890 4500
rect 10550 4358 10890 4444
rect 10550 4302 10622 4358
rect 10678 4302 10764 4358
rect 10820 4302 10890 4358
rect 10550 4216 10890 4302
rect 10550 4160 10622 4216
rect 10678 4160 10764 4216
rect 10820 4160 10890 4216
rect 10550 4074 10890 4160
rect 10550 4018 10622 4074
rect 10678 4018 10764 4074
rect 10820 4018 10890 4074
rect 10550 3932 10890 4018
rect 10550 3876 10622 3932
rect 10678 3876 10764 3932
rect 10820 3876 10890 3932
rect 10550 3790 10890 3876
rect 10550 3734 10622 3790
rect 10678 3734 10764 3790
rect 10820 3734 10890 3790
rect 10550 3648 10890 3734
rect 10550 3592 10622 3648
rect 10678 3592 10764 3648
rect 10820 3592 10890 3648
rect 10550 3506 10890 3592
rect 10550 3450 10622 3506
rect 10678 3450 10764 3506
rect 10820 3450 10890 3506
rect 10550 3364 10890 3450
rect 10550 3308 10622 3364
rect 10678 3308 10764 3364
rect 10820 3308 10890 3364
rect 10550 3222 10890 3308
rect 10550 3166 10622 3222
rect 10678 3166 10764 3222
rect 10820 3166 10890 3222
rect 10550 3080 10890 3166
rect 10550 3024 10622 3080
rect 10678 3024 10764 3080
rect 10820 3024 10890 3080
rect 10550 2938 10890 3024
rect 10550 2882 10622 2938
rect 10678 2882 10764 2938
rect 10820 2882 10890 2938
rect 10550 2796 10890 2882
rect 10550 2740 10622 2796
rect 10678 2740 10764 2796
rect 10820 2740 10890 2796
rect 10550 2654 10890 2740
rect 10550 2598 10622 2654
rect 10678 2598 10764 2654
rect 10820 2598 10890 2654
rect 10550 2512 10890 2598
rect 10550 2456 10622 2512
rect 10678 2456 10764 2512
rect 10820 2456 10890 2512
rect 10550 2370 10890 2456
rect 10550 2314 10622 2370
rect 10678 2314 10764 2370
rect 10820 2314 10890 2370
rect 10550 2228 10890 2314
rect 10550 2172 10622 2228
rect 10678 2172 10764 2228
rect 10820 2172 10890 2228
rect 10550 2086 10890 2172
rect 10550 2030 10622 2086
rect 10678 2030 10764 2086
rect 10820 2030 10890 2086
rect 10550 1944 10890 2030
rect 10550 1888 10622 1944
rect 10678 1888 10764 1944
rect 10820 1888 10890 1944
rect 10550 1802 10890 1888
rect 10550 1746 10622 1802
rect 10678 1746 10764 1802
rect 10820 1746 10890 1802
rect 10550 1660 10890 1746
rect 10550 1604 10622 1660
rect 10678 1604 10764 1660
rect 10820 1604 10890 1660
rect 10550 1518 10890 1604
rect 10550 1462 10622 1518
rect 10678 1462 10764 1518
rect 10820 1462 10890 1518
rect 10550 1376 10890 1462
rect 10550 1320 10622 1376
rect 10678 1320 10764 1376
rect 10820 1320 10890 1376
rect 10550 1234 10890 1320
rect 10550 1178 10622 1234
rect 10678 1178 10764 1234
rect 10820 1178 10890 1234
rect 10550 1092 10890 1178
rect 10550 1036 10622 1092
rect 10678 1036 10764 1092
rect 10820 1036 10890 1092
rect 10550 950 10890 1036
rect 10550 894 10622 950
rect 10678 894 10764 950
rect 10820 894 10890 950
rect 10550 808 10890 894
rect 10550 752 10622 808
rect 10678 752 10764 808
rect 10820 752 10890 808
rect 10550 666 10890 752
rect 10550 610 10622 666
rect 10678 610 10764 666
rect 10820 610 10890 666
rect 10550 524 10890 610
rect 10550 468 10622 524
rect 10678 468 10764 524
rect 10820 468 10890 524
rect 10550 458 10890 468
rect 11090 12310 11430 12320
rect 11090 12254 11162 12310
rect 11218 12254 11304 12310
rect 11360 12254 11430 12310
rect 11090 12168 11430 12254
rect 11090 12112 11162 12168
rect 11218 12112 11304 12168
rect 11360 12112 11430 12168
rect 11090 12026 11430 12112
rect 11090 11970 11162 12026
rect 11218 11970 11304 12026
rect 11360 11970 11430 12026
rect 11090 11884 11430 11970
rect 11090 11828 11162 11884
rect 11218 11828 11304 11884
rect 11360 11828 11430 11884
rect 11090 11742 11430 11828
rect 11090 11686 11162 11742
rect 11218 11686 11304 11742
rect 11360 11686 11430 11742
rect 11090 11600 11430 11686
rect 11090 11544 11162 11600
rect 11218 11544 11304 11600
rect 11360 11544 11430 11600
rect 11090 11458 11430 11544
rect 11090 11402 11162 11458
rect 11218 11402 11304 11458
rect 11360 11402 11430 11458
rect 11090 11316 11430 11402
rect 11090 11260 11162 11316
rect 11218 11260 11304 11316
rect 11360 11260 11430 11316
rect 11090 11174 11430 11260
rect 11090 11118 11162 11174
rect 11218 11118 11304 11174
rect 11360 11118 11430 11174
rect 11090 11032 11430 11118
rect 11090 10976 11162 11032
rect 11218 10976 11304 11032
rect 11360 10976 11430 11032
rect 11090 10890 11430 10976
rect 11090 10834 11162 10890
rect 11218 10834 11304 10890
rect 11360 10834 11430 10890
rect 11090 10748 11430 10834
rect 11090 10692 11162 10748
rect 11218 10692 11304 10748
rect 11360 10692 11430 10748
rect 11090 10606 11430 10692
rect 11090 10550 11162 10606
rect 11218 10550 11304 10606
rect 11360 10550 11430 10606
rect 11090 10464 11430 10550
rect 11090 10408 11162 10464
rect 11218 10408 11304 10464
rect 11360 10408 11430 10464
rect 11090 10322 11430 10408
rect 11090 10266 11162 10322
rect 11218 10266 11304 10322
rect 11360 10266 11430 10322
rect 11090 10180 11430 10266
rect 11090 10124 11162 10180
rect 11218 10124 11304 10180
rect 11360 10124 11430 10180
rect 11090 10038 11430 10124
rect 11090 9982 11162 10038
rect 11218 9982 11304 10038
rect 11360 9982 11430 10038
rect 11090 9896 11430 9982
rect 11090 9840 11162 9896
rect 11218 9840 11304 9896
rect 11360 9840 11430 9896
rect 11090 9754 11430 9840
rect 11090 9698 11162 9754
rect 11218 9698 11304 9754
rect 11360 9698 11430 9754
rect 11090 9612 11430 9698
rect 11090 9556 11162 9612
rect 11218 9556 11304 9612
rect 11360 9556 11430 9612
rect 11090 9470 11430 9556
rect 11090 9414 11162 9470
rect 11218 9414 11304 9470
rect 11360 9414 11430 9470
rect 11090 9328 11430 9414
rect 11090 9272 11162 9328
rect 11218 9272 11304 9328
rect 11360 9272 11430 9328
rect 11090 9186 11430 9272
rect 11090 9130 11162 9186
rect 11218 9130 11304 9186
rect 11360 9130 11430 9186
rect 11090 9044 11430 9130
rect 11090 8988 11162 9044
rect 11218 8988 11304 9044
rect 11360 8988 11430 9044
rect 11090 8902 11430 8988
rect 11090 8846 11162 8902
rect 11218 8846 11304 8902
rect 11360 8846 11430 8902
rect 11090 8760 11430 8846
rect 11090 8704 11162 8760
rect 11218 8704 11304 8760
rect 11360 8704 11430 8760
rect 11090 8618 11430 8704
rect 11090 8562 11162 8618
rect 11218 8562 11304 8618
rect 11360 8562 11430 8618
rect 11090 8476 11430 8562
rect 11090 8420 11162 8476
rect 11218 8420 11304 8476
rect 11360 8420 11430 8476
rect 11090 8334 11430 8420
rect 11090 8278 11162 8334
rect 11218 8278 11304 8334
rect 11360 8278 11430 8334
rect 11090 8192 11430 8278
rect 11090 8136 11162 8192
rect 11218 8136 11304 8192
rect 11360 8136 11430 8192
rect 11090 8050 11430 8136
rect 11090 7994 11162 8050
rect 11218 7994 11304 8050
rect 11360 7994 11430 8050
rect 11090 7908 11430 7994
rect 11090 7852 11162 7908
rect 11218 7852 11304 7908
rect 11360 7852 11430 7908
rect 11090 7766 11430 7852
rect 11090 7710 11162 7766
rect 11218 7710 11304 7766
rect 11360 7710 11430 7766
rect 11090 7624 11430 7710
rect 11090 7568 11162 7624
rect 11218 7568 11304 7624
rect 11360 7568 11430 7624
rect 11090 7482 11430 7568
rect 11090 7426 11162 7482
rect 11218 7426 11304 7482
rect 11360 7426 11430 7482
rect 11090 7340 11430 7426
rect 11090 7284 11162 7340
rect 11218 7284 11304 7340
rect 11360 7284 11430 7340
rect 11090 7198 11430 7284
rect 11090 7142 11162 7198
rect 11218 7142 11304 7198
rect 11360 7142 11430 7198
rect 11090 7056 11430 7142
rect 11090 7000 11162 7056
rect 11218 7000 11304 7056
rect 11360 7000 11430 7056
rect 11090 6914 11430 7000
rect 11090 6858 11162 6914
rect 11218 6858 11304 6914
rect 11360 6858 11430 6914
rect 11090 6772 11430 6858
rect 11090 6716 11162 6772
rect 11218 6716 11304 6772
rect 11360 6716 11430 6772
rect 11090 6630 11430 6716
rect 11090 6574 11162 6630
rect 11218 6574 11304 6630
rect 11360 6574 11430 6630
rect 11090 6488 11430 6574
rect 11090 6432 11162 6488
rect 11218 6432 11304 6488
rect 11360 6432 11430 6488
rect 11090 6346 11430 6432
rect 11090 6290 11162 6346
rect 11218 6290 11304 6346
rect 11360 6290 11430 6346
rect 11090 6204 11430 6290
rect 11090 6148 11162 6204
rect 11218 6148 11304 6204
rect 11360 6148 11430 6204
rect 11090 6062 11430 6148
rect 11090 6006 11162 6062
rect 11218 6006 11304 6062
rect 11360 6006 11430 6062
rect 11090 5920 11430 6006
rect 11090 5864 11162 5920
rect 11218 5864 11304 5920
rect 11360 5864 11430 5920
rect 11090 5778 11430 5864
rect 11090 5722 11162 5778
rect 11218 5722 11304 5778
rect 11360 5722 11430 5778
rect 11090 5636 11430 5722
rect 11090 5580 11162 5636
rect 11218 5580 11304 5636
rect 11360 5580 11430 5636
rect 11090 5494 11430 5580
rect 11090 5438 11162 5494
rect 11218 5438 11304 5494
rect 11360 5438 11430 5494
rect 11090 5352 11430 5438
rect 11090 5296 11162 5352
rect 11218 5296 11304 5352
rect 11360 5296 11430 5352
rect 11090 5210 11430 5296
rect 11090 5154 11162 5210
rect 11218 5154 11304 5210
rect 11360 5154 11430 5210
rect 11090 5068 11430 5154
rect 11090 5012 11162 5068
rect 11218 5012 11304 5068
rect 11360 5012 11430 5068
rect 11090 4926 11430 5012
rect 11090 4870 11162 4926
rect 11218 4870 11304 4926
rect 11360 4870 11430 4926
rect 11090 4784 11430 4870
rect 11090 4728 11162 4784
rect 11218 4728 11304 4784
rect 11360 4728 11430 4784
rect 11090 4642 11430 4728
rect 11090 4586 11162 4642
rect 11218 4586 11304 4642
rect 11360 4586 11430 4642
rect 11090 4500 11430 4586
rect 11090 4444 11162 4500
rect 11218 4444 11304 4500
rect 11360 4444 11430 4500
rect 11090 4358 11430 4444
rect 11090 4302 11162 4358
rect 11218 4302 11304 4358
rect 11360 4302 11430 4358
rect 11090 4216 11430 4302
rect 11090 4160 11162 4216
rect 11218 4160 11304 4216
rect 11360 4160 11430 4216
rect 11090 4074 11430 4160
rect 11090 4018 11162 4074
rect 11218 4018 11304 4074
rect 11360 4018 11430 4074
rect 11090 3932 11430 4018
rect 11090 3876 11162 3932
rect 11218 3876 11304 3932
rect 11360 3876 11430 3932
rect 11090 3790 11430 3876
rect 11090 3734 11162 3790
rect 11218 3734 11304 3790
rect 11360 3734 11430 3790
rect 11090 3648 11430 3734
rect 11090 3592 11162 3648
rect 11218 3592 11304 3648
rect 11360 3592 11430 3648
rect 11090 3506 11430 3592
rect 11090 3450 11162 3506
rect 11218 3450 11304 3506
rect 11360 3450 11430 3506
rect 11090 3364 11430 3450
rect 11090 3308 11162 3364
rect 11218 3308 11304 3364
rect 11360 3308 11430 3364
rect 11090 3222 11430 3308
rect 11090 3166 11162 3222
rect 11218 3166 11304 3222
rect 11360 3166 11430 3222
rect 11090 3080 11430 3166
rect 11090 3024 11162 3080
rect 11218 3024 11304 3080
rect 11360 3024 11430 3080
rect 11090 2938 11430 3024
rect 11090 2882 11162 2938
rect 11218 2882 11304 2938
rect 11360 2882 11430 2938
rect 11090 2796 11430 2882
rect 11090 2740 11162 2796
rect 11218 2740 11304 2796
rect 11360 2740 11430 2796
rect 11090 2654 11430 2740
rect 11090 2598 11162 2654
rect 11218 2598 11304 2654
rect 11360 2598 11430 2654
rect 11090 2512 11430 2598
rect 11090 2456 11162 2512
rect 11218 2456 11304 2512
rect 11360 2456 11430 2512
rect 11090 2370 11430 2456
rect 11090 2314 11162 2370
rect 11218 2314 11304 2370
rect 11360 2314 11430 2370
rect 11090 2228 11430 2314
rect 11090 2172 11162 2228
rect 11218 2172 11304 2228
rect 11360 2172 11430 2228
rect 11090 2086 11430 2172
rect 11090 2030 11162 2086
rect 11218 2030 11304 2086
rect 11360 2030 11430 2086
rect 11090 1944 11430 2030
rect 11090 1888 11162 1944
rect 11218 1888 11304 1944
rect 11360 1888 11430 1944
rect 11090 1802 11430 1888
rect 11090 1746 11162 1802
rect 11218 1746 11304 1802
rect 11360 1746 11430 1802
rect 11090 1660 11430 1746
rect 11090 1604 11162 1660
rect 11218 1604 11304 1660
rect 11360 1604 11430 1660
rect 11090 1518 11430 1604
rect 11090 1462 11162 1518
rect 11218 1462 11304 1518
rect 11360 1462 11430 1518
rect 11090 1376 11430 1462
rect 11090 1320 11162 1376
rect 11218 1320 11304 1376
rect 11360 1320 11430 1376
rect 11090 1234 11430 1320
rect 11090 1178 11162 1234
rect 11218 1178 11304 1234
rect 11360 1178 11430 1234
rect 11090 1092 11430 1178
rect 11090 1036 11162 1092
rect 11218 1036 11304 1092
rect 11360 1036 11430 1092
rect 11090 950 11430 1036
rect 11090 894 11162 950
rect 11218 894 11304 950
rect 11360 894 11430 950
rect 11090 808 11430 894
rect 11090 752 11162 808
rect 11218 752 11304 808
rect 11360 752 11430 808
rect 11090 666 11430 752
rect 11090 610 11162 666
rect 11218 610 11304 666
rect 11360 610 11430 666
rect 11090 524 11430 610
rect 11090 468 11162 524
rect 11218 468 11304 524
rect 11360 468 11430 524
rect 11090 458 11430 468
rect 11630 12310 11970 12320
rect 11630 12254 11702 12310
rect 11758 12254 11844 12310
rect 11900 12254 11970 12310
rect 11630 12168 11970 12254
rect 11630 12112 11702 12168
rect 11758 12112 11844 12168
rect 11900 12112 11970 12168
rect 11630 12026 11970 12112
rect 11630 11970 11702 12026
rect 11758 11970 11844 12026
rect 11900 11970 11970 12026
rect 11630 11884 11970 11970
rect 11630 11828 11702 11884
rect 11758 11828 11844 11884
rect 11900 11828 11970 11884
rect 11630 11742 11970 11828
rect 11630 11686 11702 11742
rect 11758 11686 11844 11742
rect 11900 11686 11970 11742
rect 11630 11600 11970 11686
rect 11630 11544 11702 11600
rect 11758 11544 11844 11600
rect 11900 11544 11970 11600
rect 11630 11458 11970 11544
rect 11630 11402 11702 11458
rect 11758 11402 11844 11458
rect 11900 11402 11970 11458
rect 11630 11316 11970 11402
rect 11630 11260 11702 11316
rect 11758 11260 11844 11316
rect 11900 11260 11970 11316
rect 11630 11174 11970 11260
rect 11630 11118 11702 11174
rect 11758 11118 11844 11174
rect 11900 11118 11970 11174
rect 11630 11032 11970 11118
rect 11630 10976 11702 11032
rect 11758 10976 11844 11032
rect 11900 10976 11970 11032
rect 11630 10890 11970 10976
rect 11630 10834 11702 10890
rect 11758 10834 11844 10890
rect 11900 10834 11970 10890
rect 11630 10748 11970 10834
rect 11630 10692 11702 10748
rect 11758 10692 11844 10748
rect 11900 10692 11970 10748
rect 11630 10606 11970 10692
rect 11630 10550 11702 10606
rect 11758 10550 11844 10606
rect 11900 10550 11970 10606
rect 11630 10464 11970 10550
rect 11630 10408 11702 10464
rect 11758 10408 11844 10464
rect 11900 10408 11970 10464
rect 11630 10322 11970 10408
rect 11630 10266 11702 10322
rect 11758 10266 11844 10322
rect 11900 10266 11970 10322
rect 11630 10180 11970 10266
rect 11630 10124 11702 10180
rect 11758 10124 11844 10180
rect 11900 10124 11970 10180
rect 11630 10038 11970 10124
rect 11630 9982 11702 10038
rect 11758 9982 11844 10038
rect 11900 9982 11970 10038
rect 11630 9896 11970 9982
rect 11630 9840 11702 9896
rect 11758 9840 11844 9896
rect 11900 9840 11970 9896
rect 11630 9754 11970 9840
rect 11630 9698 11702 9754
rect 11758 9698 11844 9754
rect 11900 9698 11970 9754
rect 11630 9612 11970 9698
rect 11630 9556 11702 9612
rect 11758 9556 11844 9612
rect 11900 9556 11970 9612
rect 11630 9470 11970 9556
rect 11630 9414 11702 9470
rect 11758 9414 11844 9470
rect 11900 9414 11970 9470
rect 11630 9328 11970 9414
rect 11630 9272 11702 9328
rect 11758 9272 11844 9328
rect 11900 9272 11970 9328
rect 11630 9186 11970 9272
rect 11630 9130 11702 9186
rect 11758 9130 11844 9186
rect 11900 9130 11970 9186
rect 11630 9044 11970 9130
rect 11630 8988 11702 9044
rect 11758 8988 11844 9044
rect 11900 8988 11970 9044
rect 11630 8902 11970 8988
rect 11630 8846 11702 8902
rect 11758 8846 11844 8902
rect 11900 8846 11970 8902
rect 11630 8760 11970 8846
rect 11630 8704 11702 8760
rect 11758 8704 11844 8760
rect 11900 8704 11970 8760
rect 11630 8618 11970 8704
rect 11630 8562 11702 8618
rect 11758 8562 11844 8618
rect 11900 8562 11970 8618
rect 11630 8476 11970 8562
rect 11630 8420 11702 8476
rect 11758 8420 11844 8476
rect 11900 8420 11970 8476
rect 11630 8334 11970 8420
rect 11630 8278 11702 8334
rect 11758 8278 11844 8334
rect 11900 8278 11970 8334
rect 11630 8192 11970 8278
rect 11630 8136 11702 8192
rect 11758 8136 11844 8192
rect 11900 8136 11970 8192
rect 11630 8050 11970 8136
rect 11630 7994 11702 8050
rect 11758 7994 11844 8050
rect 11900 7994 11970 8050
rect 11630 7908 11970 7994
rect 11630 7852 11702 7908
rect 11758 7852 11844 7908
rect 11900 7852 11970 7908
rect 11630 7766 11970 7852
rect 11630 7710 11702 7766
rect 11758 7710 11844 7766
rect 11900 7710 11970 7766
rect 11630 7624 11970 7710
rect 11630 7568 11702 7624
rect 11758 7568 11844 7624
rect 11900 7568 11970 7624
rect 11630 7482 11970 7568
rect 11630 7426 11702 7482
rect 11758 7426 11844 7482
rect 11900 7426 11970 7482
rect 11630 7340 11970 7426
rect 11630 7284 11702 7340
rect 11758 7284 11844 7340
rect 11900 7284 11970 7340
rect 11630 7198 11970 7284
rect 11630 7142 11702 7198
rect 11758 7142 11844 7198
rect 11900 7142 11970 7198
rect 11630 7056 11970 7142
rect 11630 7000 11702 7056
rect 11758 7000 11844 7056
rect 11900 7000 11970 7056
rect 11630 6914 11970 7000
rect 11630 6858 11702 6914
rect 11758 6858 11844 6914
rect 11900 6858 11970 6914
rect 11630 6772 11970 6858
rect 11630 6716 11702 6772
rect 11758 6716 11844 6772
rect 11900 6716 11970 6772
rect 11630 6630 11970 6716
rect 11630 6574 11702 6630
rect 11758 6574 11844 6630
rect 11900 6574 11970 6630
rect 11630 6488 11970 6574
rect 11630 6432 11702 6488
rect 11758 6432 11844 6488
rect 11900 6432 11970 6488
rect 11630 6346 11970 6432
rect 11630 6290 11702 6346
rect 11758 6290 11844 6346
rect 11900 6290 11970 6346
rect 11630 6204 11970 6290
rect 11630 6148 11702 6204
rect 11758 6148 11844 6204
rect 11900 6148 11970 6204
rect 11630 6062 11970 6148
rect 11630 6006 11702 6062
rect 11758 6006 11844 6062
rect 11900 6006 11970 6062
rect 11630 5920 11970 6006
rect 11630 5864 11702 5920
rect 11758 5864 11844 5920
rect 11900 5864 11970 5920
rect 11630 5778 11970 5864
rect 11630 5722 11702 5778
rect 11758 5722 11844 5778
rect 11900 5722 11970 5778
rect 11630 5636 11970 5722
rect 11630 5580 11702 5636
rect 11758 5580 11844 5636
rect 11900 5580 11970 5636
rect 11630 5494 11970 5580
rect 11630 5438 11702 5494
rect 11758 5438 11844 5494
rect 11900 5438 11970 5494
rect 11630 5352 11970 5438
rect 11630 5296 11702 5352
rect 11758 5296 11844 5352
rect 11900 5296 11970 5352
rect 11630 5210 11970 5296
rect 11630 5154 11702 5210
rect 11758 5154 11844 5210
rect 11900 5154 11970 5210
rect 11630 5068 11970 5154
rect 11630 5012 11702 5068
rect 11758 5012 11844 5068
rect 11900 5012 11970 5068
rect 11630 4926 11970 5012
rect 11630 4870 11702 4926
rect 11758 4870 11844 4926
rect 11900 4870 11970 4926
rect 11630 4784 11970 4870
rect 11630 4728 11702 4784
rect 11758 4728 11844 4784
rect 11900 4728 11970 4784
rect 11630 4642 11970 4728
rect 11630 4586 11702 4642
rect 11758 4586 11844 4642
rect 11900 4586 11970 4642
rect 11630 4500 11970 4586
rect 11630 4444 11702 4500
rect 11758 4444 11844 4500
rect 11900 4444 11970 4500
rect 11630 4358 11970 4444
rect 11630 4302 11702 4358
rect 11758 4302 11844 4358
rect 11900 4302 11970 4358
rect 11630 4216 11970 4302
rect 11630 4160 11702 4216
rect 11758 4160 11844 4216
rect 11900 4160 11970 4216
rect 11630 4074 11970 4160
rect 11630 4018 11702 4074
rect 11758 4018 11844 4074
rect 11900 4018 11970 4074
rect 11630 3932 11970 4018
rect 11630 3876 11702 3932
rect 11758 3876 11844 3932
rect 11900 3876 11970 3932
rect 11630 3790 11970 3876
rect 11630 3734 11702 3790
rect 11758 3734 11844 3790
rect 11900 3734 11970 3790
rect 11630 3648 11970 3734
rect 11630 3592 11702 3648
rect 11758 3592 11844 3648
rect 11900 3592 11970 3648
rect 11630 3506 11970 3592
rect 11630 3450 11702 3506
rect 11758 3450 11844 3506
rect 11900 3450 11970 3506
rect 11630 3364 11970 3450
rect 11630 3308 11702 3364
rect 11758 3308 11844 3364
rect 11900 3308 11970 3364
rect 11630 3222 11970 3308
rect 11630 3166 11702 3222
rect 11758 3166 11844 3222
rect 11900 3166 11970 3222
rect 11630 3080 11970 3166
rect 11630 3024 11702 3080
rect 11758 3024 11844 3080
rect 11900 3024 11970 3080
rect 11630 2938 11970 3024
rect 11630 2882 11702 2938
rect 11758 2882 11844 2938
rect 11900 2882 11970 2938
rect 11630 2796 11970 2882
rect 11630 2740 11702 2796
rect 11758 2740 11844 2796
rect 11900 2740 11970 2796
rect 11630 2654 11970 2740
rect 11630 2598 11702 2654
rect 11758 2598 11844 2654
rect 11900 2598 11970 2654
rect 11630 2512 11970 2598
rect 11630 2456 11702 2512
rect 11758 2456 11844 2512
rect 11900 2456 11970 2512
rect 11630 2370 11970 2456
rect 11630 2314 11702 2370
rect 11758 2314 11844 2370
rect 11900 2314 11970 2370
rect 11630 2228 11970 2314
rect 11630 2172 11702 2228
rect 11758 2172 11844 2228
rect 11900 2172 11970 2228
rect 11630 2086 11970 2172
rect 11630 2030 11702 2086
rect 11758 2030 11844 2086
rect 11900 2030 11970 2086
rect 11630 1944 11970 2030
rect 11630 1888 11702 1944
rect 11758 1888 11844 1944
rect 11900 1888 11970 1944
rect 11630 1802 11970 1888
rect 11630 1746 11702 1802
rect 11758 1746 11844 1802
rect 11900 1746 11970 1802
rect 11630 1660 11970 1746
rect 11630 1604 11702 1660
rect 11758 1604 11844 1660
rect 11900 1604 11970 1660
rect 11630 1518 11970 1604
rect 11630 1462 11702 1518
rect 11758 1462 11844 1518
rect 11900 1462 11970 1518
rect 11630 1376 11970 1462
rect 11630 1320 11702 1376
rect 11758 1320 11844 1376
rect 11900 1320 11970 1376
rect 11630 1234 11970 1320
rect 11630 1178 11702 1234
rect 11758 1178 11844 1234
rect 11900 1178 11970 1234
rect 11630 1092 11970 1178
rect 11630 1036 11702 1092
rect 11758 1036 11844 1092
rect 11900 1036 11970 1092
rect 11630 950 11970 1036
rect 11630 894 11702 950
rect 11758 894 11844 950
rect 11900 894 11970 950
rect 11630 808 11970 894
rect 11630 752 11702 808
rect 11758 752 11844 808
rect 11900 752 11970 808
rect 11630 666 11970 752
rect 11630 610 11702 666
rect 11758 610 11844 666
rect 11900 610 11970 666
rect 11630 524 11970 610
rect 11630 468 11702 524
rect 11758 468 11844 524
rect 11900 468 11970 524
rect 11630 458 11970 468
rect 12400 12302 12526 12320
rect 12582 12302 12650 12358
rect 12706 12302 12774 12358
rect 12830 12302 12898 12358
rect 12954 12302 13022 12358
rect 13078 12302 13200 12358
rect 12400 12234 13200 12302
rect 12400 12178 12526 12234
rect 12582 12178 12650 12234
rect 12706 12178 12774 12234
rect 12830 12178 12898 12234
rect 12954 12178 13022 12234
rect 13078 12178 13200 12234
rect 12400 12110 13200 12178
rect 12400 12054 12526 12110
rect 12582 12054 12650 12110
rect 12706 12054 12774 12110
rect 12830 12054 12898 12110
rect 12954 12054 13022 12110
rect 13078 12054 13200 12110
rect 12400 11986 13200 12054
rect 12400 11930 12526 11986
rect 12582 11930 12650 11986
rect 12706 11930 12774 11986
rect 12830 11930 12898 11986
rect 12954 11930 13022 11986
rect 13078 11930 13200 11986
rect 12400 11862 13200 11930
rect 12400 11806 12526 11862
rect 12582 11806 12650 11862
rect 12706 11806 12774 11862
rect 12830 11806 12898 11862
rect 12954 11806 13022 11862
rect 13078 11806 13200 11862
rect 12400 11738 13200 11806
rect 12400 11682 12526 11738
rect 12582 11682 12650 11738
rect 12706 11682 12774 11738
rect 12830 11682 12898 11738
rect 12954 11682 13022 11738
rect 13078 11682 13200 11738
rect 12400 11614 13200 11682
rect 12400 11558 12526 11614
rect 12582 11558 12650 11614
rect 12706 11558 12774 11614
rect 12830 11558 12898 11614
rect 12954 11558 13022 11614
rect 13078 11558 13200 11614
rect 12400 11490 13200 11558
rect 12400 11434 12526 11490
rect 12582 11434 12650 11490
rect 12706 11434 12774 11490
rect 12830 11434 12898 11490
rect 12954 11434 13022 11490
rect 13078 11434 13200 11490
rect 12400 11366 13200 11434
rect 12400 11310 12526 11366
rect 12582 11310 12650 11366
rect 12706 11310 12774 11366
rect 12830 11310 12898 11366
rect 12954 11310 13022 11366
rect 13078 11310 13200 11366
rect 12400 11242 13200 11310
rect 12400 11186 12526 11242
rect 12582 11186 12650 11242
rect 12706 11186 12774 11242
rect 12830 11186 12898 11242
rect 12954 11186 13022 11242
rect 13078 11186 13200 11242
rect 12400 11118 13200 11186
rect 12400 11062 12526 11118
rect 12582 11062 12650 11118
rect 12706 11062 12774 11118
rect 12830 11062 12898 11118
rect 12954 11062 13022 11118
rect 13078 11062 13200 11118
rect 12400 10994 13200 11062
rect 12400 10938 12526 10994
rect 12582 10938 12650 10994
rect 12706 10938 12774 10994
rect 12830 10938 12898 10994
rect 12954 10938 13022 10994
rect 13078 10938 13200 10994
rect 12400 10870 13200 10938
rect 12400 10814 12526 10870
rect 12582 10814 12650 10870
rect 12706 10814 12774 10870
rect 12830 10814 12898 10870
rect 12954 10814 13022 10870
rect 13078 10814 13200 10870
rect 12400 10746 13200 10814
rect 12400 10690 12526 10746
rect 12582 10690 12650 10746
rect 12706 10690 12774 10746
rect 12830 10690 12898 10746
rect 12954 10690 13022 10746
rect 13078 10690 13200 10746
rect 12400 10622 13200 10690
rect 12400 10566 12526 10622
rect 12582 10566 12650 10622
rect 12706 10566 12774 10622
rect 12830 10566 12898 10622
rect 12954 10566 13022 10622
rect 13078 10566 13200 10622
rect 12400 10498 13200 10566
rect 12400 10442 12526 10498
rect 12582 10442 12650 10498
rect 12706 10442 12774 10498
rect 12830 10442 12898 10498
rect 12954 10442 13022 10498
rect 13078 10442 13200 10498
rect 12400 10374 13200 10442
rect 12400 10318 12526 10374
rect 12582 10318 12650 10374
rect 12706 10318 12774 10374
rect 12830 10318 12898 10374
rect 12954 10318 13022 10374
rect 13078 10318 13200 10374
rect 12400 10250 13200 10318
rect 12400 10194 12526 10250
rect 12582 10194 12650 10250
rect 12706 10194 12774 10250
rect 12830 10194 12898 10250
rect 12954 10194 13022 10250
rect 13078 10194 13200 10250
rect 12400 10126 13200 10194
rect 12400 10070 12526 10126
rect 12582 10070 12650 10126
rect 12706 10070 12774 10126
rect 12830 10070 12898 10126
rect 12954 10070 13022 10126
rect 13078 10070 13200 10126
rect 12400 10002 13200 10070
rect 12400 9946 12526 10002
rect 12582 9946 12650 10002
rect 12706 9946 12774 10002
rect 12830 9946 12898 10002
rect 12954 9946 13022 10002
rect 13078 9946 13200 10002
rect 12400 9878 13200 9946
rect 12400 9822 12526 9878
rect 12582 9822 12650 9878
rect 12706 9822 12774 9878
rect 12830 9822 12898 9878
rect 12954 9822 13022 9878
rect 13078 9822 13200 9878
rect 12400 9754 13200 9822
rect 12400 9698 12526 9754
rect 12582 9698 12650 9754
rect 12706 9698 12774 9754
rect 12830 9698 12898 9754
rect 12954 9698 13022 9754
rect 13078 9698 13200 9754
rect 12400 9630 13200 9698
rect 12400 9574 12526 9630
rect 12582 9574 12650 9630
rect 12706 9574 12774 9630
rect 12830 9574 12898 9630
rect 12954 9574 13022 9630
rect 13078 9574 13200 9630
rect 12400 9506 13200 9574
rect 12400 9450 12526 9506
rect 12582 9450 12650 9506
rect 12706 9450 12774 9506
rect 12830 9450 12898 9506
rect 12954 9450 13022 9506
rect 13078 9450 13200 9506
rect 12400 9382 13200 9450
rect 12400 9326 12526 9382
rect 12582 9326 12650 9382
rect 12706 9326 12774 9382
rect 12830 9326 12898 9382
rect 12954 9326 13022 9382
rect 13078 9326 13200 9382
rect 12400 9258 13200 9326
rect 12400 9202 12526 9258
rect 12582 9202 12650 9258
rect 12706 9202 12774 9258
rect 12830 9202 12898 9258
rect 12954 9202 13022 9258
rect 13078 9202 13200 9258
rect 12400 9134 13200 9202
rect 12400 9078 12526 9134
rect 12582 9078 12650 9134
rect 12706 9078 12774 9134
rect 12830 9078 12898 9134
rect 12954 9078 13022 9134
rect 13078 9078 13200 9134
rect 12400 9010 13200 9078
rect 12400 8954 12526 9010
rect 12582 8954 12650 9010
rect 12706 8954 12774 9010
rect 12830 8954 12898 9010
rect 12954 8954 13022 9010
rect 13078 8954 13200 9010
rect 12400 8886 13200 8954
rect 12400 8830 12526 8886
rect 12582 8830 12650 8886
rect 12706 8830 12774 8886
rect 12830 8830 12898 8886
rect 12954 8830 13022 8886
rect 13078 8830 13200 8886
rect 12400 8762 13200 8830
rect 12400 8706 12526 8762
rect 12582 8706 12650 8762
rect 12706 8706 12774 8762
rect 12830 8706 12898 8762
rect 12954 8706 13022 8762
rect 13078 8706 13200 8762
rect 12400 8638 13200 8706
rect 12400 8582 12526 8638
rect 12582 8582 12650 8638
rect 12706 8582 12774 8638
rect 12830 8582 12898 8638
rect 12954 8582 13022 8638
rect 13078 8582 13200 8638
rect 12400 8514 13200 8582
rect 12400 8458 12526 8514
rect 12582 8458 12650 8514
rect 12706 8458 12774 8514
rect 12830 8458 12898 8514
rect 12954 8458 13022 8514
rect 13078 8458 13200 8514
rect 12400 8390 13200 8458
rect 12400 8334 12526 8390
rect 12582 8334 12650 8390
rect 12706 8334 12774 8390
rect 12830 8334 12898 8390
rect 12954 8334 13022 8390
rect 13078 8334 13200 8390
rect 12400 8266 13200 8334
rect 12400 8210 12526 8266
rect 12582 8210 12650 8266
rect 12706 8210 12774 8266
rect 12830 8210 12898 8266
rect 12954 8210 13022 8266
rect 13078 8210 13200 8266
rect 12400 8142 13200 8210
rect 12400 8086 12526 8142
rect 12582 8086 12650 8142
rect 12706 8086 12774 8142
rect 12830 8086 12898 8142
rect 12954 8086 13022 8142
rect 13078 8086 13200 8142
rect 12400 8018 13200 8086
rect 12400 7962 12526 8018
rect 12582 7962 12650 8018
rect 12706 7962 12774 8018
rect 12830 7962 12898 8018
rect 12954 7962 13022 8018
rect 13078 7962 13200 8018
rect 12400 7894 13200 7962
rect 12400 7838 12526 7894
rect 12582 7838 12650 7894
rect 12706 7838 12774 7894
rect 12830 7838 12898 7894
rect 12954 7838 13022 7894
rect 13078 7838 13200 7894
rect 12400 7770 13200 7838
rect 12400 7714 12526 7770
rect 12582 7714 12650 7770
rect 12706 7714 12774 7770
rect 12830 7714 12898 7770
rect 12954 7714 13022 7770
rect 13078 7714 13200 7770
rect 12400 7646 13200 7714
rect 12400 7590 12526 7646
rect 12582 7590 12650 7646
rect 12706 7590 12774 7646
rect 12830 7590 12898 7646
rect 12954 7590 13022 7646
rect 13078 7590 13200 7646
rect 12400 7522 13200 7590
rect 12400 7466 12526 7522
rect 12582 7466 12650 7522
rect 12706 7466 12774 7522
rect 12830 7466 12898 7522
rect 12954 7466 13022 7522
rect 13078 7466 13200 7522
rect 12400 7398 13200 7466
rect 12400 7342 12526 7398
rect 12582 7342 12650 7398
rect 12706 7342 12774 7398
rect 12830 7342 12898 7398
rect 12954 7342 13022 7398
rect 13078 7342 13200 7398
rect 12400 7274 13200 7342
rect 12400 7218 12526 7274
rect 12582 7218 12650 7274
rect 12706 7218 12774 7274
rect 12830 7218 12898 7274
rect 12954 7218 13022 7274
rect 13078 7218 13200 7274
rect 12400 7150 13200 7218
rect 12400 7094 12526 7150
rect 12582 7094 12650 7150
rect 12706 7094 12774 7150
rect 12830 7094 12898 7150
rect 12954 7094 13022 7150
rect 13078 7094 13200 7150
rect 12400 7026 13200 7094
rect 12400 6970 12526 7026
rect 12582 6970 12650 7026
rect 12706 6970 12774 7026
rect 12830 6970 12898 7026
rect 12954 6970 13022 7026
rect 13078 6970 13200 7026
rect 12400 6902 13200 6970
rect 12400 6846 12526 6902
rect 12582 6846 12650 6902
rect 12706 6846 12774 6902
rect 12830 6846 12898 6902
rect 12954 6846 13022 6902
rect 13078 6846 13200 6902
rect 12400 6778 13200 6846
rect 12400 6722 12526 6778
rect 12582 6722 12650 6778
rect 12706 6722 12774 6778
rect 12830 6722 12898 6778
rect 12954 6722 13022 6778
rect 13078 6722 13200 6778
rect 12400 6654 13200 6722
rect 12400 6598 12526 6654
rect 12582 6598 12650 6654
rect 12706 6598 12774 6654
rect 12830 6598 12898 6654
rect 12954 6598 13022 6654
rect 13078 6598 13200 6654
rect 12400 6530 13200 6598
rect 12400 6474 12526 6530
rect 12582 6474 12650 6530
rect 12706 6474 12774 6530
rect 12830 6474 12898 6530
rect 12954 6474 13022 6530
rect 13078 6474 13200 6530
rect 12400 6406 13200 6474
rect 12400 6350 12526 6406
rect 12582 6350 12650 6406
rect 12706 6350 12774 6406
rect 12830 6350 12898 6406
rect 12954 6350 13022 6406
rect 13078 6350 13200 6406
rect 12400 6282 13200 6350
rect 12400 6226 12526 6282
rect 12582 6226 12650 6282
rect 12706 6226 12774 6282
rect 12830 6226 12898 6282
rect 12954 6226 13022 6282
rect 13078 6226 13200 6282
rect 12400 6158 13200 6226
rect 12400 6102 12526 6158
rect 12582 6102 12650 6158
rect 12706 6102 12774 6158
rect 12830 6102 12898 6158
rect 12954 6102 13022 6158
rect 13078 6102 13200 6158
rect 12400 6034 13200 6102
rect 12400 5978 12526 6034
rect 12582 5978 12650 6034
rect 12706 5978 12774 6034
rect 12830 5978 12898 6034
rect 12954 5978 13022 6034
rect 13078 5978 13200 6034
rect 12400 5910 13200 5978
rect 12400 5854 12526 5910
rect 12582 5854 12650 5910
rect 12706 5854 12774 5910
rect 12830 5854 12898 5910
rect 12954 5854 13022 5910
rect 13078 5854 13200 5910
rect 12400 5786 13200 5854
rect 12400 5730 12526 5786
rect 12582 5730 12650 5786
rect 12706 5730 12774 5786
rect 12830 5730 12898 5786
rect 12954 5730 13022 5786
rect 13078 5730 13200 5786
rect 12400 5662 13200 5730
rect 12400 5606 12526 5662
rect 12582 5606 12650 5662
rect 12706 5606 12774 5662
rect 12830 5606 12898 5662
rect 12954 5606 13022 5662
rect 13078 5606 13200 5662
rect 12400 5538 13200 5606
rect 12400 5482 12526 5538
rect 12582 5482 12650 5538
rect 12706 5482 12774 5538
rect 12830 5482 12898 5538
rect 12954 5482 13022 5538
rect 13078 5482 13200 5538
rect 12400 5414 13200 5482
rect 12400 5358 12526 5414
rect 12582 5358 12650 5414
rect 12706 5358 12774 5414
rect 12830 5358 12898 5414
rect 12954 5358 13022 5414
rect 13078 5358 13200 5414
rect 12400 5290 13200 5358
rect 12400 5234 12526 5290
rect 12582 5234 12650 5290
rect 12706 5234 12774 5290
rect 12830 5234 12898 5290
rect 12954 5234 13022 5290
rect 13078 5234 13200 5290
rect 12400 5166 13200 5234
rect 12400 5110 12526 5166
rect 12582 5110 12650 5166
rect 12706 5110 12774 5166
rect 12830 5110 12898 5166
rect 12954 5110 13022 5166
rect 13078 5110 13200 5166
rect 12400 5042 13200 5110
rect 12400 4986 12526 5042
rect 12582 4986 12650 5042
rect 12706 4986 12774 5042
rect 12830 4986 12898 5042
rect 12954 4986 13022 5042
rect 13078 4986 13200 5042
rect 12400 4918 13200 4986
rect 12400 4862 12526 4918
rect 12582 4862 12650 4918
rect 12706 4862 12774 4918
rect 12830 4862 12898 4918
rect 12954 4862 13022 4918
rect 13078 4862 13200 4918
rect 12400 4794 13200 4862
rect 12400 4738 12526 4794
rect 12582 4738 12650 4794
rect 12706 4738 12774 4794
rect 12830 4738 12898 4794
rect 12954 4738 13022 4794
rect 13078 4738 13200 4794
rect 12400 4670 13200 4738
rect 12400 4614 12526 4670
rect 12582 4614 12650 4670
rect 12706 4614 12774 4670
rect 12830 4614 12898 4670
rect 12954 4614 13022 4670
rect 13078 4614 13200 4670
rect 12400 4546 13200 4614
rect 12400 4490 12526 4546
rect 12582 4490 12650 4546
rect 12706 4490 12774 4546
rect 12830 4490 12898 4546
rect 12954 4490 13022 4546
rect 13078 4490 13200 4546
rect 12400 4422 13200 4490
rect 12400 4366 12526 4422
rect 12582 4366 12650 4422
rect 12706 4366 12774 4422
rect 12830 4366 12898 4422
rect 12954 4366 13022 4422
rect 13078 4366 13200 4422
rect 12400 4298 13200 4366
rect 12400 4242 12526 4298
rect 12582 4242 12650 4298
rect 12706 4242 12774 4298
rect 12830 4242 12898 4298
rect 12954 4242 13022 4298
rect 13078 4242 13200 4298
rect 12400 4174 13200 4242
rect 12400 4118 12526 4174
rect 12582 4118 12650 4174
rect 12706 4118 12774 4174
rect 12830 4118 12898 4174
rect 12954 4118 13022 4174
rect 13078 4118 13200 4174
rect 12400 4050 13200 4118
rect 12400 3994 12526 4050
rect 12582 3994 12650 4050
rect 12706 3994 12774 4050
rect 12830 3994 12898 4050
rect 12954 3994 13022 4050
rect 13078 3994 13200 4050
rect 12400 3926 13200 3994
rect 12400 3870 12526 3926
rect 12582 3870 12650 3926
rect 12706 3870 12774 3926
rect 12830 3870 12898 3926
rect 12954 3870 13022 3926
rect 13078 3870 13200 3926
rect 12400 3802 13200 3870
rect 12400 3746 12526 3802
rect 12582 3746 12650 3802
rect 12706 3746 12774 3802
rect 12830 3746 12898 3802
rect 12954 3746 13022 3802
rect 13078 3746 13200 3802
rect 12400 3678 13200 3746
rect 12400 3622 12526 3678
rect 12582 3622 12650 3678
rect 12706 3622 12774 3678
rect 12830 3622 12898 3678
rect 12954 3622 13022 3678
rect 13078 3622 13200 3678
rect 12400 3554 13200 3622
rect 12400 3498 12526 3554
rect 12582 3498 12650 3554
rect 12706 3498 12774 3554
rect 12830 3498 12898 3554
rect 12954 3498 13022 3554
rect 13078 3498 13200 3554
rect 12400 3430 13200 3498
rect 12400 3374 12526 3430
rect 12582 3374 12650 3430
rect 12706 3374 12774 3430
rect 12830 3374 12898 3430
rect 12954 3374 13022 3430
rect 13078 3374 13200 3430
rect 12400 3306 13200 3374
rect 12400 3250 12526 3306
rect 12582 3250 12650 3306
rect 12706 3250 12774 3306
rect 12830 3250 12898 3306
rect 12954 3250 13022 3306
rect 13078 3250 13200 3306
rect 12400 3182 13200 3250
rect 12400 3126 12526 3182
rect 12582 3126 12650 3182
rect 12706 3126 12774 3182
rect 12830 3126 12898 3182
rect 12954 3126 13022 3182
rect 13078 3126 13200 3182
rect 12400 3058 13200 3126
rect 12400 3002 12526 3058
rect 12582 3002 12650 3058
rect 12706 3002 12774 3058
rect 12830 3002 12898 3058
rect 12954 3002 13022 3058
rect 13078 3002 13200 3058
rect 12400 2934 13200 3002
rect 12400 2878 12526 2934
rect 12582 2878 12650 2934
rect 12706 2878 12774 2934
rect 12830 2878 12898 2934
rect 12954 2878 13022 2934
rect 13078 2878 13200 2934
rect 12400 2810 13200 2878
rect 12400 2754 12526 2810
rect 12582 2754 12650 2810
rect 12706 2754 12774 2810
rect 12830 2754 12898 2810
rect 12954 2754 13022 2810
rect 13078 2754 13200 2810
rect 12400 2686 13200 2754
rect 12400 2630 12526 2686
rect 12582 2630 12650 2686
rect 12706 2630 12774 2686
rect 12830 2630 12898 2686
rect 12954 2630 13022 2686
rect 13078 2630 13200 2686
rect 12400 2562 13200 2630
rect 12400 2506 12526 2562
rect 12582 2506 12650 2562
rect 12706 2506 12774 2562
rect 12830 2506 12898 2562
rect 12954 2506 13022 2562
rect 13078 2506 13200 2562
rect 12400 2438 13200 2506
rect 12400 2382 12526 2438
rect 12582 2382 12650 2438
rect 12706 2382 12774 2438
rect 12830 2382 12898 2438
rect 12954 2382 13022 2438
rect 13078 2382 13200 2438
rect 12400 2314 13200 2382
rect 12400 2258 12526 2314
rect 12582 2258 12650 2314
rect 12706 2258 12774 2314
rect 12830 2258 12898 2314
rect 12954 2258 13022 2314
rect 13078 2258 13200 2314
rect 12400 2190 13200 2258
rect 12400 2134 12526 2190
rect 12582 2134 12650 2190
rect 12706 2134 12774 2190
rect 12830 2134 12898 2190
rect 12954 2134 13022 2190
rect 13078 2134 13200 2190
rect 12400 2066 13200 2134
rect 12400 2010 12526 2066
rect 12582 2010 12650 2066
rect 12706 2010 12774 2066
rect 12830 2010 12898 2066
rect 12954 2010 13022 2066
rect 13078 2010 13200 2066
rect 12400 1942 13200 2010
rect 12400 1886 12526 1942
rect 12582 1886 12650 1942
rect 12706 1886 12774 1942
rect 12830 1886 12898 1942
rect 12954 1886 13022 1942
rect 13078 1886 13200 1942
rect 12400 1818 13200 1886
rect 12400 1762 12526 1818
rect 12582 1762 12650 1818
rect 12706 1762 12774 1818
rect 12830 1762 12898 1818
rect 12954 1762 13022 1818
rect 13078 1762 13200 1818
rect 12400 1694 13200 1762
rect 12400 1638 12526 1694
rect 12582 1638 12650 1694
rect 12706 1638 12774 1694
rect 12830 1638 12898 1694
rect 12954 1638 13022 1694
rect 13078 1638 13200 1694
rect 12400 1570 13200 1638
rect 12400 1514 12526 1570
rect 12582 1514 12650 1570
rect 12706 1514 12774 1570
rect 12830 1514 12898 1570
rect 12954 1514 13022 1570
rect 13078 1514 13200 1570
rect 12400 1446 13200 1514
rect 12400 1390 12526 1446
rect 12582 1390 12650 1446
rect 12706 1390 12774 1446
rect 12830 1390 12898 1446
rect 12954 1390 13022 1446
rect 13078 1390 13200 1446
rect 12400 1322 13200 1390
rect 12400 1266 12526 1322
rect 12582 1266 12650 1322
rect 12706 1266 12774 1322
rect 12830 1266 12898 1322
rect 12954 1266 13022 1322
rect 13078 1266 13200 1322
rect 12400 1198 13200 1266
rect 12400 1142 12526 1198
rect 12582 1142 12650 1198
rect 12706 1142 12774 1198
rect 12830 1142 12898 1198
rect 12954 1142 13022 1198
rect 13078 1142 13200 1198
rect 12400 1074 13200 1142
rect 12400 1018 12526 1074
rect 12582 1018 12650 1074
rect 12706 1018 12774 1074
rect 12830 1018 12898 1074
rect 12954 1018 13022 1074
rect 13078 1018 13200 1074
rect 12400 950 13200 1018
rect 12400 894 12526 950
rect 12582 894 12650 950
rect 12706 894 12774 950
rect 12830 894 12898 950
rect 12954 894 13022 950
rect 13078 894 13200 950
rect 12400 826 13200 894
rect 12400 770 12526 826
rect 12582 770 12650 826
rect 12706 770 12774 826
rect 12830 770 12898 826
rect 12954 770 13022 826
rect 13078 770 13200 826
rect 12400 702 13200 770
rect 12400 646 12526 702
rect 12582 646 12650 702
rect 12706 646 12774 702
rect 12830 646 12898 702
rect 12954 646 13022 702
rect 13078 646 13200 702
rect 12400 578 13200 646
rect 12400 522 12526 578
rect 12582 522 12650 578
rect 12706 522 12774 578
rect 12830 522 12898 578
rect 12954 522 13022 578
rect 13078 522 13200 578
rect 12400 458 13200 522
rect -400 454 13200 458
rect -400 398 -286 454
rect -230 398 -162 454
rect -106 398 -38 454
rect 18 398 86 454
rect 142 398 210 454
rect 266 398 12526 454
rect 12582 398 12650 454
rect 12706 398 12774 454
rect 12830 398 12898 454
rect 12954 398 13022 454
rect 13078 398 13200 454
rect -400 330 13200 398
rect -400 274 -286 330
rect -230 274 -162 330
rect -106 274 -38 330
rect 18 274 86 330
rect 142 274 210 330
rect 266 302 12526 330
rect 266 274 415 302
rect -400 246 415 274
rect 471 246 557 302
rect 613 246 699 302
rect 755 246 841 302
rect 897 246 983 302
rect 1039 246 1125 302
rect 1181 246 1267 302
rect 1323 246 1409 302
rect 1465 246 1551 302
rect 1607 246 1693 302
rect 1749 246 1835 302
rect 1891 246 1977 302
rect 2033 246 2119 302
rect 2175 246 2261 302
rect 2317 246 2403 302
rect 2459 246 2545 302
rect 2601 246 2687 302
rect 2743 246 2829 302
rect 2885 246 2971 302
rect 3027 246 3113 302
rect 3169 246 3255 302
rect 3311 246 3397 302
rect 3453 246 3539 302
rect 3595 246 3681 302
rect 3737 246 3823 302
rect 3879 246 3965 302
rect 4021 246 4107 302
rect 4163 246 4249 302
rect 4305 246 4391 302
rect 4447 246 4533 302
rect 4589 246 4675 302
rect 4731 246 4817 302
rect 4873 246 4959 302
rect 5015 246 5101 302
rect 5157 246 5243 302
rect 5299 246 5385 302
rect 5441 246 5527 302
rect 5583 246 5669 302
rect 5725 246 5811 302
rect 5867 246 5953 302
rect 6009 246 6095 302
rect 6151 246 6237 302
rect 6293 246 6379 302
rect 6435 246 6521 302
rect 6577 246 6663 302
rect 6719 246 6805 302
rect 6861 246 6947 302
rect 7003 246 7089 302
rect 7145 246 7231 302
rect 7287 246 7373 302
rect 7429 246 7515 302
rect 7571 246 7657 302
rect 7713 246 7799 302
rect 7855 246 7941 302
rect 7997 246 8083 302
rect 8139 246 8225 302
rect 8281 246 8367 302
rect 8423 246 8509 302
rect 8565 246 8651 302
rect 8707 246 8793 302
rect 8849 246 8935 302
rect 8991 246 9077 302
rect 9133 246 9219 302
rect 9275 246 9361 302
rect 9417 246 9503 302
rect 9559 246 9645 302
rect 9701 246 9787 302
rect 9843 246 9929 302
rect 9985 246 10071 302
rect 10127 246 10213 302
rect 10269 246 10355 302
rect 10411 246 10497 302
rect 10553 246 10639 302
rect 10695 246 10781 302
rect 10837 246 10923 302
rect 10979 246 11065 302
rect 11121 246 11207 302
rect 11263 246 11349 302
rect 11405 246 11491 302
rect 11547 246 11633 302
rect 11689 246 11775 302
rect 11831 246 11917 302
rect 11973 246 12059 302
rect 12115 246 12201 302
rect 12257 246 12343 302
rect 12399 274 12526 302
rect 12582 274 12650 330
rect 12706 274 12774 330
rect 12830 274 12898 330
rect 12954 274 13022 330
rect 13078 274 13200 330
rect 12399 246 13200 274
rect -400 206 13200 246
rect -400 150 -286 206
rect -230 150 -162 206
rect -106 150 -38 206
rect 18 150 86 206
rect 142 150 210 206
rect 266 160 12526 206
rect 266 150 415 160
rect -400 104 415 150
rect 471 104 557 160
rect 613 104 699 160
rect 755 104 841 160
rect 897 104 983 160
rect 1039 104 1125 160
rect 1181 104 1267 160
rect 1323 104 1409 160
rect 1465 104 1551 160
rect 1607 104 1693 160
rect 1749 104 1835 160
rect 1891 104 1977 160
rect 2033 104 2119 160
rect 2175 104 2261 160
rect 2317 104 2403 160
rect 2459 104 2545 160
rect 2601 104 2687 160
rect 2743 104 2829 160
rect 2885 104 2971 160
rect 3027 104 3113 160
rect 3169 104 3255 160
rect 3311 104 3397 160
rect 3453 104 3539 160
rect 3595 104 3681 160
rect 3737 104 3823 160
rect 3879 104 3965 160
rect 4021 104 4107 160
rect 4163 104 4249 160
rect 4305 104 4391 160
rect 4447 104 4533 160
rect 4589 104 4675 160
rect 4731 104 4817 160
rect 4873 104 4959 160
rect 5015 104 5101 160
rect 5157 104 5243 160
rect 5299 104 5385 160
rect 5441 104 5527 160
rect 5583 104 5669 160
rect 5725 104 5811 160
rect 5867 104 5953 160
rect 6009 104 6095 160
rect 6151 104 6237 160
rect 6293 104 6379 160
rect 6435 104 6521 160
rect 6577 104 6663 160
rect 6719 104 6805 160
rect 6861 104 6947 160
rect 7003 104 7089 160
rect 7145 104 7231 160
rect 7287 104 7373 160
rect 7429 104 7515 160
rect 7571 104 7657 160
rect 7713 104 7799 160
rect 7855 104 7941 160
rect 7997 104 8083 160
rect 8139 104 8225 160
rect 8281 104 8367 160
rect 8423 104 8509 160
rect 8565 104 8651 160
rect 8707 104 8793 160
rect 8849 104 8935 160
rect 8991 104 9077 160
rect 9133 104 9219 160
rect 9275 104 9361 160
rect 9417 104 9503 160
rect 9559 104 9645 160
rect 9701 104 9787 160
rect 9843 104 9929 160
rect 9985 104 10071 160
rect 10127 104 10213 160
rect 10269 104 10355 160
rect 10411 104 10497 160
rect 10553 104 10639 160
rect 10695 104 10781 160
rect 10837 104 10923 160
rect 10979 104 11065 160
rect 11121 104 11207 160
rect 11263 104 11349 160
rect 11405 104 11491 160
rect 11547 104 11633 160
rect 11689 104 11775 160
rect 11831 104 11917 160
rect 11973 104 12059 160
rect 12115 104 12201 160
rect 12257 104 12343 160
rect 12399 150 12526 160
rect 12582 150 12650 206
rect 12706 150 12774 206
rect 12830 150 12898 206
rect 12954 150 13022 206
rect 13078 150 13200 206
rect 12399 104 13200 150
rect -400 0 13200 104
<< via4 >>
rect -254 12893 -198 12949
rect -130 12893 -74 12949
rect -6 12893 50 12949
rect 118 12893 174 12949
rect 242 12893 298 12949
rect 366 12893 422 12949
rect 490 12893 546 12949
rect 614 12893 670 12949
rect 738 12893 794 12949
rect 862 12893 918 12949
rect 986 12893 1042 12949
rect 1110 12893 1166 12949
rect 1234 12893 1290 12949
rect 1358 12893 1414 12949
rect 1482 12893 1538 12949
rect 1606 12893 1662 12949
rect 1730 12893 1786 12949
rect 1854 12893 1910 12949
rect 1978 12893 2034 12949
rect 2102 12893 2158 12949
rect 2226 12893 2282 12949
rect 2350 12893 2406 12949
rect 2474 12893 2530 12949
rect 2598 12893 2654 12949
rect 2722 12893 2778 12949
rect 2846 12893 2902 12949
rect 2970 12893 3026 12949
rect 3094 12893 3150 12949
rect 3218 12893 3274 12949
rect 3342 12893 3398 12949
rect 3466 12893 3522 12949
rect 3590 12893 3646 12949
rect 3714 12893 3770 12949
rect 3838 12893 3894 12949
rect 3962 12893 4018 12949
rect 4086 12893 4142 12949
rect 4210 12893 4266 12949
rect 4334 12893 4390 12949
rect 4458 12893 4514 12949
rect 4582 12893 4638 12949
rect 4706 12893 4762 12949
rect 4830 12893 4886 12949
rect 4954 12893 5010 12949
rect 5078 12893 5134 12949
rect 5202 12893 5258 12949
rect 5326 12893 5382 12949
rect 5450 12893 5506 12949
rect 5574 12893 5630 12949
rect 5698 12893 5754 12949
rect 5822 12893 5878 12949
rect 5946 12893 6002 12949
rect 6070 12893 6126 12949
rect 6194 12893 6250 12949
rect 6318 12893 6374 12949
rect 6442 12893 6498 12949
rect 6566 12893 6622 12949
rect 6690 12893 6746 12949
rect 6814 12893 6870 12949
rect 6938 12893 6994 12949
rect 7062 12893 7118 12949
rect 7186 12893 7242 12949
rect 7310 12893 7366 12949
rect 7434 12893 7490 12949
rect 7558 12893 7614 12949
rect 7682 12893 7738 12949
rect 7806 12893 7862 12949
rect 7930 12893 7986 12949
rect 8054 12893 8110 12949
rect 8178 12893 8234 12949
rect 8302 12893 8358 12949
rect 8426 12893 8482 12949
rect 8550 12893 8606 12949
rect 8674 12893 8730 12949
rect 8798 12893 8854 12949
rect 8922 12893 8978 12949
rect 9046 12893 9102 12949
rect 9170 12893 9226 12949
rect 9294 12893 9350 12949
rect 9418 12893 9474 12949
rect 9542 12893 9598 12949
rect 9666 12893 9722 12949
rect 9790 12893 9846 12949
rect 9914 12893 9970 12949
rect 10038 12893 10094 12949
rect 10162 12893 10218 12949
rect 10286 12893 10342 12949
rect 10410 12893 10466 12949
rect 10534 12893 10590 12949
rect 10658 12893 10714 12949
rect 10782 12893 10838 12949
rect 10906 12893 10962 12949
rect 11030 12893 11086 12949
rect 11154 12893 11210 12949
rect 11278 12893 11334 12949
rect 11402 12893 11458 12949
rect 11526 12893 11582 12949
rect 11650 12893 11706 12949
rect 11774 12893 11830 12949
rect 11898 12893 11954 12949
rect 12022 12893 12078 12949
rect 12146 12893 12202 12949
rect 12270 12893 12326 12949
rect 12394 12893 12450 12949
rect 12518 12893 12574 12949
rect 12642 12893 12698 12949
rect 12766 12893 12822 12949
rect 12890 12893 12946 12949
rect 13014 12893 13070 12949
rect -254 12769 -198 12825
rect -130 12769 -74 12825
rect -6 12769 50 12825
rect 118 12769 174 12825
rect 242 12769 298 12825
rect 366 12769 422 12825
rect 490 12769 546 12825
rect 614 12769 670 12825
rect 738 12769 794 12825
rect 862 12769 918 12825
rect 986 12769 1042 12825
rect 1110 12769 1166 12825
rect 1234 12769 1290 12825
rect 1358 12769 1414 12825
rect 1482 12769 1538 12825
rect 1606 12769 1662 12825
rect 1730 12769 1786 12825
rect 1854 12769 1910 12825
rect 1978 12769 2034 12825
rect 2102 12769 2158 12825
rect 2226 12769 2282 12825
rect 2350 12769 2406 12825
rect 2474 12769 2530 12825
rect 2598 12769 2654 12825
rect 2722 12769 2778 12825
rect 2846 12769 2902 12825
rect 2970 12769 3026 12825
rect 3094 12769 3150 12825
rect 3218 12769 3274 12825
rect 3342 12769 3398 12825
rect 3466 12769 3522 12825
rect 3590 12769 3646 12825
rect 3714 12769 3770 12825
rect 3838 12769 3894 12825
rect 3962 12769 4018 12825
rect 4086 12769 4142 12825
rect 4210 12769 4266 12825
rect 4334 12769 4390 12825
rect 4458 12769 4514 12825
rect 4582 12769 4638 12825
rect 4706 12769 4762 12825
rect 4830 12769 4886 12825
rect 4954 12769 5010 12825
rect 5078 12769 5134 12825
rect 5202 12769 5258 12825
rect 5326 12769 5382 12825
rect 5450 12769 5506 12825
rect 5574 12769 5630 12825
rect 5698 12769 5754 12825
rect 5822 12769 5878 12825
rect 5946 12769 6002 12825
rect 6070 12769 6126 12825
rect 6194 12769 6250 12825
rect 6318 12769 6374 12825
rect 6442 12769 6498 12825
rect 6566 12769 6622 12825
rect 6690 12769 6746 12825
rect 6814 12769 6870 12825
rect 6938 12769 6994 12825
rect 7062 12769 7118 12825
rect 7186 12769 7242 12825
rect 7310 12769 7366 12825
rect 7434 12769 7490 12825
rect 7558 12769 7614 12825
rect 7682 12769 7738 12825
rect 7806 12769 7862 12825
rect 7930 12769 7986 12825
rect 8054 12769 8110 12825
rect 8178 12769 8234 12825
rect 8302 12769 8358 12825
rect 8426 12769 8482 12825
rect 8550 12769 8606 12825
rect 8674 12769 8730 12825
rect 8798 12769 8854 12825
rect 8922 12769 8978 12825
rect 9046 12769 9102 12825
rect 9170 12769 9226 12825
rect 9294 12769 9350 12825
rect 9418 12769 9474 12825
rect 9542 12769 9598 12825
rect 9666 12769 9722 12825
rect 9790 12769 9846 12825
rect 9914 12769 9970 12825
rect 10038 12769 10094 12825
rect 10162 12769 10218 12825
rect 10286 12769 10342 12825
rect 10410 12769 10466 12825
rect 10534 12769 10590 12825
rect 10658 12769 10714 12825
rect 10782 12769 10838 12825
rect 10906 12769 10962 12825
rect 11030 12769 11086 12825
rect 11154 12769 11210 12825
rect 11278 12769 11334 12825
rect 11402 12769 11458 12825
rect 11526 12769 11582 12825
rect 11650 12769 11706 12825
rect 11774 12769 11830 12825
rect 11898 12769 11954 12825
rect 12022 12769 12078 12825
rect 12146 12769 12202 12825
rect 12270 12769 12326 12825
rect 12394 12769 12450 12825
rect 12518 12769 12574 12825
rect 12642 12769 12698 12825
rect 12766 12769 12822 12825
rect 12890 12769 12946 12825
rect 13014 12769 13070 12825
rect -254 12645 -198 12701
rect -130 12645 -74 12701
rect -6 12645 50 12701
rect 118 12645 174 12701
rect 242 12645 298 12701
rect 366 12645 422 12701
rect 490 12645 546 12701
rect 614 12645 670 12701
rect 738 12645 794 12701
rect 862 12645 918 12701
rect 986 12645 1042 12701
rect 1110 12645 1166 12701
rect 1234 12645 1290 12701
rect 1358 12645 1414 12701
rect 1482 12645 1538 12701
rect 1606 12645 1662 12701
rect 1730 12645 1786 12701
rect 1854 12645 1910 12701
rect 1978 12645 2034 12701
rect 2102 12645 2158 12701
rect 2226 12645 2282 12701
rect 2350 12645 2406 12701
rect 2474 12645 2530 12701
rect 2598 12645 2654 12701
rect 2722 12645 2778 12701
rect 2846 12645 2902 12701
rect 2970 12645 3026 12701
rect 3094 12645 3150 12701
rect 3218 12645 3274 12701
rect 3342 12645 3398 12701
rect 3466 12645 3522 12701
rect 3590 12645 3646 12701
rect 3714 12645 3770 12701
rect 3838 12645 3894 12701
rect 3962 12645 4018 12701
rect 4086 12645 4142 12701
rect 4210 12645 4266 12701
rect 4334 12645 4390 12701
rect 4458 12645 4514 12701
rect 4582 12645 4638 12701
rect 4706 12645 4762 12701
rect 4830 12645 4886 12701
rect 4954 12645 5010 12701
rect 5078 12645 5134 12701
rect 5202 12645 5258 12701
rect 5326 12645 5382 12701
rect 5450 12645 5506 12701
rect 5574 12645 5630 12701
rect 5698 12645 5754 12701
rect 5822 12645 5878 12701
rect 5946 12645 6002 12701
rect 6070 12645 6126 12701
rect 6194 12645 6250 12701
rect 6318 12645 6374 12701
rect 6442 12645 6498 12701
rect 6566 12645 6622 12701
rect 6690 12645 6746 12701
rect 6814 12645 6870 12701
rect 6938 12645 6994 12701
rect 7062 12645 7118 12701
rect 7186 12645 7242 12701
rect 7310 12645 7366 12701
rect 7434 12645 7490 12701
rect 7558 12645 7614 12701
rect 7682 12645 7738 12701
rect 7806 12645 7862 12701
rect 7930 12645 7986 12701
rect 8054 12645 8110 12701
rect 8178 12645 8234 12701
rect 8302 12645 8358 12701
rect 8426 12645 8482 12701
rect 8550 12645 8606 12701
rect 8674 12645 8730 12701
rect 8798 12645 8854 12701
rect 8922 12645 8978 12701
rect 9046 12645 9102 12701
rect 9170 12645 9226 12701
rect 9294 12645 9350 12701
rect 9418 12645 9474 12701
rect 9542 12645 9598 12701
rect 9666 12645 9722 12701
rect 9790 12645 9846 12701
rect 9914 12645 9970 12701
rect 10038 12645 10094 12701
rect 10162 12645 10218 12701
rect 10286 12645 10342 12701
rect 10410 12645 10466 12701
rect 10534 12645 10590 12701
rect 10658 12645 10714 12701
rect 10782 12645 10838 12701
rect 10906 12645 10962 12701
rect 11030 12645 11086 12701
rect 11154 12645 11210 12701
rect 11278 12645 11334 12701
rect 11402 12645 11458 12701
rect 11526 12645 11582 12701
rect 11650 12645 11706 12701
rect 11774 12645 11830 12701
rect 11898 12645 11954 12701
rect 12022 12645 12078 12701
rect 12146 12645 12202 12701
rect 12270 12645 12326 12701
rect 12394 12645 12450 12701
rect 12518 12645 12574 12701
rect 12642 12645 12698 12701
rect 12766 12645 12822 12701
rect 12890 12645 12946 12701
rect 13014 12645 13070 12701
rect -254 12521 -198 12577
rect -130 12521 -74 12577
rect -6 12521 50 12577
rect 118 12521 174 12577
rect 242 12521 298 12577
rect 366 12521 422 12577
rect 490 12521 546 12577
rect 614 12521 670 12577
rect 738 12521 794 12577
rect 862 12521 918 12577
rect 986 12521 1042 12577
rect 1110 12521 1166 12577
rect 1234 12521 1290 12577
rect 1358 12521 1414 12577
rect 1482 12521 1538 12577
rect 1606 12521 1662 12577
rect 1730 12521 1786 12577
rect 1854 12521 1910 12577
rect 1978 12521 2034 12577
rect 2102 12521 2158 12577
rect 2226 12521 2282 12577
rect 2350 12521 2406 12577
rect 2474 12521 2530 12577
rect 2598 12521 2654 12577
rect 2722 12521 2778 12577
rect 2846 12521 2902 12577
rect 2970 12521 3026 12577
rect 3094 12521 3150 12577
rect 3218 12521 3274 12577
rect 3342 12521 3398 12577
rect 3466 12521 3522 12577
rect 3590 12521 3646 12577
rect 3714 12521 3770 12577
rect 3838 12521 3894 12577
rect 3962 12521 4018 12577
rect 4086 12521 4142 12577
rect 4210 12521 4266 12577
rect 4334 12521 4390 12577
rect 4458 12521 4514 12577
rect 4582 12521 4638 12577
rect 4706 12521 4762 12577
rect 4830 12521 4886 12577
rect 4954 12521 5010 12577
rect 5078 12521 5134 12577
rect 5202 12521 5258 12577
rect 5326 12521 5382 12577
rect 5450 12521 5506 12577
rect 5574 12521 5630 12577
rect 5698 12521 5754 12577
rect 5822 12521 5878 12577
rect 5946 12521 6002 12577
rect 6070 12521 6126 12577
rect 6194 12521 6250 12577
rect 6318 12521 6374 12577
rect 6442 12521 6498 12577
rect 6566 12521 6622 12577
rect 6690 12521 6746 12577
rect 6814 12521 6870 12577
rect 6938 12521 6994 12577
rect 7062 12521 7118 12577
rect 7186 12521 7242 12577
rect 7310 12521 7366 12577
rect 7434 12521 7490 12577
rect 7558 12521 7614 12577
rect 7682 12521 7738 12577
rect 7806 12521 7862 12577
rect 7930 12521 7986 12577
rect 8054 12521 8110 12577
rect 8178 12521 8234 12577
rect 8302 12521 8358 12577
rect 8426 12521 8482 12577
rect 8550 12521 8606 12577
rect 8674 12521 8730 12577
rect 8798 12521 8854 12577
rect 8922 12521 8978 12577
rect 9046 12521 9102 12577
rect 9170 12521 9226 12577
rect 9294 12521 9350 12577
rect 9418 12521 9474 12577
rect 9542 12521 9598 12577
rect 9666 12521 9722 12577
rect 9790 12521 9846 12577
rect 9914 12521 9970 12577
rect 10038 12521 10094 12577
rect 10162 12521 10218 12577
rect 10286 12521 10342 12577
rect 10410 12521 10466 12577
rect 10534 12521 10590 12577
rect 10658 12521 10714 12577
rect 10782 12521 10838 12577
rect 10906 12521 10962 12577
rect 11030 12521 11086 12577
rect 11154 12521 11210 12577
rect 11278 12521 11334 12577
rect 11402 12521 11458 12577
rect 11526 12521 11582 12577
rect 11650 12521 11706 12577
rect 11774 12521 11830 12577
rect 11898 12521 11954 12577
rect 12022 12521 12078 12577
rect 12146 12521 12202 12577
rect 12270 12521 12326 12577
rect 12394 12521 12450 12577
rect 12518 12521 12574 12577
rect 12642 12521 12698 12577
rect 12766 12521 12822 12577
rect 12890 12521 12946 12577
rect 13014 12521 13070 12577
rect -286 12302 -230 12358
rect -162 12302 -106 12358
rect -38 12302 18 12358
rect 86 12302 142 12358
rect 210 12302 266 12358
rect -286 12178 -230 12234
rect -162 12178 -106 12234
rect -38 12178 18 12234
rect 86 12178 142 12234
rect 210 12178 266 12234
rect -286 12054 -230 12110
rect -162 12054 -106 12110
rect -38 12054 18 12110
rect 86 12054 142 12110
rect 210 12054 266 12110
rect -286 11930 -230 11986
rect -162 11930 -106 11986
rect -38 11930 18 11986
rect 86 11930 142 11986
rect 210 11930 266 11986
rect -286 11806 -230 11862
rect -162 11806 -106 11862
rect -38 11806 18 11862
rect 86 11806 142 11862
rect 210 11806 266 11862
rect -286 11682 -230 11738
rect -162 11682 -106 11738
rect -38 11682 18 11738
rect 86 11682 142 11738
rect 210 11682 266 11738
rect -286 11558 -230 11614
rect -162 11558 -106 11614
rect -38 11558 18 11614
rect 86 11558 142 11614
rect 210 11558 266 11614
rect -286 11434 -230 11490
rect -162 11434 -106 11490
rect -38 11434 18 11490
rect 86 11434 142 11490
rect 210 11434 266 11490
rect -286 11310 -230 11366
rect -162 11310 -106 11366
rect -38 11310 18 11366
rect 86 11310 142 11366
rect 210 11310 266 11366
rect -286 11186 -230 11242
rect -162 11186 -106 11242
rect -38 11186 18 11242
rect 86 11186 142 11242
rect 210 11186 266 11242
rect -286 11062 -230 11118
rect -162 11062 -106 11118
rect -38 11062 18 11118
rect 86 11062 142 11118
rect 210 11062 266 11118
rect -286 10938 -230 10994
rect -162 10938 -106 10994
rect -38 10938 18 10994
rect 86 10938 142 10994
rect 210 10938 266 10994
rect -286 10814 -230 10870
rect -162 10814 -106 10870
rect -38 10814 18 10870
rect 86 10814 142 10870
rect 210 10814 266 10870
rect -286 10690 -230 10746
rect -162 10690 -106 10746
rect -38 10690 18 10746
rect 86 10690 142 10746
rect 210 10690 266 10746
rect -286 10566 -230 10622
rect -162 10566 -106 10622
rect -38 10566 18 10622
rect 86 10566 142 10622
rect 210 10566 266 10622
rect -286 10442 -230 10498
rect -162 10442 -106 10498
rect -38 10442 18 10498
rect 86 10442 142 10498
rect 210 10442 266 10498
rect -286 10318 -230 10374
rect -162 10318 -106 10374
rect -38 10318 18 10374
rect 86 10318 142 10374
rect 210 10318 266 10374
rect -286 10194 -230 10250
rect -162 10194 -106 10250
rect -38 10194 18 10250
rect 86 10194 142 10250
rect 210 10194 266 10250
rect -286 10070 -230 10126
rect -162 10070 -106 10126
rect -38 10070 18 10126
rect 86 10070 142 10126
rect 210 10070 266 10126
rect -286 9946 -230 10002
rect -162 9946 -106 10002
rect -38 9946 18 10002
rect 86 9946 142 10002
rect 210 9946 266 10002
rect -286 9822 -230 9878
rect -162 9822 -106 9878
rect -38 9822 18 9878
rect 86 9822 142 9878
rect 210 9822 266 9878
rect -286 9698 -230 9754
rect -162 9698 -106 9754
rect -38 9698 18 9754
rect 86 9698 142 9754
rect 210 9698 266 9754
rect -286 9574 -230 9630
rect -162 9574 -106 9630
rect -38 9574 18 9630
rect 86 9574 142 9630
rect 210 9574 266 9630
rect -286 9450 -230 9506
rect -162 9450 -106 9506
rect -38 9450 18 9506
rect 86 9450 142 9506
rect 210 9450 266 9506
rect -286 9326 -230 9382
rect -162 9326 -106 9382
rect -38 9326 18 9382
rect 86 9326 142 9382
rect 210 9326 266 9382
rect -286 9202 -230 9258
rect -162 9202 -106 9258
rect -38 9202 18 9258
rect 86 9202 142 9258
rect 210 9202 266 9258
rect -286 9078 -230 9134
rect -162 9078 -106 9134
rect -38 9078 18 9134
rect 86 9078 142 9134
rect 210 9078 266 9134
rect -286 8954 -230 9010
rect -162 8954 -106 9010
rect -38 8954 18 9010
rect 86 8954 142 9010
rect 210 8954 266 9010
rect -286 8830 -230 8886
rect -162 8830 -106 8886
rect -38 8830 18 8886
rect 86 8830 142 8886
rect 210 8830 266 8886
rect -286 8706 -230 8762
rect -162 8706 -106 8762
rect -38 8706 18 8762
rect 86 8706 142 8762
rect 210 8706 266 8762
rect -286 8582 -230 8638
rect -162 8582 -106 8638
rect -38 8582 18 8638
rect 86 8582 142 8638
rect 210 8582 266 8638
rect -286 8458 -230 8514
rect -162 8458 -106 8514
rect -38 8458 18 8514
rect 86 8458 142 8514
rect 210 8458 266 8514
rect -286 8334 -230 8390
rect -162 8334 -106 8390
rect -38 8334 18 8390
rect 86 8334 142 8390
rect 210 8334 266 8390
rect -286 8210 -230 8266
rect -162 8210 -106 8266
rect -38 8210 18 8266
rect 86 8210 142 8266
rect 210 8210 266 8266
rect -286 8086 -230 8142
rect -162 8086 -106 8142
rect -38 8086 18 8142
rect 86 8086 142 8142
rect 210 8086 266 8142
rect -286 7962 -230 8018
rect -162 7962 -106 8018
rect -38 7962 18 8018
rect 86 7962 142 8018
rect 210 7962 266 8018
rect -286 7838 -230 7894
rect -162 7838 -106 7894
rect -38 7838 18 7894
rect 86 7838 142 7894
rect 210 7838 266 7894
rect -286 7714 -230 7770
rect -162 7714 -106 7770
rect -38 7714 18 7770
rect 86 7714 142 7770
rect 210 7714 266 7770
rect -286 7590 -230 7646
rect -162 7590 -106 7646
rect -38 7590 18 7646
rect 86 7590 142 7646
rect 210 7590 266 7646
rect -286 7466 -230 7522
rect -162 7466 -106 7522
rect -38 7466 18 7522
rect 86 7466 142 7522
rect 210 7466 266 7522
rect -286 7342 -230 7398
rect -162 7342 -106 7398
rect -38 7342 18 7398
rect 86 7342 142 7398
rect 210 7342 266 7398
rect -286 7218 -230 7274
rect -162 7218 -106 7274
rect -38 7218 18 7274
rect 86 7218 142 7274
rect 210 7218 266 7274
rect -286 7094 -230 7150
rect -162 7094 -106 7150
rect -38 7094 18 7150
rect 86 7094 142 7150
rect 210 7094 266 7150
rect -286 6970 -230 7026
rect -162 6970 -106 7026
rect -38 6970 18 7026
rect 86 6970 142 7026
rect 210 6970 266 7026
rect -286 6846 -230 6902
rect -162 6846 -106 6902
rect -38 6846 18 6902
rect 86 6846 142 6902
rect 210 6846 266 6902
rect -286 6722 -230 6778
rect -162 6722 -106 6778
rect -38 6722 18 6778
rect 86 6722 142 6778
rect 210 6722 266 6778
rect -286 6598 -230 6654
rect -162 6598 -106 6654
rect -38 6598 18 6654
rect 86 6598 142 6654
rect 210 6598 266 6654
rect -286 6474 -230 6530
rect -162 6474 -106 6530
rect -38 6474 18 6530
rect 86 6474 142 6530
rect 210 6474 266 6530
rect -286 6350 -230 6406
rect -162 6350 -106 6406
rect -38 6350 18 6406
rect 86 6350 142 6406
rect 210 6350 266 6406
rect -286 6226 -230 6282
rect -162 6226 -106 6282
rect -38 6226 18 6282
rect 86 6226 142 6282
rect 210 6226 266 6282
rect -286 6102 -230 6158
rect -162 6102 -106 6158
rect -38 6102 18 6158
rect 86 6102 142 6158
rect 210 6102 266 6158
rect -286 5978 -230 6034
rect -162 5978 -106 6034
rect -38 5978 18 6034
rect 86 5978 142 6034
rect 210 5978 266 6034
rect -286 5854 -230 5910
rect -162 5854 -106 5910
rect -38 5854 18 5910
rect 86 5854 142 5910
rect 210 5854 266 5910
rect -286 5730 -230 5786
rect -162 5730 -106 5786
rect -38 5730 18 5786
rect 86 5730 142 5786
rect 210 5730 266 5786
rect -286 5606 -230 5662
rect -162 5606 -106 5662
rect -38 5606 18 5662
rect 86 5606 142 5662
rect 210 5606 266 5662
rect -286 5482 -230 5538
rect -162 5482 -106 5538
rect -38 5482 18 5538
rect 86 5482 142 5538
rect 210 5482 266 5538
rect -286 5358 -230 5414
rect -162 5358 -106 5414
rect -38 5358 18 5414
rect 86 5358 142 5414
rect 210 5358 266 5414
rect -286 5234 -230 5290
rect -162 5234 -106 5290
rect -38 5234 18 5290
rect 86 5234 142 5290
rect 210 5234 266 5290
rect -286 5110 -230 5166
rect -162 5110 -106 5166
rect -38 5110 18 5166
rect 86 5110 142 5166
rect 210 5110 266 5166
rect -286 4986 -230 5042
rect -162 4986 -106 5042
rect -38 4986 18 5042
rect 86 4986 142 5042
rect 210 4986 266 5042
rect -286 4862 -230 4918
rect -162 4862 -106 4918
rect -38 4862 18 4918
rect 86 4862 142 4918
rect 210 4862 266 4918
rect -286 4738 -230 4794
rect -162 4738 -106 4794
rect -38 4738 18 4794
rect 86 4738 142 4794
rect 210 4738 266 4794
rect -286 4614 -230 4670
rect -162 4614 -106 4670
rect -38 4614 18 4670
rect 86 4614 142 4670
rect 210 4614 266 4670
rect -286 4490 -230 4546
rect -162 4490 -106 4546
rect -38 4490 18 4546
rect 86 4490 142 4546
rect 210 4490 266 4546
rect -286 4366 -230 4422
rect -162 4366 -106 4422
rect -38 4366 18 4422
rect 86 4366 142 4422
rect 210 4366 266 4422
rect -286 4242 -230 4298
rect -162 4242 -106 4298
rect -38 4242 18 4298
rect 86 4242 142 4298
rect 210 4242 266 4298
rect -286 4118 -230 4174
rect -162 4118 -106 4174
rect -38 4118 18 4174
rect 86 4118 142 4174
rect 210 4118 266 4174
rect -286 3994 -230 4050
rect -162 3994 -106 4050
rect -38 3994 18 4050
rect 86 3994 142 4050
rect 210 3994 266 4050
rect -286 3870 -230 3926
rect -162 3870 -106 3926
rect -38 3870 18 3926
rect 86 3870 142 3926
rect 210 3870 266 3926
rect -286 3746 -230 3802
rect -162 3746 -106 3802
rect -38 3746 18 3802
rect 86 3746 142 3802
rect 210 3746 266 3802
rect -286 3622 -230 3678
rect -162 3622 -106 3678
rect -38 3622 18 3678
rect 86 3622 142 3678
rect 210 3622 266 3678
rect -286 3498 -230 3554
rect -162 3498 -106 3554
rect -38 3498 18 3554
rect 86 3498 142 3554
rect 210 3498 266 3554
rect -286 3374 -230 3430
rect -162 3374 -106 3430
rect -38 3374 18 3430
rect 86 3374 142 3430
rect 210 3374 266 3430
rect -286 3250 -230 3306
rect -162 3250 -106 3306
rect -38 3250 18 3306
rect 86 3250 142 3306
rect 210 3250 266 3306
rect -286 3126 -230 3182
rect -162 3126 -106 3182
rect -38 3126 18 3182
rect 86 3126 142 3182
rect 210 3126 266 3182
rect -286 3002 -230 3058
rect -162 3002 -106 3058
rect -38 3002 18 3058
rect 86 3002 142 3058
rect 210 3002 266 3058
rect -286 2878 -230 2934
rect -162 2878 -106 2934
rect -38 2878 18 2934
rect 86 2878 142 2934
rect 210 2878 266 2934
rect -286 2754 -230 2810
rect -162 2754 -106 2810
rect -38 2754 18 2810
rect 86 2754 142 2810
rect 210 2754 266 2810
rect -286 2630 -230 2686
rect -162 2630 -106 2686
rect -38 2630 18 2686
rect 86 2630 142 2686
rect 210 2630 266 2686
rect -286 2506 -230 2562
rect -162 2506 -106 2562
rect -38 2506 18 2562
rect 86 2506 142 2562
rect 210 2506 266 2562
rect -286 2382 -230 2438
rect -162 2382 -106 2438
rect -38 2382 18 2438
rect 86 2382 142 2438
rect 210 2382 266 2438
rect -286 2258 -230 2314
rect -162 2258 -106 2314
rect -38 2258 18 2314
rect 86 2258 142 2314
rect 210 2258 266 2314
rect -286 2134 -230 2190
rect -162 2134 -106 2190
rect -38 2134 18 2190
rect 86 2134 142 2190
rect 210 2134 266 2190
rect -286 2010 -230 2066
rect -162 2010 -106 2066
rect -38 2010 18 2066
rect 86 2010 142 2066
rect 210 2010 266 2066
rect -286 1886 -230 1942
rect -162 1886 -106 1942
rect -38 1886 18 1942
rect 86 1886 142 1942
rect 210 1886 266 1942
rect -286 1762 -230 1818
rect -162 1762 -106 1818
rect -38 1762 18 1818
rect 86 1762 142 1818
rect 210 1762 266 1818
rect -286 1638 -230 1694
rect -162 1638 -106 1694
rect -38 1638 18 1694
rect 86 1638 142 1694
rect 210 1638 266 1694
rect -286 1514 -230 1570
rect -162 1514 -106 1570
rect -38 1514 18 1570
rect 86 1514 142 1570
rect 210 1514 266 1570
rect -286 1390 -230 1446
rect -162 1390 -106 1446
rect -38 1390 18 1446
rect 86 1390 142 1446
rect 210 1390 266 1446
rect -286 1266 -230 1322
rect -162 1266 -106 1322
rect -38 1266 18 1322
rect 86 1266 142 1322
rect 210 1266 266 1322
rect -286 1142 -230 1198
rect -162 1142 -106 1198
rect -38 1142 18 1198
rect 86 1142 142 1198
rect 210 1142 266 1198
rect -286 1018 -230 1074
rect -162 1018 -106 1074
rect -38 1018 18 1074
rect 86 1018 142 1074
rect 210 1018 266 1074
rect -286 894 -230 950
rect -162 894 -106 950
rect -38 894 18 950
rect 86 894 142 950
rect 210 894 266 950
rect -286 770 -230 826
rect -162 770 -106 826
rect -38 770 18 826
rect 86 770 142 826
rect 210 770 266 826
rect -286 646 -230 702
rect -162 646 -106 702
rect -38 646 18 702
rect 86 646 142 702
rect 210 646 266 702
rect -286 522 -230 578
rect -162 522 -106 578
rect -38 522 18 578
rect 86 522 142 578
rect 210 522 266 578
rect 903 12254 959 12310
rect 1045 12254 1101 12310
rect 903 12112 959 12168
rect 1045 12112 1101 12168
rect 903 11970 959 12026
rect 1045 11970 1101 12026
rect 903 11828 959 11884
rect 1045 11828 1101 11884
rect 903 11686 959 11742
rect 1045 11686 1101 11742
rect 903 11544 959 11600
rect 1045 11544 1101 11600
rect 903 11402 959 11458
rect 1045 11402 1101 11458
rect 903 11260 959 11316
rect 1045 11260 1101 11316
rect 903 11118 959 11174
rect 1045 11118 1101 11174
rect 903 10976 959 11032
rect 1045 10976 1101 11032
rect 903 10834 959 10890
rect 1045 10834 1101 10890
rect 903 10692 959 10748
rect 1045 10692 1101 10748
rect 903 10550 959 10606
rect 1045 10550 1101 10606
rect 903 10408 959 10464
rect 1045 10408 1101 10464
rect 903 10266 959 10322
rect 1045 10266 1101 10322
rect 903 10124 959 10180
rect 1045 10124 1101 10180
rect 903 9982 959 10038
rect 1045 9982 1101 10038
rect 903 9840 959 9896
rect 1045 9840 1101 9896
rect 903 9698 959 9754
rect 1045 9698 1101 9754
rect 903 9556 959 9612
rect 1045 9556 1101 9612
rect 903 9414 959 9470
rect 1045 9414 1101 9470
rect 903 9272 959 9328
rect 1045 9272 1101 9328
rect 903 9130 959 9186
rect 1045 9130 1101 9186
rect 903 8988 959 9044
rect 1045 8988 1101 9044
rect 903 8846 959 8902
rect 1045 8846 1101 8902
rect 903 8704 959 8760
rect 1045 8704 1101 8760
rect 903 8562 959 8618
rect 1045 8562 1101 8618
rect 903 8420 959 8476
rect 1045 8420 1101 8476
rect 903 8278 959 8334
rect 1045 8278 1101 8334
rect 903 8136 959 8192
rect 1045 8136 1101 8192
rect 903 7994 959 8050
rect 1045 7994 1101 8050
rect 903 7852 959 7908
rect 1045 7852 1101 7908
rect 903 7710 959 7766
rect 1045 7710 1101 7766
rect 903 7568 959 7624
rect 1045 7568 1101 7624
rect 903 7426 959 7482
rect 1045 7426 1101 7482
rect 903 7284 959 7340
rect 1045 7284 1101 7340
rect 903 7142 959 7198
rect 1045 7142 1101 7198
rect 903 7000 959 7056
rect 1045 7000 1101 7056
rect 903 6858 959 6914
rect 1045 6858 1101 6914
rect 903 6716 959 6772
rect 1045 6716 1101 6772
rect 903 6574 959 6630
rect 1045 6574 1101 6630
rect 903 6432 959 6488
rect 1045 6432 1101 6488
rect 903 6290 959 6346
rect 1045 6290 1101 6346
rect 903 6148 959 6204
rect 1045 6148 1101 6204
rect 903 6006 959 6062
rect 1045 6006 1101 6062
rect 903 5864 959 5920
rect 1045 5864 1101 5920
rect 903 5722 959 5778
rect 1045 5722 1101 5778
rect 903 5580 959 5636
rect 1045 5580 1101 5636
rect 903 5438 959 5494
rect 1045 5438 1101 5494
rect 903 5296 959 5352
rect 1045 5296 1101 5352
rect 903 5154 959 5210
rect 1045 5154 1101 5210
rect 903 5012 959 5068
rect 1045 5012 1101 5068
rect 903 4870 959 4926
rect 1045 4870 1101 4926
rect 903 4728 959 4784
rect 1045 4728 1101 4784
rect 903 4586 959 4642
rect 1045 4586 1101 4642
rect 903 4444 959 4500
rect 1045 4444 1101 4500
rect 903 4302 959 4358
rect 1045 4302 1101 4358
rect 903 4160 959 4216
rect 1045 4160 1101 4216
rect 903 4018 959 4074
rect 1045 4018 1101 4074
rect 903 3876 959 3932
rect 1045 3876 1101 3932
rect 903 3734 959 3790
rect 1045 3734 1101 3790
rect 903 3592 959 3648
rect 1045 3592 1101 3648
rect 903 3450 959 3506
rect 1045 3450 1101 3506
rect 903 3308 959 3364
rect 1045 3308 1101 3364
rect 903 3166 959 3222
rect 1045 3166 1101 3222
rect 903 3024 959 3080
rect 1045 3024 1101 3080
rect 903 2882 959 2938
rect 1045 2882 1101 2938
rect 903 2740 959 2796
rect 1045 2740 1101 2796
rect 903 2598 959 2654
rect 1045 2598 1101 2654
rect 903 2456 959 2512
rect 1045 2456 1101 2512
rect 903 2314 959 2370
rect 1045 2314 1101 2370
rect 903 2172 959 2228
rect 1045 2172 1101 2228
rect 903 2030 959 2086
rect 1045 2030 1101 2086
rect 903 1888 959 1944
rect 1045 1888 1101 1944
rect 903 1746 959 1802
rect 1045 1746 1101 1802
rect 903 1604 959 1660
rect 1045 1604 1101 1660
rect 903 1462 959 1518
rect 1045 1462 1101 1518
rect 903 1320 959 1376
rect 1045 1320 1101 1376
rect 903 1178 959 1234
rect 1045 1178 1101 1234
rect 903 1036 959 1092
rect 1045 1036 1101 1092
rect 903 894 959 950
rect 1045 894 1101 950
rect 903 752 959 808
rect 1045 752 1101 808
rect 903 610 959 666
rect 1045 610 1101 666
rect 903 468 959 524
rect 1045 468 1101 524
rect 1444 12254 1500 12310
rect 1586 12254 1642 12310
rect 1444 12112 1500 12168
rect 1586 12112 1642 12168
rect 1444 11970 1500 12026
rect 1586 11970 1642 12026
rect 1444 11828 1500 11884
rect 1586 11828 1642 11884
rect 1444 11686 1500 11742
rect 1586 11686 1642 11742
rect 1444 11544 1500 11600
rect 1586 11544 1642 11600
rect 1444 11402 1500 11458
rect 1586 11402 1642 11458
rect 1444 11260 1500 11316
rect 1586 11260 1642 11316
rect 1444 11118 1500 11174
rect 1586 11118 1642 11174
rect 1444 10976 1500 11032
rect 1586 10976 1642 11032
rect 1444 10834 1500 10890
rect 1586 10834 1642 10890
rect 1444 10692 1500 10748
rect 1586 10692 1642 10748
rect 1444 10550 1500 10606
rect 1586 10550 1642 10606
rect 1444 10408 1500 10464
rect 1586 10408 1642 10464
rect 1444 10266 1500 10322
rect 1586 10266 1642 10322
rect 1444 10124 1500 10180
rect 1586 10124 1642 10180
rect 1444 9982 1500 10038
rect 1586 9982 1642 10038
rect 1444 9840 1500 9896
rect 1586 9840 1642 9896
rect 1444 9698 1500 9754
rect 1586 9698 1642 9754
rect 1444 9556 1500 9612
rect 1586 9556 1642 9612
rect 1444 9414 1500 9470
rect 1586 9414 1642 9470
rect 1444 9272 1500 9328
rect 1586 9272 1642 9328
rect 1444 9130 1500 9186
rect 1586 9130 1642 9186
rect 1444 8988 1500 9044
rect 1586 8988 1642 9044
rect 1444 8846 1500 8902
rect 1586 8846 1642 8902
rect 1444 8704 1500 8760
rect 1586 8704 1642 8760
rect 1444 8562 1500 8618
rect 1586 8562 1642 8618
rect 1444 8420 1500 8476
rect 1586 8420 1642 8476
rect 1444 8278 1500 8334
rect 1586 8278 1642 8334
rect 1444 8136 1500 8192
rect 1586 8136 1642 8192
rect 1444 7994 1500 8050
rect 1586 7994 1642 8050
rect 1444 7852 1500 7908
rect 1586 7852 1642 7908
rect 1444 7710 1500 7766
rect 1586 7710 1642 7766
rect 1444 7568 1500 7624
rect 1586 7568 1642 7624
rect 1444 7426 1500 7482
rect 1586 7426 1642 7482
rect 1444 7284 1500 7340
rect 1586 7284 1642 7340
rect 1444 7142 1500 7198
rect 1586 7142 1642 7198
rect 1444 7000 1500 7056
rect 1586 7000 1642 7056
rect 1444 6858 1500 6914
rect 1586 6858 1642 6914
rect 1444 6716 1500 6772
rect 1586 6716 1642 6772
rect 1444 6574 1500 6630
rect 1586 6574 1642 6630
rect 1444 6432 1500 6488
rect 1586 6432 1642 6488
rect 1444 6290 1500 6346
rect 1586 6290 1642 6346
rect 1444 6148 1500 6204
rect 1586 6148 1642 6204
rect 1444 6006 1500 6062
rect 1586 6006 1642 6062
rect 1444 5864 1500 5920
rect 1586 5864 1642 5920
rect 1444 5722 1500 5778
rect 1586 5722 1642 5778
rect 1444 5580 1500 5636
rect 1586 5580 1642 5636
rect 1444 5438 1500 5494
rect 1586 5438 1642 5494
rect 1444 5296 1500 5352
rect 1586 5296 1642 5352
rect 1444 5154 1500 5210
rect 1586 5154 1642 5210
rect 1444 5012 1500 5068
rect 1586 5012 1642 5068
rect 1444 4870 1500 4926
rect 1586 4870 1642 4926
rect 1444 4728 1500 4784
rect 1586 4728 1642 4784
rect 1444 4586 1500 4642
rect 1586 4586 1642 4642
rect 1444 4444 1500 4500
rect 1586 4444 1642 4500
rect 1444 4302 1500 4358
rect 1586 4302 1642 4358
rect 1444 4160 1500 4216
rect 1586 4160 1642 4216
rect 1444 4018 1500 4074
rect 1586 4018 1642 4074
rect 1444 3876 1500 3932
rect 1586 3876 1642 3932
rect 1444 3734 1500 3790
rect 1586 3734 1642 3790
rect 1444 3592 1500 3648
rect 1586 3592 1642 3648
rect 1444 3450 1500 3506
rect 1586 3450 1642 3506
rect 1444 3308 1500 3364
rect 1586 3308 1642 3364
rect 1444 3166 1500 3222
rect 1586 3166 1642 3222
rect 1444 3024 1500 3080
rect 1586 3024 1642 3080
rect 1444 2882 1500 2938
rect 1586 2882 1642 2938
rect 1444 2740 1500 2796
rect 1586 2740 1642 2796
rect 1444 2598 1500 2654
rect 1586 2598 1642 2654
rect 1444 2456 1500 2512
rect 1586 2456 1642 2512
rect 1444 2314 1500 2370
rect 1586 2314 1642 2370
rect 1444 2172 1500 2228
rect 1586 2172 1642 2228
rect 1444 2030 1500 2086
rect 1586 2030 1642 2086
rect 1444 1888 1500 1944
rect 1586 1888 1642 1944
rect 1444 1746 1500 1802
rect 1586 1746 1642 1802
rect 1444 1604 1500 1660
rect 1586 1604 1642 1660
rect 1444 1462 1500 1518
rect 1586 1462 1642 1518
rect 1444 1320 1500 1376
rect 1586 1320 1642 1376
rect 1444 1178 1500 1234
rect 1586 1178 1642 1234
rect 1444 1036 1500 1092
rect 1586 1036 1642 1092
rect 1444 894 1500 950
rect 1586 894 1642 950
rect 1444 752 1500 808
rect 1586 752 1642 808
rect 1444 610 1500 666
rect 1586 610 1642 666
rect 1444 468 1500 524
rect 1586 468 1642 524
rect 1984 12254 2040 12310
rect 2126 12254 2182 12310
rect 1984 12112 2040 12168
rect 2126 12112 2182 12168
rect 1984 11970 2040 12026
rect 2126 11970 2182 12026
rect 1984 11828 2040 11884
rect 2126 11828 2182 11884
rect 1984 11686 2040 11742
rect 2126 11686 2182 11742
rect 1984 11544 2040 11600
rect 2126 11544 2182 11600
rect 1984 11402 2040 11458
rect 2126 11402 2182 11458
rect 1984 11260 2040 11316
rect 2126 11260 2182 11316
rect 1984 11118 2040 11174
rect 2126 11118 2182 11174
rect 1984 10976 2040 11032
rect 2126 10976 2182 11032
rect 1984 10834 2040 10890
rect 2126 10834 2182 10890
rect 1984 10692 2040 10748
rect 2126 10692 2182 10748
rect 1984 10550 2040 10606
rect 2126 10550 2182 10606
rect 1984 10408 2040 10464
rect 2126 10408 2182 10464
rect 1984 10266 2040 10322
rect 2126 10266 2182 10322
rect 1984 10124 2040 10180
rect 2126 10124 2182 10180
rect 1984 9982 2040 10038
rect 2126 9982 2182 10038
rect 1984 9840 2040 9896
rect 2126 9840 2182 9896
rect 1984 9698 2040 9754
rect 2126 9698 2182 9754
rect 1984 9556 2040 9612
rect 2126 9556 2182 9612
rect 1984 9414 2040 9470
rect 2126 9414 2182 9470
rect 1984 9272 2040 9328
rect 2126 9272 2182 9328
rect 1984 9130 2040 9186
rect 2126 9130 2182 9186
rect 1984 8988 2040 9044
rect 2126 8988 2182 9044
rect 1984 8846 2040 8902
rect 2126 8846 2182 8902
rect 1984 8704 2040 8760
rect 2126 8704 2182 8760
rect 1984 8562 2040 8618
rect 2126 8562 2182 8618
rect 1984 8420 2040 8476
rect 2126 8420 2182 8476
rect 1984 8278 2040 8334
rect 2126 8278 2182 8334
rect 1984 8136 2040 8192
rect 2126 8136 2182 8192
rect 1984 7994 2040 8050
rect 2126 7994 2182 8050
rect 1984 7852 2040 7908
rect 2126 7852 2182 7908
rect 1984 7710 2040 7766
rect 2126 7710 2182 7766
rect 1984 7568 2040 7624
rect 2126 7568 2182 7624
rect 1984 7426 2040 7482
rect 2126 7426 2182 7482
rect 1984 7284 2040 7340
rect 2126 7284 2182 7340
rect 1984 7142 2040 7198
rect 2126 7142 2182 7198
rect 1984 7000 2040 7056
rect 2126 7000 2182 7056
rect 1984 6858 2040 6914
rect 2126 6858 2182 6914
rect 1984 6716 2040 6772
rect 2126 6716 2182 6772
rect 1984 6574 2040 6630
rect 2126 6574 2182 6630
rect 1984 6432 2040 6488
rect 2126 6432 2182 6488
rect 1984 6290 2040 6346
rect 2126 6290 2182 6346
rect 1984 6148 2040 6204
rect 2126 6148 2182 6204
rect 1984 6006 2040 6062
rect 2126 6006 2182 6062
rect 1984 5864 2040 5920
rect 2126 5864 2182 5920
rect 1984 5722 2040 5778
rect 2126 5722 2182 5778
rect 1984 5580 2040 5636
rect 2126 5580 2182 5636
rect 1984 5438 2040 5494
rect 2126 5438 2182 5494
rect 1984 5296 2040 5352
rect 2126 5296 2182 5352
rect 1984 5154 2040 5210
rect 2126 5154 2182 5210
rect 1984 5012 2040 5068
rect 2126 5012 2182 5068
rect 1984 4870 2040 4926
rect 2126 4870 2182 4926
rect 1984 4728 2040 4784
rect 2126 4728 2182 4784
rect 1984 4586 2040 4642
rect 2126 4586 2182 4642
rect 1984 4444 2040 4500
rect 2126 4444 2182 4500
rect 1984 4302 2040 4358
rect 2126 4302 2182 4358
rect 1984 4160 2040 4216
rect 2126 4160 2182 4216
rect 1984 4018 2040 4074
rect 2126 4018 2182 4074
rect 1984 3876 2040 3932
rect 2126 3876 2182 3932
rect 1984 3734 2040 3790
rect 2126 3734 2182 3790
rect 1984 3592 2040 3648
rect 2126 3592 2182 3648
rect 1984 3450 2040 3506
rect 2126 3450 2182 3506
rect 1984 3308 2040 3364
rect 2126 3308 2182 3364
rect 1984 3166 2040 3222
rect 2126 3166 2182 3222
rect 1984 3024 2040 3080
rect 2126 3024 2182 3080
rect 1984 2882 2040 2938
rect 2126 2882 2182 2938
rect 1984 2740 2040 2796
rect 2126 2740 2182 2796
rect 1984 2598 2040 2654
rect 2126 2598 2182 2654
rect 1984 2456 2040 2512
rect 2126 2456 2182 2512
rect 1984 2314 2040 2370
rect 2126 2314 2182 2370
rect 1984 2172 2040 2228
rect 2126 2172 2182 2228
rect 1984 2030 2040 2086
rect 2126 2030 2182 2086
rect 1984 1888 2040 1944
rect 2126 1888 2182 1944
rect 1984 1746 2040 1802
rect 2126 1746 2182 1802
rect 1984 1604 2040 1660
rect 2126 1604 2182 1660
rect 1984 1462 2040 1518
rect 2126 1462 2182 1518
rect 1984 1320 2040 1376
rect 2126 1320 2182 1376
rect 1984 1178 2040 1234
rect 2126 1178 2182 1234
rect 1984 1036 2040 1092
rect 2126 1036 2182 1092
rect 1984 894 2040 950
rect 2126 894 2182 950
rect 1984 752 2040 808
rect 2126 752 2182 808
rect 1984 610 2040 666
rect 2126 610 2182 666
rect 1984 468 2040 524
rect 2126 468 2182 524
rect 2521 12254 2577 12310
rect 2663 12254 2719 12310
rect 2521 12112 2577 12168
rect 2663 12112 2719 12168
rect 2521 11970 2577 12026
rect 2663 11970 2719 12026
rect 2521 11828 2577 11884
rect 2663 11828 2719 11884
rect 2521 11686 2577 11742
rect 2663 11686 2719 11742
rect 2521 11544 2577 11600
rect 2663 11544 2719 11600
rect 2521 11402 2577 11458
rect 2663 11402 2719 11458
rect 2521 11260 2577 11316
rect 2663 11260 2719 11316
rect 2521 11118 2577 11174
rect 2663 11118 2719 11174
rect 2521 10976 2577 11032
rect 2663 10976 2719 11032
rect 2521 10834 2577 10890
rect 2663 10834 2719 10890
rect 2521 10692 2577 10748
rect 2663 10692 2719 10748
rect 2521 10550 2577 10606
rect 2663 10550 2719 10606
rect 2521 10408 2577 10464
rect 2663 10408 2719 10464
rect 2521 10266 2577 10322
rect 2663 10266 2719 10322
rect 2521 10124 2577 10180
rect 2663 10124 2719 10180
rect 2521 9982 2577 10038
rect 2663 9982 2719 10038
rect 2521 9840 2577 9896
rect 2663 9840 2719 9896
rect 2521 9698 2577 9754
rect 2663 9698 2719 9754
rect 2521 9556 2577 9612
rect 2663 9556 2719 9612
rect 2521 9414 2577 9470
rect 2663 9414 2719 9470
rect 2521 9272 2577 9328
rect 2663 9272 2719 9328
rect 2521 9130 2577 9186
rect 2663 9130 2719 9186
rect 2521 8988 2577 9044
rect 2663 8988 2719 9044
rect 2521 8846 2577 8902
rect 2663 8846 2719 8902
rect 2521 8704 2577 8760
rect 2663 8704 2719 8760
rect 2521 8562 2577 8618
rect 2663 8562 2719 8618
rect 2521 8420 2577 8476
rect 2663 8420 2719 8476
rect 2521 8278 2577 8334
rect 2663 8278 2719 8334
rect 2521 8136 2577 8192
rect 2663 8136 2719 8192
rect 2521 7994 2577 8050
rect 2663 7994 2719 8050
rect 2521 7852 2577 7908
rect 2663 7852 2719 7908
rect 2521 7710 2577 7766
rect 2663 7710 2719 7766
rect 2521 7568 2577 7624
rect 2663 7568 2719 7624
rect 2521 7426 2577 7482
rect 2663 7426 2719 7482
rect 2521 7284 2577 7340
rect 2663 7284 2719 7340
rect 2521 7142 2577 7198
rect 2663 7142 2719 7198
rect 2521 7000 2577 7056
rect 2663 7000 2719 7056
rect 2521 6858 2577 6914
rect 2663 6858 2719 6914
rect 2521 6716 2577 6772
rect 2663 6716 2719 6772
rect 2521 6574 2577 6630
rect 2663 6574 2719 6630
rect 2521 6432 2577 6488
rect 2663 6432 2719 6488
rect 2521 6290 2577 6346
rect 2663 6290 2719 6346
rect 2521 6148 2577 6204
rect 2663 6148 2719 6204
rect 2521 6006 2577 6062
rect 2663 6006 2719 6062
rect 2521 5864 2577 5920
rect 2663 5864 2719 5920
rect 2521 5722 2577 5778
rect 2663 5722 2719 5778
rect 2521 5580 2577 5636
rect 2663 5580 2719 5636
rect 2521 5438 2577 5494
rect 2663 5438 2719 5494
rect 2521 5296 2577 5352
rect 2663 5296 2719 5352
rect 2521 5154 2577 5210
rect 2663 5154 2719 5210
rect 2521 5012 2577 5068
rect 2663 5012 2719 5068
rect 2521 4870 2577 4926
rect 2663 4870 2719 4926
rect 2521 4728 2577 4784
rect 2663 4728 2719 4784
rect 2521 4586 2577 4642
rect 2663 4586 2719 4642
rect 2521 4444 2577 4500
rect 2663 4444 2719 4500
rect 2521 4302 2577 4358
rect 2663 4302 2719 4358
rect 2521 4160 2577 4216
rect 2663 4160 2719 4216
rect 2521 4018 2577 4074
rect 2663 4018 2719 4074
rect 2521 3876 2577 3932
rect 2663 3876 2719 3932
rect 2521 3734 2577 3790
rect 2663 3734 2719 3790
rect 2521 3592 2577 3648
rect 2663 3592 2719 3648
rect 2521 3450 2577 3506
rect 2663 3450 2719 3506
rect 2521 3308 2577 3364
rect 2663 3308 2719 3364
rect 2521 3166 2577 3222
rect 2663 3166 2719 3222
rect 2521 3024 2577 3080
rect 2663 3024 2719 3080
rect 2521 2882 2577 2938
rect 2663 2882 2719 2938
rect 2521 2740 2577 2796
rect 2663 2740 2719 2796
rect 2521 2598 2577 2654
rect 2663 2598 2719 2654
rect 2521 2456 2577 2512
rect 2663 2456 2719 2512
rect 2521 2314 2577 2370
rect 2663 2314 2719 2370
rect 2521 2172 2577 2228
rect 2663 2172 2719 2228
rect 2521 2030 2577 2086
rect 2663 2030 2719 2086
rect 2521 1888 2577 1944
rect 2663 1888 2719 1944
rect 2521 1746 2577 1802
rect 2663 1746 2719 1802
rect 2521 1604 2577 1660
rect 2663 1604 2719 1660
rect 2521 1462 2577 1518
rect 2663 1462 2719 1518
rect 2521 1320 2577 1376
rect 2663 1320 2719 1376
rect 2521 1178 2577 1234
rect 2663 1178 2719 1234
rect 2521 1036 2577 1092
rect 2663 1036 2719 1092
rect 2521 894 2577 950
rect 2663 894 2719 950
rect 2521 752 2577 808
rect 2663 752 2719 808
rect 2521 610 2577 666
rect 2663 610 2719 666
rect 2521 468 2577 524
rect 2663 468 2719 524
rect 3058 12254 3114 12310
rect 3200 12254 3256 12310
rect 3058 12112 3114 12168
rect 3200 12112 3256 12168
rect 3058 11970 3114 12026
rect 3200 11970 3256 12026
rect 3058 11828 3114 11884
rect 3200 11828 3256 11884
rect 3058 11686 3114 11742
rect 3200 11686 3256 11742
rect 3058 11544 3114 11600
rect 3200 11544 3256 11600
rect 3058 11402 3114 11458
rect 3200 11402 3256 11458
rect 3058 11260 3114 11316
rect 3200 11260 3256 11316
rect 3058 11118 3114 11174
rect 3200 11118 3256 11174
rect 3058 10976 3114 11032
rect 3200 10976 3256 11032
rect 3058 10834 3114 10890
rect 3200 10834 3256 10890
rect 3058 10692 3114 10748
rect 3200 10692 3256 10748
rect 3058 10550 3114 10606
rect 3200 10550 3256 10606
rect 3058 10408 3114 10464
rect 3200 10408 3256 10464
rect 3058 10266 3114 10322
rect 3200 10266 3256 10322
rect 3058 10124 3114 10180
rect 3200 10124 3256 10180
rect 3058 9982 3114 10038
rect 3200 9982 3256 10038
rect 3058 9840 3114 9896
rect 3200 9840 3256 9896
rect 3058 9698 3114 9754
rect 3200 9698 3256 9754
rect 3058 9556 3114 9612
rect 3200 9556 3256 9612
rect 3058 9414 3114 9470
rect 3200 9414 3256 9470
rect 3058 9272 3114 9328
rect 3200 9272 3256 9328
rect 3058 9130 3114 9186
rect 3200 9130 3256 9186
rect 3058 8988 3114 9044
rect 3200 8988 3256 9044
rect 3058 8846 3114 8902
rect 3200 8846 3256 8902
rect 3058 8704 3114 8760
rect 3200 8704 3256 8760
rect 3058 8562 3114 8618
rect 3200 8562 3256 8618
rect 3058 8420 3114 8476
rect 3200 8420 3256 8476
rect 3058 8278 3114 8334
rect 3200 8278 3256 8334
rect 3058 8136 3114 8192
rect 3200 8136 3256 8192
rect 3058 7994 3114 8050
rect 3200 7994 3256 8050
rect 3058 7852 3114 7908
rect 3200 7852 3256 7908
rect 3058 7710 3114 7766
rect 3200 7710 3256 7766
rect 3058 7568 3114 7624
rect 3200 7568 3256 7624
rect 3058 7426 3114 7482
rect 3200 7426 3256 7482
rect 3058 7284 3114 7340
rect 3200 7284 3256 7340
rect 3058 7142 3114 7198
rect 3200 7142 3256 7198
rect 3058 7000 3114 7056
rect 3200 7000 3256 7056
rect 3058 6858 3114 6914
rect 3200 6858 3256 6914
rect 3058 6716 3114 6772
rect 3200 6716 3256 6772
rect 3058 6574 3114 6630
rect 3200 6574 3256 6630
rect 3058 6432 3114 6488
rect 3200 6432 3256 6488
rect 3058 6290 3114 6346
rect 3200 6290 3256 6346
rect 3058 6148 3114 6204
rect 3200 6148 3256 6204
rect 3058 6006 3114 6062
rect 3200 6006 3256 6062
rect 3058 5864 3114 5920
rect 3200 5864 3256 5920
rect 3058 5722 3114 5778
rect 3200 5722 3256 5778
rect 3058 5580 3114 5636
rect 3200 5580 3256 5636
rect 3058 5438 3114 5494
rect 3200 5438 3256 5494
rect 3058 5296 3114 5352
rect 3200 5296 3256 5352
rect 3058 5154 3114 5210
rect 3200 5154 3256 5210
rect 3058 5012 3114 5068
rect 3200 5012 3256 5068
rect 3058 4870 3114 4926
rect 3200 4870 3256 4926
rect 3058 4728 3114 4784
rect 3200 4728 3256 4784
rect 3058 4586 3114 4642
rect 3200 4586 3256 4642
rect 3058 4444 3114 4500
rect 3200 4444 3256 4500
rect 3058 4302 3114 4358
rect 3200 4302 3256 4358
rect 3058 4160 3114 4216
rect 3200 4160 3256 4216
rect 3058 4018 3114 4074
rect 3200 4018 3256 4074
rect 3058 3876 3114 3932
rect 3200 3876 3256 3932
rect 3058 3734 3114 3790
rect 3200 3734 3256 3790
rect 3058 3592 3114 3648
rect 3200 3592 3256 3648
rect 3058 3450 3114 3506
rect 3200 3450 3256 3506
rect 3058 3308 3114 3364
rect 3200 3308 3256 3364
rect 3058 3166 3114 3222
rect 3200 3166 3256 3222
rect 3058 3024 3114 3080
rect 3200 3024 3256 3080
rect 3058 2882 3114 2938
rect 3200 2882 3256 2938
rect 3058 2740 3114 2796
rect 3200 2740 3256 2796
rect 3058 2598 3114 2654
rect 3200 2598 3256 2654
rect 3058 2456 3114 2512
rect 3200 2456 3256 2512
rect 3058 2314 3114 2370
rect 3200 2314 3256 2370
rect 3058 2172 3114 2228
rect 3200 2172 3256 2228
rect 3058 2030 3114 2086
rect 3200 2030 3256 2086
rect 3058 1888 3114 1944
rect 3200 1888 3256 1944
rect 3058 1746 3114 1802
rect 3200 1746 3256 1802
rect 3058 1604 3114 1660
rect 3200 1604 3256 1660
rect 3058 1462 3114 1518
rect 3200 1462 3256 1518
rect 3058 1320 3114 1376
rect 3200 1320 3256 1376
rect 3058 1178 3114 1234
rect 3200 1178 3256 1234
rect 3058 1036 3114 1092
rect 3200 1036 3256 1092
rect 3058 894 3114 950
rect 3200 894 3256 950
rect 3058 752 3114 808
rect 3200 752 3256 808
rect 3058 610 3114 666
rect 3200 610 3256 666
rect 3058 468 3114 524
rect 3200 468 3256 524
rect 3602 12254 3658 12310
rect 3744 12254 3800 12310
rect 3602 12112 3658 12168
rect 3744 12112 3800 12168
rect 3602 11970 3658 12026
rect 3744 11970 3800 12026
rect 3602 11828 3658 11884
rect 3744 11828 3800 11884
rect 3602 11686 3658 11742
rect 3744 11686 3800 11742
rect 3602 11544 3658 11600
rect 3744 11544 3800 11600
rect 3602 11402 3658 11458
rect 3744 11402 3800 11458
rect 3602 11260 3658 11316
rect 3744 11260 3800 11316
rect 3602 11118 3658 11174
rect 3744 11118 3800 11174
rect 3602 10976 3658 11032
rect 3744 10976 3800 11032
rect 3602 10834 3658 10890
rect 3744 10834 3800 10890
rect 3602 10692 3658 10748
rect 3744 10692 3800 10748
rect 3602 10550 3658 10606
rect 3744 10550 3800 10606
rect 3602 10408 3658 10464
rect 3744 10408 3800 10464
rect 3602 10266 3658 10322
rect 3744 10266 3800 10322
rect 3602 10124 3658 10180
rect 3744 10124 3800 10180
rect 3602 9982 3658 10038
rect 3744 9982 3800 10038
rect 3602 9840 3658 9896
rect 3744 9840 3800 9896
rect 3602 9698 3658 9754
rect 3744 9698 3800 9754
rect 3602 9556 3658 9612
rect 3744 9556 3800 9612
rect 3602 9414 3658 9470
rect 3744 9414 3800 9470
rect 3602 9272 3658 9328
rect 3744 9272 3800 9328
rect 3602 9130 3658 9186
rect 3744 9130 3800 9186
rect 3602 8988 3658 9044
rect 3744 8988 3800 9044
rect 3602 8846 3658 8902
rect 3744 8846 3800 8902
rect 3602 8704 3658 8760
rect 3744 8704 3800 8760
rect 3602 8562 3658 8618
rect 3744 8562 3800 8618
rect 3602 8420 3658 8476
rect 3744 8420 3800 8476
rect 3602 8278 3658 8334
rect 3744 8278 3800 8334
rect 3602 8136 3658 8192
rect 3744 8136 3800 8192
rect 3602 7994 3658 8050
rect 3744 7994 3800 8050
rect 3602 7852 3658 7908
rect 3744 7852 3800 7908
rect 3602 7710 3658 7766
rect 3744 7710 3800 7766
rect 3602 7568 3658 7624
rect 3744 7568 3800 7624
rect 3602 7426 3658 7482
rect 3744 7426 3800 7482
rect 3602 7284 3658 7340
rect 3744 7284 3800 7340
rect 3602 7142 3658 7198
rect 3744 7142 3800 7198
rect 3602 7000 3658 7056
rect 3744 7000 3800 7056
rect 3602 6858 3658 6914
rect 3744 6858 3800 6914
rect 3602 6716 3658 6772
rect 3744 6716 3800 6772
rect 3602 6574 3658 6630
rect 3744 6574 3800 6630
rect 3602 6432 3658 6488
rect 3744 6432 3800 6488
rect 3602 6290 3658 6346
rect 3744 6290 3800 6346
rect 3602 6148 3658 6204
rect 3744 6148 3800 6204
rect 3602 6006 3658 6062
rect 3744 6006 3800 6062
rect 3602 5864 3658 5920
rect 3744 5864 3800 5920
rect 3602 5722 3658 5778
rect 3744 5722 3800 5778
rect 3602 5580 3658 5636
rect 3744 5580 3800 5636
rect 3602 5438 3658 5494
rect 3744 5438 3800 5494
rect 3602 5296 3658 5352
rect 3744 5296 3800 5352
rect 3602 5154 3658 5210
rect 3744 5154 3800 5210
rect 3602 5012 3658 5068
rect 3744 5012 3800 5068
rect 3602 4870 3658 4926
rect 3744 4870 3800 4926
rect 3602 4728 3658 4784
rect 3744 4728 3800 4784
rect 3602 4586 3658 4642
rect 3744 4586 3800 4642
rect 3602 4444 3658 4500
rect 3744 4444 3800 4500
rect 3602 4302 3658 4358
rect 3744 4302 3800 4358
rect 3602 4160 3658 4216
rect 3744 4160 3800 4216
rect 3602 4018 3658 4074
rect 3744 4018 3800 4074
rect 3602 3876 3658 3932
rect 3744 3876 3800 3932
rect 3602 3734 3658 3790
rect 3744 3734 3800 3790
rect 3602 3592 3658 3648
rect 3744 3592 3800 3648
rect 3602 3450 3658 3506
rect 3744 3450 3800 3506
rect 3602 3308 3658 3364
rect 3744 3308 3800 3364
rect 3602 3166 3658 3222
rect 3744 3166 3800 3222
rect 3602 3024 3658 3080
rect 3744 3024 3800 3080
rect 3602 2882 3658 2938
rect 3744 2882 3800 2938
rect 3602 2740 3658 2796
rect 3744 2740 3800 2796
rect 3602 2598 3658 2654
rect 3744 2598 3800 2654
rect 3602 2456 3658 2512
rect 3744 2456 3800 2512
rect 3602 2314 3658 2370
rect 3744 2314 3800 2370
rect 3602 2172 3658 2228
rect 3744 2172 3800 2228
rect 3602 2030 3658 2086
rect 3744 2030 3800 2086
rect 3602 1888 3658 1944
rect 3744 1888 3800 1944
rect 3602 1746 3658 1802
rect 3744 1746 3800 1802
rect 3602 1604 3658 1660
rect 3744 1604 3800 1660
rect 3602 1462 3658 1518
rect 3744 1462 3800 1518
rect 3602 1320 3658 1376
rect 3744 1320 3800 1376
rect 3602 1178 3658 1234
rect 3744 1178 3800 1234
rect 3602 1036 3658 1092
rect 3744 1036 3800 1092
rect 3602 894 3658 950
rect 3744 894 3800 950
rect 3602 752 3658 808
rect 3744 752 3800 808
rect 3602 610 3658 666
rect 3744 610 3800 666
rect 3602 468 3658 524
rect 3744 468 3800 524
rect 4138 12254 4194 12310
rect 4280 12254 4336 12310
rect 4138 12112 4194 12168
rect 4280 12112 4336 12168
rect 4138 11970 4194 12026
rect 4280 11970 4336 12026
rect 4138 11828 4194 11884
rect 4280 11828 4336 11884
rect 4138 11686 4194 11742
rect 4280 11686 4336 11742
rect 4138 11544 4194 11600
rect 4280 11544 4336 11600
rect 4138 11402 4194 11458
rect 4280 11402 4336 11458
rect 4138 11260 4194 11316
rect 4280 11260 4336 11316
rect 4138 11118 4194 11174
rect 4280 11118 4336 11174
rect 4138 10976 4194 11032
rect 4280 10976 4336 11032
rect 4138 10834 4194 10890
rect 4280 10834 4336 10890
rect 4138 10692 4194 10748
rect 4280 10692 4336 10748
rect 4138 10550 4194 10606
rect 4280 10550 4336 10606
rect 4138 10408 4194 10464
rect 4280 10408 4336 10464
rect 4138 10266 4194 10322
rect 4280 10266 4336 10322
rect 4138 10124 4194 10180
rect 4280 10124 4336 10180
rect 4138 9982 4194 10038
rect 4280 9982 4336 10038
rect 4138 9840 4194 9896
rect 4280 9840 4336 9896
rect 4138 9698 4194 9754
rect 4280 9698 4336 9754
rect 4138 9556 4194 9612
rect 4280 9556 4336 9612
rect 4138 9414 4194 9470
rect 4280 9414 4336 9470
rect 4138 9272 4194 9328
rect 4280 9272 4336 9328
rect 4138 9130 4194 9186
rect 4280 9130 4336 9186
rect 4138 8988 4194 9044
rect 4280 8988 4336 9044
rect 4138 8846 4194 8902
rect 4280 8846 4336 8902
rect 4138 8704 4194 8760
rect 4280 8704 4336 8760
rect 4138 8562 4194 8618
rect 4280 8562 4336 8618
rect 4138 8420 4194 8476
rect 4280 8420 4336 8476
rect 4138 8278 4194 8334
rect 4280 8278 4336 8334
rect 4138 8136 4194 8192
rect 4280 8136 4336 8192
rect 4138 7994 4194 8050
rect 4280 7994 4336 8050
rect 4138 7852 4194 7908
rect 4280 7852 4336 7908
rect 4138 7710 4194 7766
rect 4280 7710 4336 7766
rect 4138 7568 4194 7624
rect 4280 7568 4336 7624
rect 4138 7426 4194 7482
rect 4280 7426 4336 7482
rect 4138 7284 4194 7340
rect 4280 7284 4336 7340
rect 4138 7142 4194 7198
rect 4280 7142 4336 7198
rect 4138 7000 4194 7056
rect 4280 7000 4336 7056
rect 4138 6858 4194 6914
rect 4280 6858 4336 6914
rect 4138 6716 4194 6772
rect 4280 6716 4336 6772
rect 4138 6574 4194 6630
rect 4280 6574 4336 6630
rect 4138 6432 4194 6488
rect 4280 6432 4336 6488
rect 4138 6290 4194 6346
rect 4280 6290 4336 6346
rect 4138 6148 4194 6204
rect 4280 6148 4336 6204
rect 4138 6006 4194 6062
rect 4280 6006 4336 6062
rect 4138 5864 4194 5920
rect 4280 5864 4336 5920
rect 4138 5722 4194 5778
rect 4280 5722 4336 5778
rect 4138 5580 4194 5636
rect 4280 5580 4336 5636
rect 4138 5438 4194 5494
rect 4280 5438 4336 5494
rect 4138 5296 4194 5352
rect 4280 5296 4336 5352
rect 4138 5154 4194 5210
rect 4280 5154 4336 5210
rect 4138 5012 4194 5068
rect 4280 5012 4336 5068
rect 4138 4870 4194 4926
rect 4280 4870 4336 4926
rect 4138 4728 4194 4784
rect 4280 4728 4336 4784
rect 4138 4586 4194 4642
rect 4280 4586 4336 4642
rect 4138 4444 4194 4500
rect 4280 4444 4336 4500
rect 4138 4302 4194 4358
rect 4280 4302 4336 4358
rect 4138 4160 4194 4216
rect 4280 4160 4336 4216
rect 4138 4018 4194 4074
rect 4280 4018 4336 4074
rect 4138 3876 4194 3932
rect 4280 3876 4336 3932
rect 4138 3734 4194 3790
rect 4280 3734 4336 3790
rect 4138 3592 4194 3648
rect 4280 3592 4336 3648
rect 4138 3450 4194 3506
rect 4280 3450 4336 3506
rect 4138 3308 4194 3364
rect 4280 3308 4336 3364
rect 4138 3166 4194 3222
rect 4280 3166 4336 3222
rect 4138 3024 4194 3080
rect 4280 3024 4336 3080
rect 4138 2882 4194 2938
rect 4280 2882 4336 2938
rect 4138 2740 4194 2796
rect 4280 2740 4336 2796
rect 4138 2598 4194 2654
rect 4280 2598 4336 2654
rect 4138 2456 4194 2512
rect 4280 2456 4336 2512
rect 4138 2314 4194 2370
rect 4280 2314 4336 2370
rect 4138 2172 4194 2228
rect 4280 2172 4336 2228
rect 4138 2030 4194 2086
rect 4280 2030 4336 2086
rect 4138 1888 4194 1944
rect 4280 1888 4336 1944
rect 4138 1746 4194 1802
rect 4280 1746 4336 1802
rect 4138 1604 4194 1660
rect 4280 1604 4336 1660
rect 4138 1462 4194 1518
rect 4280 1462 4336 1518
rect 4138 1320 4194 1376
rect 4280 1320 4336 1376
rect 4138 1178 4194 1234
rect 4280 1178 4336 1234
rect 4138 1036 4194 1092
rect 4280 1036 4336 1092
rect 4138 894 4194 950
rect 4280 894 4336 950
rect 4138 752 4194 808
rect 4280 752 4336 808
rect 4138 610 4194 666
rect 4280 610 4336 666
rect 4138 468 4194 524
rect 4280 468 4336 524
rect 4678 12254 4734 12310
rect 4820 12254 4876 12310
rect 4678 12112 4734 12168
rect 4820 12112 4876 12168
rect 4678 11970 4734 12026
rect 4820 11970 4876 12026
rect 4678 11828 4734 11884
rect 4820 11828 4876 11884
rect 4678 11686 4734 11742
rect 4820 11686 4876 11742
rect 4678 11544 4734 11600
rect 4820 11544 4876 11600
rect 4678 11402 4734 11458
rect 4820 11402 4876 11458
rect 4678 11260 4734 11316
rect 4820 11260 4876 11316
rect 4678 11118 4734 11174
rect 4820 11118 4876 11174
rect 4678 10976 4734 11032
rect 4820 10976 4876 11032
rect 4678 10834 4734 10890
rect 4820 10834 4876 10890
rect 4678 10692 4734 10748
rect 4820 10692 4876 10748
rect 4678 10550 4734 10606
rect 4820 10550 4876 10606
rect 4678 10408 4734 10464
rect 4820 10408 4876 10464
rect 4678 10266 4734 10322
rect 4820 10266 4876 10322
rect 4678 10124 4734 10180
rect 4820 10124 4876 10180
rect 4678 9982 4734 10038
rect 4820 9982 4876 10038
rect 4678 9840 4734 9896
rect 4820 9840 4876 9896
rect 4678 9698 4734 9754
rect 4820 9698 4876 9754
rect 4678 9556 4734 9612
rect 4820 9556 4876 9612
rect 4678 9414 4734 9470
rect 4820 9414 4876 9470
rect 4678 9272 4734 9328
rect 4820 9272 4876 9328
rect 4678 9130 4734 9186
rect 4820 9130 4876 9186
rect 4678 8988 4734 9044
rect 4820 8988 4876 9044
rect 4678 8846 4734 8902
rect 4820 8846 4876 8902
rect 4678 8704 4734 8760
rect 4820 8704 4876 8760
rect 4678 8562 4734 8618
rect 4820 8562 4876 8618
rect 4678 8420 4734 8476
rect 4820 8420 4876 8476
rect 4678 8278 4734 8334
rect 4820 8278 4876 8334
rect 4678 8136 4734 8192
rect 4820 8136 4876 8192
rect 4678 7994 4734 8050
rect 4820 7994 4876 8050
rect 4678 7852 4734 7908
rect 4820 7852 4876 7908
rect 4678 7710 4734 7766
rect 4820 7710 4876 7766
rect 4678 7568 4734 7624
rect 4820 7568 4876 7624
rect 4678 7426 4734 7482
rect 4820 7426 4876 7482
rect 4678 7284 4734 7340
rect 4820 7284 4876 7340
rect 4678 7142 4734 7198
rect 4820 7142 4876 7198
rect 4678 7000 4734 7056
rect 4820 7000 4876 7056
rect 4678 6858 4734 6914
rect 4820 6858 4876 6914
rect 4678 6716 4734 6772
rect 4820 6716 4876 6772
rect 4678 6574 4734 6630
rect 4820 6574 4876 6630
rect 4678 6432 4734 6488
rect 4820 6432 4876 6488
rect 4678 6290 4734 6346
rect 4820 6290 4876 6346
rect 4678 6148 4734 6204
rect 4820 6148 4876 6204
rect 4678 6006 4734 6062
rect 4820 6006 4876 6062
rect 4678 5864 4734 5920
rect 4820 5864 4876 5920
rect 4678 5722 4734 5778
rect 4820 5722 4876 5778
rect 4678 5580 4734 5636
rect 4820 5580 4876 5636
rect 4678 5438 4734 5494
rect 4820 5438 4876 5494
rect 4678 5296 4734 5352
rect 4820 5296 4876 5352
rect 4678 5154 4734 5210
rect 4820 5154 4876 5210
rect 4678 5012 4734 5068
rect 4820 5012 4876 5068
rect 4678 4870 4734 4926
rect 4820 4870 4876 4926
rect 4678 4728 4734 4784
rect 4820 4728 4876 4784
rect 4678 4586 4734 4642
rect 4820 4586 4876 4642
rect 4678 4444 4734 4500
rect 4820 4444 4876 4500
rect 4678 4302 4734 4358
rect 4820 4302 4876 4358
rect 4678 4160 4734 4216
rect 4820 4160 4876 4216
rect 4678 4018 4734 4074
rect 4820 4018 4876 4074
rect 4678 3876 4734 3932
rect 4820 3876 4876 3932
rect 4678 3734 4734 3790
rect 4820 3734 4876 3790
rect 4678 3592 4734 3648
rect 4820 3592 4876 3648
rect 4678 3450 4734 3506
rect 4820 3450 4876 3506
rect 4678 3308 4734 3364
rect 4820 3308 4876 3364
rect 4678 3166 4734 3222
rect 4820 3166 4876 3222
rect 4678 3024 4734 3080
rect 4820 3024 4876 3080
rect 4678 2882 4734 2938
rect 4820 2882 4876 2938
rect 4678 2740 4734 2796
rect 4820 2740 4876 2796
rect 4678 2598 4734 2654
rect 4820 2598 4876 2654
rect 4678 2456 4734 2512
rect 4820 2456 4876 2512
rect 4678 2314 4734 2370
rect 4820 2314 4876 2370
rect 4678 2172 4734 2228
rect 4820 2172 4876 2228
rect 4678 2030 4734 2086
rect 4820 2030 4876 2086
rect 4678 1888 4734 1944
rect 4820 1888 4876 1944
rect 4678 1746 4734 1802
rect 4820 1746 4876 1802
rect 4678 1604 4734 1660
rect 4820 1604 4876 1660
rect 4678 1462 4734 1518
rect 4820 1462 4876 1518
rect 4678 1320 4734 1376
rect 4820 1320 4876 1376
rect 4678 1178 4734 1234
rect 4820 1178 4876 1234
rect 4678 1036 4734 1092
rect 4820 1036 4876 1092
rect 4678 894 4734 950
rect 4820 894 4876 950
rect 4678 752 4734 808
rect 4820 752 4876 808
rect 4678 610 4734 666
rect 4820 610 4876 666
rect 4678 468 4734 524
rect 4820 468 4876 524
rect 5215 12254 5271 12310
rect 5357 12254 5413 12310
rect 5215 12112 5271 12168
rect 5357 12112 5413 12168
rect 5215 11970 5271 12026
rect 5357 11970 5413 12026
rect 5215 11828 5271 11884
rect 5357 11828 5413 11884
rect 5215 11686 5271 11742
rect 5357 11686 5413 11742
rect 5215 11544 5271 11600
rect 5357 11544 5413 11600
rect 5215 11402 5271 11458
rect 5357 11402 5413 11458
rect 5215 11260 5271 11316
rect 5357 11260 5413 11316
rect 5215 11118 5271 11174
rect 5357 11118 5413 11174
rect 5215 10976 5271 11032
rect 5357 10976 5413 11032
rect 5215 10834 5271 10890
rect 5357 10834 5413 10890
rect 5215 10692 5271 10748
rect 5357 10692 5413 10748
rect 5215 10550 5271 10606
rect 5357 10550 5413 10606
rect 5215 10408 5271 10464
rect 5357 10408 5413 10464
rect 5215 10266 5271 10322
rect 5357 10266 5413 10322
rect 5215 10124 5271 10180
rect 5357 10124 5413 10180
rect 5215 9982 5271 10038
rect 5357 9982 5413 10038
rect 5215 9840 5271 9896
rect 5357 9840 5413 9896
rect 5215 9698 5271 9754
rect 5357 9698 5413 9754
rect 5215 9556 5271 9612
rect 5357 9556 5413 9612
rect 5215 9414 5271 9470
rect 5357 9414 5413 9470
rect 5215 9272 5271 9328
rect 5357 9272 5413 9328
rect 5215 9130 5271 9186
rect 5357 9130 5413 9186
rect 5215 8988 5271 9044
rect 5357 8988 5413 9044
rect 5215 8846 5271 8902
rect 5357 8846 5413 8902
rect 5215 8704 5271 8760
rect 5357 8704 5413 8760
rect 5215 8562 5271 8618
rect 5357 8562 5413 8618
rect 5215 8420 5271 8476
rect 5357 8420 5413 8476
rect 5215 8278 5271 8334
rect 5357 8278 5413 8334
rect 5215 8136 5271 8192
rect 5357 8136 5413 8192
rect 5215 7994 5271 8050
rect 5357 7994 5413 8050
rect 5215 7852 5271 7908
rect 5357 7852 5413 7908
rect 5215 7710 5271 7766
rect 5357 7710 5413 7766
rect 5215 7568 5271 7624
rect 5357 7568 5413 7624
rect 5215 7426 5271 7482
rect 5357 7426 5413 7482
rect 5215 7284 5271 7340
rect 5357 7284 5413 7340
rect 5215 7142 5271 7198
rect 5357 7142 5413 7198
rect 5215 7000 5271 7056
rect 5357 7000 5413 7056
rect 5215 6858 5271 6914
rect 5357 6858 5413 6914
rect 5215 6716 5271 6772
rect 5357 6716 5413 6772
rect 5215 6574 5271 6630
rect 5357 6574 5413 6630
rect 5215 6432 5271 6488
rect 5357 6432 5413 6488
rect 5215 6290 5271 6346
rect 5357 6290 5413 6346
rect 5215 6148 5271 6204
rect 5357 6148 5413 6204
rect 5215 6006 5271 6062
rect 5357 6006 5413 6062
rect 5215 5864 5271 5920
rect 5357 5864 5413 5920
rect 5215 5722 5271 5778
rect 5357 5722 5413 5778
rect 5215 5580 5271 5636
rect 5357 5580 5413 5636
rect 5215 5438 5271 5494
rect 5357 5438 5413 5494
rect 5215 5296 5271 5352
rect 5357 5296 5413 5352
rect 5215 5154 5271 5210
rect 5357 5154 5413 5210
rect 5215 5012 5271 5068
rect 5357 5012 5413 5068
rect 5215 4870 5271 4926
rect 5357 4870 5413 4926
rect 5215 4728 5271 4784
rect 5357 4728 5413 4784
rect 5215 4586 5271 4642
rect 5357 4586 5413 4642
rect 5215 4444 5271 4500
rect 5357 4444 5413 4500
rect 5215 4302 5271 4358
rect 5357 4302 5413 4358
rect 5215 4160 5271 4216
rect 5357 4160 5413 4216
rect 5215 4018 5271 4074
rect 5357 4018 5413 4074
rect 5215 3876 5271 3932
rect 5357 3876 5413 3932
rect 5215 3734 5271 3790
rect 5357 3734 5413 3790
rect 5215 3592 5271 3648
rect 5357 3592 5413 3648
rect 5215 3450 5271 3506
rect 5357 3450 5413 3506
rect 5215 3308 5271 3364
rect 5357 3308 5413 3364
rect 5215 3166 5271 3222
rect 5357 3166 5413 3222
rect 5215 3024 5271 3080
rect 5357 3024 5413 3080
rect 5215 2882 5271 2938
rect 5357 2882 5413 2938
rect 5215 2740 5271 2796
rect 5357 2740 5413 2796
rect 5215 2598 5271 2654
rect 5357 2598 5413 2654
rect 5215 2456 5271 2512
rect 5357 2456 5413 2512
rect 5215 2314 5271 2370
rect 5357 2314 5413 2370
rect 5215 2172 5271 2228
rect 5357 2172 5413 2228
rect 5215 2030 5271 2086
rect 5357 2030 5413 2086
rect 5215 1888 5271 1944
rect 5357 1888 5413 1944
rect 5215 1746 5271 1802
rect 5357 1746 5413 1802
rect 5215 1604 5271 1660
rect 5357 1604 5413 1660
rect 5215 1462 5271 1518
rect 5357 1462 5413 1518
rect 5215 1320 5271 1376
rect 5357 1320 5413 1376
rect 5215 1178 5271 1234
rect 5357 1178 5413 1234
rect 5215 1036 5271 1092
rect 5357 1036 5413 1092
rect 5215 894 5271 950
rect 5357 894 5413 950
rect 5215 752 5271 808
rect 5357 752 5413 808
rect 5215 610 5271 666
rect 5357 610 5413 666
rect 5215 468 5271 524
rect 5357 468 5413 524
rect 5760 12254 5816 12310
rect 5902 12254 5958 12310
rect 5760 12112 5816 12168
rect 5902 12112 5958 12168
rect 5760 11970 5816 12026
rect 5902 11970 5958 12026
rect 5760 11828 5816 11884
rect 5902 11828 5958 11884
rect 5760 11686 5816 11742
rect 5902 11686 5958 11742
rect 5760 11544 5816 11600
rect 5902 11544 5958 11600
rect 5760 11402 5816 11458
rect 5902 11402 5958 11458
rect 5760 11260 5816 11316
rect 5902 11260 5958 11316
rect 5760 11118 5816 11174
rect 5902 11118 5958 11174
rect 5760 10976 5816 11032
rect 5902 10976 5958 11032
rect 5760 10834 5816 10890
rect 5902 10834 5958 10890
rect 5760 10692 5816 10748
rect 5902 10692 5958 10748
rect 5760 10550 5816 10606
rect 5902 10550 5958 10606
rect 5760 10408 5816 10464
rect 5902 10408 5958 10464
rect 5760 10266 5816 10322
rect 5902 10266 5958 10322
rect 5760 10124 5816 10180
rect 5902 10124 5958 10180
rect 5760 9982 5816 10038
rect 5902 9982 5958 10038
rect 5760 9840 5816 9896
rect 5902 9840 5958 9896
rect 5760 9698 5816 9754
rect 5902 9698 5958 9754
rect 5760 9556 5816 9612
rect 5902 9556 5958 9612
rect 5760 9414 5816 9470
rect 5902 9414 5958 9470
rect 5760 9272 5816 9328
rect 5902 9272 5958 9328
rect 5760 9130 5816 9186
rect 5902 9130 5958 9186
rect 5760 8988 5816 9044
rect 5902 8988 5958 9044
rect 5760 8846 5816 8902
rect 5902 8846 5958 8902
rect 5760 8704 5816 8760
rect 5902 8704 5958 8760
rect 5760 8562 5816 8618
rect 5902 8562 5958 8618
rect 5760 8420 5816 8476
rect 5902 8420 5958 8476
rect 5760 8278 5816 8334
rect 5902 8278 5958 8334
rect 5760 8136 5816 8192
rect 5902 8136 5958 8192
rect 5760 7994 5816 8050
rect 5902 7994 5958 8050
rect 5760 7852 5816 7908
rect 5902 7852 5958 7908
rect 5760 7710 5816 7766
rect 5902 7710 5958 7766
rect 5760 7568 5816 7624
rect 5902 7568 5958 7624
rect 5760 7426 5816 7482
rect 5902 7426 5958 7482
rect 5760 7284 5816 7340
rect 5902 7284 5958 7340
rect 5760 7142 5816 7198
rect 5902 7142 5958 7198
rect 5760 7000 5816 7056
rect 5902 7000 5958 7056
rect 5760 6858 5816 6914
rect 5902 6858 5958 6914
rect 5760 6716 5816 6772
rect 5902 6716 5958 6772
rect 5760 6574 5816 6630
rect 5902 6574 5958 6630
rect 5760 6432 5816 6488
rect 5902 6432 5958 6488
rect 5760 6290 5816 6346
rect 5902 6290 5958 6346
rect 5760 6148 5816 6204
rect 5902 6148 5958 6204
rect 5760 6006 5816 6062
rect 5902 6006 5958 6062
rect 5760 5864 5816 5920
rect 5902 5864 5958 5920
rect 5760 5722 5816 5778
rect 5902 5722 5958 5778
rect 5760 5580 5816 5636
rect 5902 5580 5958 5636
rect 5760 5438 5816 5494
rect 5902 5438 5958 5494
rect 5760 5296 5816 5352
rect 5902 5296 5958 5352
rect 5760 5154 5816 5210
rect 5902 5154 5958 5210
rect 5760 5012 5816 5068
rect 5902 5012 5958 5068
rect 5760 4870 5816 4926
rect 5902 4870 5958 4926
rect 5760 4728 5816 4784
rect 5902 4728 5958 4784
rect 5760 4586 5816 4642
rect 5902 4586 5958 4642
rect 5760 4444 5816 4500
rect 5902 4444 5958 4500
rect 5760 4302 5816 4358
rect 5902 4302 5958 4358
rect 5760 4160 5816 4216
rect 5902 4160 5958 4216
rect 5760 4018 5816 4074
rect 5902 4018 5958 4074
rect 5760 3876 5816 3932
rect 5902 3876 5958 3932
rect 5760 3734 5816 3790
rect 5902 3734 5958 3790
rect 5760 3592 5816 3648
rect 5902 3592 5958 3648
rect 5760 3450 5816 3506
rect 5902 3450 5958 3506
rect 5760 3308 5816 3364
rect 5902 3308 5958 3364
rect 5760 3166 5816 3222
rect 5902 3166 5958 3222
rect 5760 3024 5816 3080
rect 5902 3024 5958 3080
rect 5760 2882 5816 2938
rect 5902 2882 5958 2938
rect 5760 2740 5816 2796
rect 5902 2740 5958 2796
rect 5760 2598 5816 2654
rect 5902 2598 5958 2654
rect 5760 2456 5816 2512
rect 5902 2456 5958 2512
rect 5760 2314 5816 2370
rect 5902 2314 5958 2370
rect 5760 2172 5816 2228
rect 5902 2172 5958 2228
rect 5760 2030 5816 2086
rect 5902 2030 5958 2086
rect 5760 1888 5816 1944
rect 5902 1888 5958 1944
rect 5760 1746 5816 1802
rect 5902 1746 5958 1802
rect 5760 1604 5816 1660
rect 5902 1604 5958 1660
rect 5760 1462 5816 1518
rect 5902 1462 5958 1518
rect 5760 1320 5816 1376
rect 5902 1320 5958 1376
rect 5760 1178 5816 1234
rect 5902 1178 5958 1234
rect 5760 1036 5816 1092
rect 5902 1036 5958 1092
rect 5760 894 5816 950
rect 5902 894 5958 950
rect 5760 752 5816 808
rect 5902 752 5958 808
rect 5760 610 5816 666
rect 5902 610 5958 666
rect 5760 468 5816 524
rect 5902 468 5958 524
rect 6300 12254 6356 12310
rect 6442 12254 6498 12310
rect 6300 12112 6356 12168
rect 6442 12112 6498 12168
rect 6300 11970 6356 12026
rect 6442 11970 6498 12026
rect 6300 11828 6356 11884
rect 6442 11828 6498 11884
rect 6300 11686 6356 11742
rect 6442 11686 6498 11742
rect 6300 11544 6356 11600
rect 6442 11544 6498 11600
rect 6300 11402 6356 11458
rect 6442 11402 6498 11458
rect 6300 11260 6356 11316
rect 6442 11260 6498 11316
rect 6300 11118 6356 11174
rect 6442 11118 6498 11174
rect 6300 10976 6356 11032
rect 6442 10976 6498 11032
rect 6300 10834 6356 10890
rect 6442 10834 6498 10890
rect 6300 10692 6356 10748
rect 6442 10692 6498 10748
rect 6300 10550 6356 10606
rect 6442 10550 6498 10606
rect 6300 10408 6356 10464
rect 6442 10408 6498 10464
rect 6300 10266 6356 10322
rect 6442 10266 6498 10322
rect 6300 10124 6356 10180
rect 6442 10124 6498 10180
rect 6300 9982 6356 10038
rect 6442 9982 6498 10038
rect 6300 9840 6356 9896
rect 6442 9840 6498 9896
rect 6300 9698 6356 9754
rect 6442 9698 6498 9754
rect 6300 9556 6356 9612
rect 6442 9556 6498 9612
rect 6300 9414 6356 9470
rect 6442 9414 6498 9470
rect 6300 9272 6356 9328
rect 6442 9272 6498 9328
rect 6300 9130 6356 9186
rect 6442 9130 6498 9186
rect 6300 8988 6356 9044
rect 6442 8988 6498 9044
rect 6300 8846 6356 8902
rect 6442 8846 6498 8902
rect 6300 8704 6356 8760
rect 6442 8704 6498 8760
rect 6300 8562 6356 8618
rect 6442 8562 6498 8618
rect 6300 8420 6356 8476
rect 6442 8420 6498 8476
rect 6300 8278 6356 8334
rect 6442 8278 6498 8334
rect 6300 8136 6356 8192
rect 6442 8136 6498 8192
rect 6300 7994 6356 8050
rect 6442 7994 6498 8050
rect 6300 7852 6356 7908
rect 6442 7852 6498 7908
rect 6300 7710 6356 7766
rect 6442 7710 6498 7766
rect 6300 7568 6356 7624
rect 6442 7568 6498 7624
rect 6300 7426 6356 7482
rect 6442 7426 6498 7482
rect 6300 7284 6356 7340
rect 6442 7284 6498 7340
rect 6300 7142 6356 7198
rect 6442 7142 6498 7198
rect 6300 7000 6356 7056
rect 6442 7000 6498 7056
rect 6300 6858 6356 6914
rect 6442 6858 6498 6914
rect 6300 6716 6356 6772
rect 6442 6716 6498 6772
rect 6300 6574 6356 6630
rect 6442 6574 6498 6630
rect 6300 6432 6356 6488
rect 6442 6432 6498 6488
rect 6300 6290 6356 6346
rect 6442 6290 6498 6346
rect 6300 6148 6356 6204
rect 6442 6148 6498 6204
rect 6300 6006 6356 6062
rect 6442 6006 6498 6062
rect 6300 5864 6356 5920
rect 6442 5864 6498 5920
rect 6300 5722 6356 5778
rect 6442 5722 6498 5778
rect 6300 5580 6356 5636
rect 6442 5580 6498 5636
rect 6300 5438 6356 5494
rect 6442 5438 6498 5494
rect 6300 5296 6356 5352
rect 6442 5296 6498 5352
rect 6300 5154 6356 5210
rect 6442 5154 6498 5210
rect 6300 5012 6356 5068
rect 6442 5012 6498 5068
rect 6300 4870 6356 4926
rect 6442 4870 6498 4926
rect 6300 4728 6356 4784
rect 6442 4728 6498 4784
rect 6300 4586 6356 4642
rect 6442 4586 6498 4642
rect 6300 4444 6356 4500
rect 6442 4444 6498 4500
rect 6300 4302 6356 4358
rect 6442 4302 6498 4358
rect 6300 4160 6356 4216
rect 6442 4160 6498 4216
rect 6300 4018 6356 4074
rect 6442 4018 6498 4074
rect 6300 3876 6356 3932
rect 6442 3876 6498 3932
rect 6300 3734 6356 3790
rect 6442 3734 6498 3790
rect 6300 3592 6356 3648
rect 6442 3592 6498 3648
rect 6300 3450 6356 3506
rect 6442 3450 6498 3506
rect 6300 3308 6356 3364
rect 6442 3308 6498 3364
rect 6300 3166 6356 3222
rect 6442 3166 6498 3222
rect 6300 3024 6356 3080
rect 6442 3024 6498 3080
rect 6300 2882 6356 2938
rect 6442 2882 6498 2938
rect 6300 2740 6356 2796
rect 6442 2740 6498 2796
rect 6300 2598 6356 2654
rect 6442 2598 6498 2654
rect 6300 2456 6356 2512
rect 6442 2456 6498 2512
rect 6300 2314 6356 2370
rect 6442 2314 6498 2370
rect 6300 2172 6356 2228
rect 6442 2172 6498 2228
rect 6300 2030 6356 2086
rect 6442 2030 6498 2086
rect 6300 1888 6356 1944
rect 6442 1888 6498 1944
rect 6300 1746 6356 1802
rect 6442 1746 6498 1802
rect 6300 1604 6356 1660
rect 6442 1604 6498 1660
rect 6300 1462 6356 1518
rect 6442 1462 6498 1518
rect 6300 1320 6356 1376
rect 6442 1320 6498 1376
rect 6300 1178 6356 1234
rect 6442 1178 6498 1234
rect 6300 1036 6356 1092
rect 6442 1036 6498 1092
rect 6300 894 6356 950
rect 6442 894 6498 950
rect 6300 752 6356 808
rect 6442 752 6498 808
rect 6300 610 6356 666
rect 6442 610 6498 666
rect 6300 468 6356 524
rect 6442 468 6498 524
rect 6845 12254 6901 12310
rect 6987 12254 7043 12310
rect 6845 12112 6901 12168
rect 6987 12112 7043 12168
rect 6845 11970 6901 12026
rect 6987 11970 7043 12026
rect 6845 11828 6901 11884
rect 6987 11828 7043 11884
rect 6845 11686 6901 11742
rect 6987 11686 7043 11742
rect 6845 11544 6901 11600
rect 6987 11544 7043 11600
rect 6845 11402 6901 11458
rect 6987 11402 7043 11458
rect 6845 11260 6901 11316
rect 6987 11260 7043 11316
rect 6845 11118 6901 11174
rect 6987 11118 7043 11174
rect 6845 10976 6901 11032
rect 6987 10976 7043 11032
rect 6845 10834 6901 10890
rect 6987 10834 7043 10890
rect 6845 10692 6901 10748
rect 6987 10692 7043 10748
rect 6845 10550 6901 10606
rect 6987 10550 7043 10606
rect 6845 10408 6901 10464
rect 6987 10408 7043 10464
rect 6845 10266 6901 10322
rect 6987 10266 7043 10322
rect 6845 10124 6901 10180
rect 6987 10124 7043 10180
rect 6845 9982 6901 10038
rect 6987 9982 7043 10038
rect 6845 9840 6901 9896
rect 6987 9840 7043 9896
rect 6845 9698 6901 9754
rect 6987 9698 7043 9754
rect 6845 9556 6901 9612
rect 6987 9556 7043 9612
rect 6845 9414 6901 9470
rect 6987 9414 7043 9470
rect 6845 9272 6901 9328
rect 6987 9272 7043 9328
rect 6845 9130 6901 9186
rect 6987 9130 7043 9186
rect 6845 8988 6901 9044
rect 6987 8988 7043 9044
rect 6845 8846 6901 8902
rect 6987 8846 7043 8902
rect 6845 8704 6901 8760
rect 6987 8704 7043 8760
rect 6845 8562 6901 8618
rect 6987 8562 7043 8618
rect 6845 8420 6901 8476
rect 6987 8420 7043 8476
rect 6845 8278 6901 8334
rect 6987 8278 7043 8334
rect 6845 8136 6901 8192
rect 6987 8136 7043 8192
rect 6845 7994 6901 8050
rect 6987 7994 7043 8050
rect 6845 7852 6901 7908
rect 6987 7852 7043 7908
rect 6845 7710 6901 7766
rect 6987 7710 7043 7766
rect 6845 7568 6901 7624
rect 6987 7568 7043 7624
rect 6845 7426 6901 7482
rect 6987 7426 7043 7482
rect 6845 7284 6901 7340
rect 6987 7284 7043 7340
rect 6845 7142 6901 7198
rect 6987 7142 7043 7198
rect 6845 7000 6901 7056
rect 6987 7000 7043 7056
rect 6845 6858 6901 6914
rect 6987 6858 7043 6914
rect 6845 6716 6901 6772
rect 6987 6716 7043 6772
rect 6845 6574 6901 6630
rect 6987 6574 7043 6630
rect 6845 6432 6901 6488
rect 6987 6432 7043 6488
rect 6845 6290 6901 6346
rect 6987 6290 7043 6346
rect 6845 6148 6901 6204
rect 6987 6148 7043 6204
rect 6845 6006 6901 6062
rect 6987 6006 7043 6062
rect 6845 5864 6901 5920
rect 6987 5864 7043 5920
rect 6845 5722 6901 5778
rect 6987 5722 7043 5778
rect 6845 5580 6901 5636
rect 6987 5580 7043 5636
rect 6845 5438 6901 5494
rect 6987 5438 7043 5494
rect 6845 5296 6901 5352
rect 6987 5296 7043 5352
rect 6845 5154 6901 5210
rect 6987 5154 7043 5210
rect 6845 5012 6901 5068
rect 6987 5012 7043 5068
rect 6845 4870 6901 4926
rect 6987 4870 7043 4926
rect 6845 4728 6901 4784
rect 6987 4728 7043 4784
rect 6845 4586 6901 4642
rect 6987 4586 7043 4642
rect 6845 4444 6901 4500
rect 6987 4444 7043 4500
rect 6845 4302 6901 4358
rect 6987 4302 7043 4358
rect 6845 4160 6901 4216
rect 6987 4160 7043 4216
rect 6845 4018 6901 4074
rect 6987 4018 7043 4074
rect 6845 3876 6901 3932
rect 6987 3876 7043 3932
rect 6845 3734 6901 3790
rect 6987 3734 7043 3790
rect 6845 3592 6901 3648
rect 6987 3592 7043 3648
rect 6845 3450 6901 3506
rect 6987 3450 7043 3506
rect 6845 3308 6901 3364
rect 6987 3308 7043 3364
rect 6845 3166 6901 3222
rect 6987 3166 7043 3222
rect 6845 3024 6901 3080
rect 6987 3024 7043 3080
rect 6845 2882 6901 2938
rect 6987 2882 7043 2938
rect 6845 2740 6901 2796
rect 6987 2740 7043 2796
rect 6845 2598 6901 2654
rect 6987 2598 7043 2654
rect 6845 2456 6901 2512
rect 6987 2456 7043 2512
rect 6845 2314 6901 2370
rect 6987 2314 7043 2370
rect 6845 2172 6901 2228
rect 6987 2172 7043 2228
rect 6845 2030 6901 2086
rect 6987 2030 7043 2086
rect 6845 1888 6901 1944
rect 6987 1888 7043 1944
rect 6845 1746 6901 1802
rect 6987 1746 7043 1802
rect 6845 1604 6901 1660
rect 6987 1604 7043 1660
rect 6845 1462 6901 1518
rect 6987 1462 7043 1518
rect 6845 1320 6901 1376
rect 6987 1320 7043 1376
rect 6845 1178 6901 1234
rect 6987 1178 7043 1234
rect 6845 1036 6901 1092
rect 6987 1036 7043 1092
rect 6845 894 6901 950
rect 6987 894 7043 950
rect 6845 752 6901 808
rect 6987 752 7043 808
rect 6845 610 6901 666
rect 6987 610 7043 666
rect 6845 468 6901 524
rect 6987 468 7043 524
rect 7382 12254 7438 12310
rect 7524 12254 7580 12310
rect 7382 12112 7438 12168
rect 7524 12112 7580 12168
rect 7382 11970 7438 12026
rect 7524 11970 7580 12026
rect 7382 11828 7438 11884
rect 7524 11828 7580 11884
rect 7382 11686 7438 11742
rect 7524 11686 7580 11742
rect 7382 11544 7438 11600
rect 7524 11544 7580 11600
rect 7382 11402 7438 11458
rect 7524 11402 7580 11458
rect 7382 11260 7438 11316
rect 7524 11260 7580 11316
rect 7382 11118 7438 11174
rect 7524 11118 7580 11174
rect 7382 10976 7438 11032
rect 7524 10976 7580 11032
rect 7382 10834 7438 10890
rect 7524 10834 7580 10890
rect 7382 10692 7438 10748
rect 7524 10692 7580 10748
rect 7382 10550 7438 10606
rect 7524 10550 7580 10606
rect 7382 10408 7438 10464
rect 7524 10408 7580 10464
rect 7382 10266 7438 10322
rect 7524 10266 7580 10322
rect 7382 10124 7438 10180
rect 7524 10124 7580 10180
rect 7382 9982 7438 10038
rect 7524 9982 7580 10038
rect 7382 9840 7438 9896
rect 7524 9840 7580 9896
rect 7382 9698 7438 9754
rect 7524 9698 7580 9754
rect 7382 9556 7438 9612
rect 7524 9556 7580 9612
rect 7382 9414 7438 9470
rect 7524 9414 7580 9470
rect 7382 9272 7438 9328
rect 7524 9272 7580 9328
rect 7382 9130 7438 9186
rect 7524 9130 7580 9186
rect 7382 8988 7438 9044
rect 7524 8988 7580 9044
rect 7382 8846 7438 8902
rect 7524 8846 7580 8902
rect 7382 8704 7438 8760
rect 7524 8704 7580 8760
rect 7382 8562 7438 8618
rect 7524 8562 7580 8618
rect 7382 8420 7438 8476
rect 7524 8420 7580 8476
rect 7382 8278 7438 8334
rect 7524 8278 7580 8334
rect 7382 8136 7438 8192
rect 7524 8136 7580 8192
rect 7382 7994 7438 8050
rect 7524 7994 7580 8050
rect 7382 7852 7438 7908
rect 7524 7852 7580 7908
rect 7382 7710 7438 7766
rect 7524 7710 7580 7766
rect 7382 7568 7438 7624
rect 7524 7568 7580 7624
rect 7382 7426 7438 7482
rect 7524 7426 7580 7482
rect 7382 7284 7438 7340
rect 7524 7284 7580 7340
rect 7382 7142 7438 7198
rect 7524 7142 7580 7198
rect 7382 7000 7438 7056
rect 7524 7000 7580 7056
rect 7382 6858 7438 6914
rect 7524 6858 7580 6914
rect 7382 6716 7438 6772
rect 7524 6716 7580 6772
rect 7382 6574 7438 6630
rect 7524 6574 7580 6630
rect 7382 6432 7438 6488
rect 7524 6432 7580 6488
rect 7382 6290 7438 6346
rect 7524 6290 7580 6346
rect 7382 6148 7438 6204
rect 7524 6148 7580 6204
rect 7382 6006 7438 6062
rect 7524 6006 7580 6062
rect 7382 5864 7438 5920
rect 7524 5864 7580 5920
rect 7382 5722 7438 5778
rect 7524 5722 7580 5778
rect 7382 5580 7438 5636
rect 7524 5580 7580 5636
rect 7382 5438 7438 5494
rect 7524 5438 7580 5494
rect 7382 5296 7438 5352
rect 7524 5296 7580 5352
rect 7382 5154 7438 5210
rect 7524 5154 7580 5210
rect 7382 5012 7438 5068
rect 7524 5012 7580 5068
rect 7382 4870 7438 4926
rect 7524 4870 7580 4926
rect 7382 4728 7438 4784
rect 7524 4728 7580 4784
rect 7382 4586 7438 4642
rect 7524 4586 7580 4642
rect 7382 4444 7438 4500
rect 7524 4444 7580 4500
rect 7382 4302 7438 4358
rect 7524 4302 7580 4358
rect 7382 4160 7438 4216
rect 7524 4160 7580 4216
rect 7382 4018 7438 4074
rect 7524 4018 7580 4074
rect 7382 3876 7438 3932
rect 7524 3876 7580 3932
rect 7382 3734 7438 3790
rect 7524 3734 7580 3790
rect 7382 3592 7438 3648
rect 7524 3592 7580 3648
rect 7382 3450 7438 3506
rect 7524 3450 7580 3506
rect 7382 3308 7438 3364
rect 7524 3308 7580 3364
rect 7382 3166 7438 3222
rect 7524 3166 7580 3222
rect 7382 3024 7438 3080
rect 7524 3024 7580 3080
rect 7382 2882 7438 2938
rect 7524 2882 7580 2938
rect 7382 2740 7438 2796
rect 7524 2740 7580 2796
rect 7382 2598 7438 2654
rect 7524 2598 7580 2654
rect 7382 2456 7438 2512
rect 7524 2456 7580 2512
rect 7382 2314 7438 2370
rect 7524 2314 7580 2370
rect 7382 2172 7438 2228
rect 7524 2172 7580 2228
rect 7382 2030 7438 2086
rect 7524 2030 7580 2086
rect 7382 1888 7438 1944
rect 7524 1888 7580 1944
rect 7382 1746 7438 1802
rect 7524 1746 7580 1802
rect 7382 1604 7438 1660
rect 7524 1604 7580 1660
rect 7382 1462 7438 1518
rect 7524 1462 7580 1518
rect 7382 1320 7438 1376
rect 7524 1320 7580 1376
rect 7382 1178 7438 1234
rect 7524 1178 7580 1234
rect 7382 1036 7438 1092
rect 7524 1036 7580 1092
rect 7382 894 7438 950
rect 7524 894 7580 950
rect 7382 752 7438 808
rect 7524 752 7580 808
rect 7382 610 7438 666
rect 7524 610 7580 666
rect 7382 468 7438 524
rect 7524 468 7580 524
rect 7919 12254 7975 12310
rect 8061 12254 8117 12310
rect 7919 12112 7975 12168
rect 8061 12112 8117 12168
rect 7919 11970 7975 12026
rect 8061 11970 8117 12026
rect 7919 11828 7975 11884
rect 8061 11828 8117 11884
rect 7919 11686 7975 11742
rect 8061 11686 8117 11742
rect 7919 11544 7975 11600
rect 8061 11544 8117 11600
rect 7919 11402 7975 11458
rect 8061 11402 8117 11458
rect 7919 11260 7975 11316
rect 8061 11260 8117 11316
rect 7919 11118 7975 11174
rect 8061 11118 8117 11174
rect 7919 10976 7975 11032
rect 8061 10976 8117 11032
rect 7919 10834 7975 10890
rect 8061 10834 8117 10890
rect 7919 10692 7975 10748
rect 8061 10692 8117 10748
rect 7919 10550 7975 10606
rect 8061 10550 8117 10606
rect 7919 10408 7975 10464
rect 8061 10408 8117 10464
rect 7919 10266 7975 10322
rect 8061 10266 8117 10322
rect 7919 10124 7975 10180
rect 8061 10124 8117 10180
rect 7919 9982 7975 10038
rect 8061 9982 8117 10038
rect 7919 9840 7975 9896
rect 8061 9840 8117 9896
rect 7919 9698 7975 9754
rect 8061 9698 8117 9754
rect 7919 9556 7975 9612
rect 8061 9556 8117 9612
rect 7919 9414 7975 9470
rect 8061 9414 8117 9470
rect 7919 9272 7975 9328
rect 8061 9272 8117 9328
rect 7919 9130 7975 9186
rect 8061 9130 8117 9186
rect 7919 8988 7975 9044
rect 8061 8988 8117 9044
rect 7919 8846 7975 8902
rect 8061 8846 8117 8902
rect 7919 8704 7975 8760
rect 8061 8704 8117 8760
rect 7919 8562 7975 8618
rect 8061 8562 8117 8618
rect 7919 8420 7975 8476
rect 8061 8420 8117 8476
rect 7919 8278 7975 8334
rect 8061 8278 8117 8334
rect 7919 8136 7975 8192
rect 8061 8136 8117 8192
rect 7919 7994 7975 8050
rect 8061 7994 8117 8050
rect 7919 7852 7975 7908
rect 8061 7852 8117 7908
rect 7919 7710 7975 7766
rect 8061 7710 8117 7766
rect 7919 7568 7975 7624
rect 8061 7568 8117 7624
rect 7919 7426 7975 7482
rect 8061 7426 8117 7482
rect 7919 7284 7975 7340
rect 8061 7284 8117 7340
rect 7919 7142 7975 7198
rect 8061 7142 8117 7198
rect 7919 7000 7975 7056
rect 8061 7000 8117 7056
rect 7919 6858 7975 6914
rect 8061 6858 8117 6914
rect 7919 6716 7975 6772
rect 8061 6716 8117 6772
rect 7919 6574 7975 6630
rect 8061 6574 8117 6630
rect 7919 6432 7975 6488
rect 8061 6432 8117 6488
rect 7919 6290 7975 6346
rect 8061 6290 8117 6346
rect 7919 6148 7975 6204
rect 8061 6148 8117 6204
rect 7919 6006 7975 6062
rect 8061 6006 8117 6062
rect 7919 5864 7975 5920
rect 8061 5864 8117 5920
rect 7919 5722 7975 5778
rect 8061 5722 8117 5778
rect 7919 5580 7975 5636
rect 8061 5580 8117 5636
rect 7919 5438 7975 5494
rect 8061 5438 8117 5494
rect 7919 5296 7975 5352
rect 8061 5296 8117 5352
rect 7919 5154 7975 5210
rect 8061 5154 8117 5210
rect 7919 5012 7975 5068
rect 8061 5012 8117 5068
rect 7919 4870 7975 4926
rect 8061 4870 8117 4926
rect 7919 4728 7975 4784
rect 8061 4728 8117 4784
rect 7919 4586 7975 4642
rect 8061 4586 8117 4642
rect 7919 4444 7975 4500
rect 8061 4444 8117 4500
rect 7919 4302 7975 4358
rect 8061 4302 8117 4358
rect 7919 4160 7975 4216
rect 8061 4160 8117 4216
rect 7919 4018 7975 4074
rect 8061 4018 8117 4074
rect 7919 3876 7975 3932
rect 8061 3876 8117 3932
rect 7919 3734 7975 3790
rect 8061 3734 8117 3790
rect 7919 3592 7975 3648
rect 8061 3592 8117 3648
rect 7919 3450 7975 3506
rect 8061 3450 8117 3506
rect 7919 3308 7975 3364
rect 8061 3308 8117 3364
rect 7919 3166 7975 3222
rect 8061 3166 8117 3222
rect 7919 3024 7975 3080
rect 8061 3024 8117 3080
rect 7919 2882 7975 2938
rect 8061 2882 8117 2938
rect 7919 2740 7975 2796
rect 8061 2740 8117 2796
rect 7919 2598 7975 2654
rect 8061 2598 8117 2654
rect 7919 2456 7975 2512
rect 8061 2456 8117 2512
rect 7919 2314 7975 2370
rect 8061 2314 8117 2370
rect 7919 2172 7975 2228
rect 8061 2172 8117 2228
rect 7919 2030 7975 2086
rect 8061 2030 8117 2086
rect 7919 1888 7975 1944
rect 8061 1888 8117 1944
rect 7919 1746 7975 1802
rect 8061 1746 8117 1802
rect 7919 1604 7975 1660
rect 8061 1604 8117 1660
rect 7919 1462 7975 1518
rect 8061 1462 8117 1518
rect 7919 1320 7975 1376
rect 8061 1320 8117 1376
rect 7919 1178 7975 1234
rect 8061 1178 8117 1234
rect 7919 1036 7975 1092
rect 8061 1036 8117 1092
rect 7919 894 7975 950
rect 8061 894 8117 950
rect 7919 752 7975 808
rect 8061 752 8117 808
rect 7919 610 7975 666
rect 8061 610 8117 666
rect 7919 468 7975 524
rect 8061 468 8117 524
rect 8462 12254 8518 12310
rect 8604 12254 8660 12310
rect 8462 12112 8518 12168
rect 8604 12112 8660 12168
rect 8462 11970 8518 12026
rect 8604 11970 8660 12026
rect 8462 11828 8518 11884
rect 8604 11828 8660 11884
rect 8462 11686 8518 11742
rect 8604 11686 8660 11742
rect 8462 11544 8518 11600
rect 8604 11544 8660 11600
rect 8462 11402 8518 11458
rect 8604 11402 8660 11458
rect 8462 11260 8518 11316
rect 8604 11260 8660 11316
rect 8462 11118 8518 11174
rect 8604 11118 8660 11174
rect 8462 10976 8518 11032
rect 8604 10976 8660 11032
rect 8462 10834 8518 10890
rect 8604 10834 8660 10890
rect 8462 10692 8518 10748
rect 8604 10692 8660 10748
rect 8462 10550 8518 10606
rect 8604 10550 8660 10606
rect 8462 10408 8518 10464
rect 8604 10408 8660 10464
rect 8462 10266 8518 10322
rect 8604 10266 8660 10322
rect 8462 10124 8518 10180
rect 8604 10124 8660 10180
rect 8462 9982 8518 10038
rect 8604 9982 8660 10038
rect 8462 9840 8518 9896
rect 8604 9840 8660 9896
rect 8462 9698 8518 9754
rect 8604 9698 8660 9754
rect 8462 9556 8518 9612
rect 8604 9556 8660 9612
rect 8462 9414 8518 9470
rect 8604 9414 8660 9470
rect 8462 9272 8518 9328
rect 8604 9272 8660 9328
rect 8462 9130 8518 9186
rect 8604 9130 8660 9186
rect 8462 8988 8518 9044
rect 8604 8988 8660 9044
rect 8462 8846 8518 8902
rect 8604 8846 8660 8902
rect 8462 8704 8518 8760
rect 8604 8704 8660 8760
rect 8462 8562 8518 8618
rect 8604 8562 8660 8618
rect 8462 8420 8518 8476
rect 8604 8420 8660 8476
rect 8462 8278 8518 8334
rect 8604 8278 8660 8334
rect 8462 8136 8518 8192
rect 8604 8136 8660 8192
rect 8462 7994 8518 8050
rect 8604 7994 8660 8050
rect 8462 7852 8518 7908
rect 8604 7852 8660 7908
rect 8462 7710 8518 7766
rect 8604 7710 8660 7766
rect 8462 7568 8518 7624
rect 8604 7568 8660 7624
rect 8462 7426 8518 7482
rect 8604 7426 8660 7482
rect 8462 7284 8518 7340
rect 8604 7284 8660 7340
rect 8462 7142 8518 7198
rect 8604 7142 8660 7198
rect 8462 7000 8518 7056
rect 8604 7000 8660 7056
rect 8462 6858 8518 6914
rect 8604 6858 8660 6914
rect 8462 6716 8518 6772
rect 8604 6716 8660 6772
rect 8462 6574 8518 6630
rect 8604 6574 8660 6630
rect 8462 6432 8518 6488
rect 8604 6432 8660 6488
rect 8462 6290 8518 6346
rect 8604 6290 8660 6346
rect 8462 6148 8518 6204
rect 8604 6148 8660 6204
rect 8462 6006 8518 6062
rect 8604 6006 8660 6062
rect 8462 5864 8518 5920
rect 8604 5864 8660 5920
rect 8462 5722 8518 5778
rect 8604 5722 8660 5778
rect 8462 5580 8518 5636
rect 8604 5580 8660 5636
rect 8462 5438 8518 5494
rect 8604 5438 8660 5494
rect 8462 5296 8518 5352
rect 8604 5296 8660 5352
rect 8462 5154 8518 5210
rect 8604 5154 8660 5210
rect 8462 5012 8518 5068
rect 8604 5012 8660 5068
rect 8462 4870 8518 4926
rect 8604 4870 8660 4926
rect 8462 4728 8518 4784
rect 8604 4728 8660 4784
rect 8462 4586 8518 4642
rect 8604 4586 8660 4642
rect 8462 4444 8518 4500
rect 8604 4444 8660 4500
rect 8462 4302 8518 4358
rect 8604 4302 8660 4358
rect 8462 4160 8518 4216
rect 8604 4160 8660 4216
rect 8462 4018 8518 4074
rect 8604 4018 8660 4074
rect 8462 3876 8518 3932
rect 8604 3876 8660 3932
rect 8462 3734 8518 3790
rect 8604 3734 8660 3790
rect 8462 3592 8518 3648
rect 8604 3592 8660 3648
rect 8462 3450 8518 3506
rect 8604 3450 8660 3506
rect 8462 3308 8518 3364
rect 8604 3308 8660 3364
rect 8462 3166 8518 3222
rect 8604 3166 8660 3222
rect 8462 3024 8518 3080
rect 8604 3024 8660 3080
rect 8462 2882 8518 2938
rect 8604 2882 8660 2938
rect 8462 2740 8518 2796
rect 8604 2740 8660 2796
rect 8462 2598 8518 2654
rect 8604 2598 8660 2654
rect 8462 2456 8518 2512
rect 8604 2456 8660 2512
rect 8462 2314 8518 2370
rect 8604 2314 8660 2370
rect 8462 2172 8518 2228
rect 8604 2172 8660 2228
rect 8462 2030 8518 2086
rect 8604 2030 8660 2086
rect 8462 1888 8518 1944
rect 8604 1888 8660 1944
rect 8462 1746 8518 1802
rect 8604 1746 8660 1802
rect 8462 1604 8518 1660
rect 8604 1604 8660 1660
rect 8462 1462 8518 1518
rect 8604 1462 8660 1518
rect 8462 1320 8518 1376
rect 8604 1320 8660 1376
rect 8462 1178 8518 1234
rect 8604 1178 8660 1234
rect 8462 1036 8518 1092
rect 8604 1036 8660 1092
rect 8462 894 8518 950
rect 8604 894 8660 950
rect 8462 752 8518 808
rect 8604 752 8660 808
rect 8462 610 8518 666
rect 8604 610 8660 666
rect 8462 468 8518 524
rect 8604 468 8660 524
rect 9004 12254 9060 12310
rect 9146 12254 9202 12310
rect 9004 12112 9060 12168
rect 9146 12112 9202 12168
rect 9004 11970 9060 12026
rect 9146 11970 9202 12026
rect 9004 11828 9060 11884
rect 9146 11828 9202 11884
rect 9004 11686 9060 11742
rect 9146 11686 9202 11742
rect 9004 11544 9060 11600
rect 9146 11544 9202 11600
rect 9004 11402 9060 11458
rect 9146 11402 9202 11458
rect 9004 11260 9060 11316
rect 9146 11260 9202 11316
rect 9004 11118 9060 11174
rect 9146 11118 9202 11174
rect 9004 10976 9060 11032
rect 9146 10976 9202 11032
rect 9004 10834 9060 10890
rect 9146 10834 9202 10890
rect 9004 10692 9060 10748
rect 9146 10692 9202 10748
rect 9004 10550 9060 10606
rect 9146 10550 9202 10606
rect 9004 10408 9060 10464
rect 9146 10408 9202 10464
rect 9004 10266 9060 10322
rect 9146 10266 9202 10322
rect 9004 10124 9060 10180
rect 9146 10124 9202 10180
rect 9004 9982 9060 10038
rect 9146 9982 9202 10038
rect 9004 9840 9060 9896
rect 9146 9840 9202 9896
rect 9004 9698 9060 9754
rect 9146 9698 9202 9754
rect 9004 9556 9060 9612
rect 9146 9556 9202 9612
rect 9004 9414 9060 9470
rect 9146 9414 9202 9470
rect 9004 9272 9060 9328
rect 9146 9272 9202 9328
rect 9004 9130 9060 9186
rect 9146 9130 9202 9186
rect 9004 8988 9060 9044
rect 9146 8988 9202 9044
rect 9004 8846 9060 8902
rect 9146 8846 9202 8902
rect 9004 8704 9060 8760
rect 9146 8704 9202 8760
rect 9004 8562 9060 8618
rect 9146 8562 9202 8618
rect 9004 8420 9060 8476
rect 9146 8420 9202 8476
rect 9004 8278 9060 8334
rect 9146 8278 9202 8334
rect 9004 8136 9060 8192
rect 9146 8136 9202 8192
rect 9004 7994 9060 8050
rect 9146 7994 9202 8050
rect 9004 7852 9060 7908
rect 9146 7852 9202 7908
rect 9004 7710 9060 7766
rect 9146 7710 9202 7766
rect 9004 7568 9060 7624
rect 9146 7568 9202 7624
rect 9004 7426 9060 7482
rect 9146 7426 9202 7482
rect 9004 7284 9060 7340
rect 9146 7284 9202 7340
rect 9004 7142 9060 7198
rect 9146 7142 9202 7198
rect 9004 7000 9060 7056
rect 9146 7000 9202 7056
rect 9004 6858 9060 6914
rect 9146 6858 9202 6914
rect 9004 6716 9060 6772
rect 9146 6716 9202 6772
rect 9004 6574 9060 6630
rect 9146 6574 9202 6630
rect 9004 6432 9060 6488
rect 9146 6432 9202 6488
rect 9004 6290 9060 6346
rect 9146 6290 9202 6346
rect 9004 6148 9060 6204
rect 9146 6148 9202 6204
rect 9004 6006 9060 6062
rect 9146 6006 9202 6062
rect 9004 5864 9060 5920
rect 9146 5864 9202 5920
rect 9004 5722 9060 5778
rect 9146 5722 9202 5778
rect 9004 5580 9060 5636
rect 9146 5580 9202 5636
rect 9004 5438 9060 5494
rect 9146 5438 9202 5494
rect 9004 5296 9060 5352
rect 9146 5296 9202 5352
rect 9004 5154 9060 5210
rect 9146 5154 9202 5210
rect 9004 5012 9060 5068
rect 9146 5012 9202 5068
rect 9004 4870 9060 4926
rect 9146 4870 9202 4926
rect 9004 4728 9060 4784
rect 9146 4728 9202 4784
rect 9004 4586 9060 4642
rect 9146 4586 9202 4642
rect 9004 4444 9060 4500
rect 9146 4444 9202 4500
rect 9004 4302 9060 4358
rect 9146 4302 9202 4358
rect 9004 4160 9060 4216
rect 9146 4160 9202 4216
rect 9004 4018 9060 4074
rect 9146 4018 9202 4074
rect 9004 3876 9060 3932
rect 9146 3876 9202 3932
rect 9004 3734 9060 3790
rect 9146 3734 9202 3790
rect 9004 3592 9060 3648
rect 9146 3592 9202 3648
rect 9004 3450 9060 3506
rect 9146 3450 9202 3506
rect 9004 3308 9060 3364
rect 9146 3308 9202 3364
rect 9004 3166 9060 3222
rect 9146 3166 9202 3222
rect 9004 3024 9060 3080
rect 9146 3024 9202 3080
rect 9004 2882 9060 2938
rect 9146 2882 9202 2938
rect 9004 2740 9060 2796
rect 9146 2740 9202 2796
rect 9004 2598 9060 2654
rect 9146 2598 9202 2654
rect 9004 2456 9060 2512
rect 9146 2456 9202 2512
rect 9004 2314 9060 2370
rect 9146 2314 9202 2370
rect 9004 2172 9060 2228
rect 9146 2172 9202 2228
rect 9004 2030 9060 2086
rect 9146 2030 9202 2086
rect 9004 1888 9060 1944
rect 9146 1888 9202 1944
rect 9004 1746 9060 1802
rect 9146 1746 9202 1802
rect 9004 1604 9060 1660
rect 9146 1604 9202 1660
rect 9004 1462 9060 1518
rect 9146 1462 9202 1518
rect 9004 1320 9060 1376
rect 9146 1320 9202 1376
rect 9004 1178 9060 1234
rect 9146 1178 9202 1234
rect 9004 1036 9060 1092
rect 9146 1036 9202 1092
rect 9004 894 9060 950
rect 9146 894 9202 950
rect 9004 752 9060 808
rect 9146 752 9202 808
rect 9004 610 9060 666
rect 9146 610 9202 666
rect 9004 468 9060 524
rect 9146 468 9202 524
rect 9547 12254 9603 12310
rect 9689 12254 9745 12310
rect 9547 12112 9603 12168
rect 9689 12112 9745 12168
rect 9547 11970 9603 12026
rect 9689 11970 9745 12026
rect 9547 11828 9603 11884
rect 9689 11828 9745 11884
rect 9547 11686 9603 11742
rect 9689 11686 9745 11742
rect 9547 11544 9603 11600
rect 9689 11544 9745 11600
rect 9547 11402 9603 11458
rect 9689 11402 9745 11458
rect 9547 11260 9603 11316
rect 9689 11260 9745 11316
rect 9547 11118 9603 11174
rect 9689 11118 9745 11174
rect 9547 10976 9603 11032
rect 9689 10976 9745 11032
rect 9547 10834 9603 10890
rect 9689 10834 9745 10890
rect 9547 10692 9603 10748
rect 9689 10692 9745 10748
rect 9547 10550 9603 10606
rect 9689 10550 9745 10606
rect 9547 10408 9603 10464
rect 9689 10408 9745 10464
rect 9547 10266 9603 10322
rect 9689 10266 9745 10322
rect 9547 10124 9603 10180
rect 9689 10124 9745 10180
rect 9547 9982 9603 10038
rect 9689 9982 9745 10038
rect 9547 9840 9603 9896
rect 9689 9840 9745 9896
rect 9547 9698 9603 9754
rect 9689 9698 9745 9754
rect 9547 9556 9603 9612
rect 9689 9556 9745 9612
rect 9547 9414 9603 9470
rect 9689 9414 9745 9470
rect 9547 9272 9603 9328
rect 9689 9272 9745 9328
rect 9547 9130 9603 9186
rect 9689 9130 9745 9186
rect 9547 8988 9603 9044
rect 9689 8988 9745 9044
rect 9547 8846 9603 8902
rect 9689 8846 9745 8902
rect 9547 8704 9603 8760
rect 9689 8704 9745 8760
rect 9547 8562 9603 8618
rect 9689 8562 9745 8618
rect 9547 8420 9603 8476
rect 9689 8420 9745 8476
rect 9547 8278 9603 8334
rect 9689 8278 9745 8334
rect 9547 8136 9603 8192
rect 9689 8136 9745 8192
rect 9547 7994 9603 8050
rect 9689 7994 9745 8050
rect 9547 7852 9603 7908
rect 9689 7852 9745 7908
rect 9547 7710 9603 7766
rect 9689 7710 9745 7766
rect 9547 7568 9603 7624
rect 9689 7568 9745 7624
rect 9547 7426 9603 7482
rect 9689 7426 9745 7482
rect 9547 7284 9603 7340
rect 9689 7284 9745 7340
rect 9547 7142 9603 7198
rect 9689 7142 9745 7198
rect 9547 7000 9603 7056
rect 9689 7000 9745 7056
rect 9547 6858 9603 6914
rect 9689 6858 9745 6914
rect 9547 6716 9603 6772
rect 9689 6716 9745 6772
rect 9547 6574 9603 6630
rect 9689 6574 9745 6630
rect 9547 6432 9603 6488
rect 9689 6432 9745 6488
rect 9547 6290 9603 6346
rect 9689 6290 9745 6346
rect 9547 6148 9603 6204
rect 9689 6148 9745 6204
rect 9547 6006 9603 6062
rect 9689 6006 9745 6062
rect 9547 5864 9603 5920
rect 9689 5864 9745 5920
rect 9547 5722 9603 5778
rect 9689 5722 9745 5778
rect 9547 5580 9603 5636
rect 9689 5580 9745 5636
rect 9547 5438 9603 5494
rect 9689 5438 9745 5494
rect 9547 5296 9603 5352
rect 9689 5296 9745 5352
rect 9547 5154 9603 5210
rect 9689 5154 9745 5210
rect 9547 5012 9603 5068
rect 9689 5012 9745 5068
rect 9547 4870 9603 4926
rect 9689 4870 9745 4926
rect 9547 4728 9603 4784
rect 9689 4728 9745 4784
rect 9547 4586 9603 4642
rect 9689 4586 9745 4642
rect 9547 4444 9603 4500
rect 9689 4444 9745 4500
rect 9547 4302 9603 4358
rect 9689 4302 9745 4358
rect 9547 4160 9603 4216
rect 9689 4160 9745 4216
rect 9547 4018 9603 4074
rect 9689 4018 9745 4074
rect 9547 3876 9603 3932
rect 9689 3876 9745 3932
rect 9547 3734 9603 3790
rect 9689 3734 9745 3790
rect 9547 3592 9603 3648
rect 9689 3592 9745 3648
rect 9547 3450 9603 3506
rect 9689 3450 9745 3506
rect 9547 3308 9603 3364
rect 9689 3308 9745 3364
rect 9547 3166 9603 3222
rect 9689 3166 9745 3222
rect 9547 3024 9603 3080
rect 9689 3024 9745 3080
rect 9547 2882 9603 2938
rect 9689 2882 9745 2938
rect 9547 2740 9603 2796
rect 9689 2740 9745 2796
rect 9547 2598 9603 2654
rect 9689 2598 9745 2654
rect 9547 2456 9603 2512
rect 9689 2456 9745 2512
rect 9547 2314 9603 2370
rect 9689 2314 9745 2370
rect 9547 2172 9603 2228
rect 9689 2172 9745 2228
rect 9547 2030 9603 2086
rect 9689 2030 9745 2086
rect 9547 1888 9603 1944
rect 9689 1888 9745 1944
rect 9547 1746 9603 1802
rect 9689 1746 9745 1802
rect 9547 1604 9603 1660
rect 9689 1604 9745 1660
rect 9547 1462 9603 1518
rect 9689 1462 9745 1518
rect 9547 1320 9603 1376
rect 9689 1320 9745 1376
rect 9547 1178 9603 1234
rect 9689 1178 9745 1234
rect 9547 1036 9603 1092
rect 9689 1036 9745 1092
rect 9547 894 9603 950
rect 9689 894 9745 950
rect 9547 752 9603 808
rect 9689 752 9745 808
rect 9547 610 9603 666
rect 9689 610 9745 666
rect 9547 468 9603 524
rect 9689 468 9745 524
rect 10081 12254 10137 12310
rect 10223 12254 10279 12310
rect 10081 12112 10137 12168
rect 10223 12112 10279 12168
rect 10081 11970 10137 12026
rect 10223 11970 10279 12026
rect 10081 11828 10137 11884
rect 10223 11828 10279 11884
rect 10081 11686 10137 11742
rect 10223 11686 10279 11742
rect 10081 11544 10137 11600
rect 10223 11544 10279 11600
rect 10081 11402 10137 11458
rect 10223 11402 10279 11458
rect 10081 11260 10137 11316
rect 10223 11260 10279 11316
rect 10081 11118 10137 11174
rect 10223 11118 10279 11174
rect 10081 10976 10137 11032
rect 10223 10976 10279 11032
rect 10081 10834 10137 10890
rect 10223 10834 10279 10890
rect 10081 10692 10137 10748
rect 10223 10692 10279 10748
rect 10081 10550 10137 10606
rect 10223 10550 10279 10606
rect 10081 10408 10137 10464
rect 10223 10408 10279 10464
rect 10081 10266 10137 10322
rect 10223 10266 10279 10322
rect 10081 10124 10137 10180
rect 10223 10124 10279 10180
rect 10081 9982 10137 10038
rect 10223 9982 10279 10038
rect 10081 9840 10137 9896
rect 10223 9840 10279 9896
rect 10081 9698 10137 9754
rect 10223 9698 10279 9754
rect 10081 9556 10137 9612
rect 10223 9556 10279 9612
rect 10081 9414 10137 9470
rect 10223 9414 10279 9470
rect 10081 9272 10137 9328
rect 10223 9272 10279 9328
rect 10081 9130 10137 9186
rect 10223 9130 10279 9186
rect 10081 8988 10137 9044
rect 10223 8988 10279 9044
rect 10081 8846 10137 8902
rect 10223 8846 10279 8902
rect 10081 8704 10137 8760
rect 10223 8704 10279 8760
rect 10081 8562 10137 8618
rect 10223 8562 10279 8618
rect 10081 8420 10137 8476
rect 10223 8420 10279 8476
rect 10081 8278 10137 8334
rect 10223 8278 10279 8334
rect 10081 8136 10137 8192
rect 10223 8136 10279 8192
rect 10081 7994 10137 8050
rect 10223 7994 10279 8050
rect 10081 7852 10137 7908
rect 10223 7852 10279 7908
rect 10081 7710 10137 7766
rect 10223 7710 10279 7766
rect 10081 7568 10137 7624
rect 10223 7568 10279 7624
rect 10081 7426 10137 7482
rect 10223 7426 10279 7482
rect 10081 7284 10137 7340
rect 10223 7284 10279 7340
rect 10081 7142 10137 7198
rect 10223 7142 10279 7198
rect 10081 7000 10137 7056
rect 10223 7000 10279 7056
rect 10081 6858 10137 6914
rect 10223 6858 10279 6914
rect 10081 6716 10137 6772
rect 10223 6716 10279 6772
rect 10081 6574 10137 6630
rect 10223 6574 10279 6630
rect 10081 6432 10137 6488
rect 10223 6432 10279 6488
rect 10081 6290 10137 6346
rect 10223 6290 10279 6346
rect 10081 6148 10137 6204
rect 10223 6148 10279 6204
rect 10081 6006 10137 6062
rect 10223 6006 10279 6062
rect 10081 5864 10137 5920
rect 10223 5864 10279 5920
rect 10081 5722 10137 5778
rect 10223 5722 10279 5778
rect 10081 5580 10137 5636
rect 10223 5580 10279 5636
rect 10081 5438 10137 5494
rect 10223 5438 10279 5494
rect 10081 5296 10137 5352
rect 10223 5296 10279 5352
rect 10081 5154 10137 5210
rect 10223 5154 10279 5210
rect 10081 5012 10137 5068
rect 10223 5012 10279 5068
rect 10081 4870 10137 4926
rect 10223 4870 10279 4926
rect 10081 4728 10137 4784
rect 10223 4728 10279 4784
rect 10081 4586 10137 4642
rect 10223 4586 10279 4642
rect 10081 4444 10137 4500
rect 10223 4444 10279 4500
rect 10081 4302 10137 4358
rect 10223 4302 10279 4358
rect 10081 4160 10137 4216
rect 10223 4160 10279 4216
rect 10081 4018 10137 4074
rect 10223 4018 10279 4074
rect 10081 3876 10137 3932
rect 10223 3876 10279 3932
rect 10081 3734 10137 3790
rect 10223 3734 10279 3790
rect 10081 3592 10137 3648
rect 10223 3592 10279 3648
rect 10081 3450 10137 3506
rect 10223 3450 10279 3506
rect 10081 3308 10137 3364
rect 10223 3308 10279 3364
rect 10081 3166 10137 3222
rect 10223 3166 10279 3222
rect 10081 3024 10137 3080
rect 10223 3024 10279 3080
rect 10081 2882 10137 2938
rect 10223 2882 10279 2938
rect 10081 2740 10137 2796
rect 10223 2740 10279 2796
rect 10081 2598 10137 2654
rect 10223 2598 10279 2654
rect 10081 2456 10137 2512
rect 10223 2456 10279 2512
rect 10081 2314 10137 2370
rect 10223 2314 10279 2370
rect 10081 2172 10137 2228
rect 10223 2172 10279 2228
rect 10081 2030 10137 2086
rect 10223 2030 10279 2086
rect 10081 1888 10137 1944
rect 10223 1888 10279 1944
rect 10081 1746 10137 1802
rect 10223 1746 10279 1802
rect 10081 1604 10137 1660
rect 10223 1604 10279 1660
rect 10081 1462 10137 1518
rect 10223 1462 10279 1518
rect 10081 1320 10137 1376
rect 10223 1320 10279 1376
rect 10081 1178 10137 1234
rect 10223 1178 10279 1234
rect 10081 1036 10137 1092
rect 10223 1036 10279 1092
rect 10081 894 10137 950
rect 10223 894 10279 950
rect 10081 752 10137 808
rect 10223 752 10279 808
rect 10081 610 10137 666
rect 10223 610 10279 666
rect 10081 468 10137 524
rect 10223 468 10279 524
rect 10622 12254 10678 12310
rect 10764 12254 10820 12310
rect 10622 12112 10678 12168
rect 10764 12112 10820 12168
rect 10622 11970 10678 12026
rect 10764 11970 10820 12026
rect 10622 11828 10678 11884
rect 10764 11828 10820 11884
rect 10622 11686 10678 11742
rect 10764 11686 10820 11742
rect 10622 11544 10678 11600
rect 10764 11544 10820 11600
rect 10622 11402 10678 11458
rect 10764 11402 10820 11458
rect 10622 11260 10678 11316
rect 10764 11260 10820 11316
rect 10622 11118 10678 11174
rect 10764 11118 10820 11174
rect 10622 10976 10678 11032
rect 10764 10976 10820 11032
rect 10622 10834 10678 10890
rect 10764 10834 10820 10890
rect 10622 10692 10678 10748
rect 10764 10692 10820 10748
rect 10622 10550 10678 10606
rect 10764 10550 10820 10606
rect 10622 10408 10678 10464
rect 10764 10408 10820 10464
rect 10622 10266 10678 10322
rect 10764 10266 10820 10322
rect 10622 10124 10678 10180
rect 10764 10124 10820 10180
rect 10622 9982 10678 10038
rect 10764 9982 10820 10038
rect 10622 9840 10678 9896
rect 10764 9840 10820 9896
rect 10622 9698 10678 9754
rect 10764 9698 10820 9754
rect 10622 9556 10678 9612
rect 10764 9556 10820 9612
rect 10622 9414 10678 9470
rect 10764 9414 10820 9470
rect 10622 9272 10678 9328
rect 10764 9272 10820 9328
rect 10622 9130 10678 9186
rect 10764 9130 10820 9186
rect 10622 8988 10678 9044
rect 10764 8988 10820 9044
rect 10622 8846 10678 8902
rect 10764 8846 10820 8902
rect 10622 8704 10678 8760
rect 10764 8704 10820 8760
rect 10622 8562 10678 8618
rect 10764 8562 10820 8618
rect 10622 8420 10678 8476
rect 10764 8420 10820 8476
rect 10622 8278 10678 8334
rect 10764 8278 10820 8334
rect 10622 8136 10678 8192
rect 10764 8136 10820 8192
rect 10622 7994 10678 8050
rect 10764 7994 10820 8050
rect 10622 7852 10678 7908
rect 10764 7852 10820 7908
rect 10622 7710 10678 7766
rect 10764 7710 10820 7766
rect 10622 7568 10678 7624
rect 10764 7568 10820 7624
rect 10622 7426 10678 7482
rect 10764 7426 10820 7482
rect 10622 7284 10678 7340
rect 10764 7284 10820 7340
rect 10622 7142 10678 7198
rect 10764 7142 10820 7198
rect 10622 7000 10678 7056
rect 10764 7000 10820 7056
rect 10622 6858 10678 6914
rect 10764 6858 10820 6914
rect 10622 6716 10678 6772
rect 10764 6716 10820 6772
rect 10622 6574 10678 6630
rect 10764 6574 10820 6630
rect 10622 6432 10678 6488
rect 10764 6432 10820 6488
rect 10622 6290 10678 6346
rect 10764 6290 10820 6346
rect 10622 6148 10678 6204
rect 10764 6148 10820 6204
rect 10622 6006 10678 6062
rect 10764 6006 10820 6062
rect 10622 5864 10678 5920
rect 10764 5864 10820 5920
rect 10622 5722 10678 5778
rect 10764 5722 10820 5778
rect 10622 5580 10678 5636
rect 10764 5580 10820 5636
rect 10622 5438 10678 5494
rect 10764 5438 10820 5494
rect 10622 5296 10678 5352
rect 10764 5296 10820 5352
rect 10622 5154 10678 5210
rect 10764 5154 10820 5210
rect 10622 5012 10678 5068
rect 10764 5012 10820 5068
rect 10622 4870 10678 4926
rect 10764 4870 10820 4926
rect 10622 4728 10678 4784
rect 10764 4728 10820 4784
rect 10622 4586 10678 4642
rect 10764 4586 10820 4642
rect 10622 4444 10678 4500
rect 10764 4444 10820 4500
rect 10622 4302 10678 4358
rect 10764 4302 10820 4358
rect 10622 4160 10678 4216
rect 10764 4160 10820 4216
rect 10622 4018 10678 4074
rect 10764 4018 10820 4074
rect 10622 3876 10678 3932
rect 10764 3876 10820 3932
rect 10622 3734 10678 3790
rect 10764 3734 10820 3790
rect 10622 3592 10678 3648
rect 10764 3592 10820 3648
rect 10622 3450 10678 3506
rect 10764 3450 10820 3506
rect 10622 3308 10678 3364
rect 10764 3308 10820 3364
rect 10622 3166 10678 3222
rect 10764 3166 10820 3222
rect 10622 3024 10678 3080
rect 10764 3024 10820 3080
rect 10622 2882 10678 2938
rect 10764 2882 10820 2938
rect 10622 2740 10678 2796
rect 10764 2740 10820 2796
rect 10622 2598 10678 2654
rect 10764 2598 10820 2654
rect 10622 2456 10678 2512
rect 10764 2456 10820 2512
rect 10622 2314 10678 2370
rect 10764 2314 10820 2370
rect 10622 2172 10678 2228
rect 10764 2172 10820 2228
rect 10622 2030 10678 2086
rect 10764 2030 10820 2086
rect 10622 1888 10678 1944
rect 10764 1888 10820 1944
rect 10622 1746 10678 1802
rect 10764 1746 10820 1802
rect 10622 1604 10678 1660
rect 10764 1604 10820 1660
rect 10622 1462 10678 1518
rect 10764 1462 10820 1518
rect 10622 1320 10678 1376
rect 10764 1320 10820 1376
rect 10622 1178 10678 1234
rect 10764 1178 10820 1234
rect 10622 1036 10678 1092
rect 10764 1036 10820 1092
rect 10622 894 10678 950
rect 10764 894 10820 950
rect 10622 752 10678 808
rect 10764 752 10820 808
rect 10622 610 10678 666
rect 10764 610 10820 666
rect 10622 468 10678 524
rect 10764 468 10820 524
rect 11162 12254 11218 12310
rect 11304 12254 11360 12310
rect 11162 12112 11218 12168
rect 11304 12112 11360 12168
rect 11162 11970 11218 12026
rect 11304 11970 11360 12026
rect 11162 11828 11218 11884
rect 11304 11828 11360 11884
rect 11162 11686 11218 11742
rect 11304 11686 11360 11742
rect 11162 11544 11218 11600
rect 11304 11544 11360 11600
rect 11162 11402 11218 11458
rect 11304 11402 11360 11458
rect 11162 11260 11218 11316
rect 11304 11260 11360 11316
rect 11162 11118 11218 11174
rect 11304 11118 11360 11174
rect 11162 10976 11218 11032
rect 11304 10976 11360 11032
rect 11162 10834 11218 10890
rect 11304 10834 11360 10890
rect 11162 10692 11218 10748
rect 11304 10692 11360 10748
rect 11162 10550 11218 10606
rect 11304 10550 11360 10606
rect 11162 10408 11218 10464
rect 11304 10408 11360 10464
rect 11162 10266 11218 10322
rect 11304 10266 11360 10322
rect 11162 10124 11218 10180
rect 11304 10124 11360 10180
rect 11162 9982 11218 10038
rect 11304 9982 11360 10038
rect 11162 9840 11218 9896
rect 11304 9840 11360 9896
rect 11162 9698 11218 9754
rect 11304 9698 11360 9754
rect 11162 9556 11218 9612
rect 11304 9556 11360 9612
rect 11162 9414 11218 9470
rect 11304 9414 11360 9470
rect 11162 9272 11218 9328
rect 11304 9272 11360 9328
rect 11162 9130 11218 9186
rect 11304 9130 11360 9186
rect 11162 8988 11218 9044
rect 11304 8988 11360 9044
rect 11162 8846 11218 8902
rect 11304 8846 11360 8902
rect 11162 8704 11218 8760
rect 11304 8704 11360 8760
rect 11162 8562 11218 8618
rect 11304 8562 11360 8618
rect 11162 8420 11218 8476
rect 11304 8420 11360 8476
rect 11162 8278 11218 8334
rect 11304 8278 11360 8334
rect 11162 8136 11218 8192
rect 11304 8136 11360 8192
rect 11162 7994 11218 8050
rect 11304 7994 11360 8050
rect 11162 7852 11218 7908
rect 11304 7852 11360 7908
rect 11162 7710 11218 7766
rect 11304 7710 11360 7766
rect 11162 7568 11218 7624
rect 11304 7568 11360 7624
rect 11162 7426 11218 7482
rect 11304 7426 11360 7482
rect 11162 7284 11218 7340
rect 11304 7284 11360 7340
rect 11162 7142 11218 7198
rect 11304 7142 11360 7198
rect 11162 7000 11218 7056
rect 11304 7000 11360 7056
rect 11162 6858 11218 6914
rect 11304 6858 11360 6914
rect 11162 6716 11218 6772
rect 11304 6716 11360 6772
rect 11162 6574 11218 6630
rect 11304 6574 11360 6630
rect 11162 6432 11218 6488
rect 11304 6432 11360 6488
rect 11162 6290 11218 6346
rect 11304 6290 11360 6346
rect 11162 6148 11218 6204
rect 11304 6148 11360 6204
rect 11162 6006 11218 6062
rect 11304 6006 11360 6062
rect 11162 5864 11218 5920
rect 11304 5864 11360 5920
rect 11162 5722 11218 5778
rect 11304 5722 11360 5778
rect 11162 5580 11218 5636
rect 11304 5580 11360 5636
rect 11162 5438 11218 5494
rect 11304 5438 11360 5494
rect 11162 5296 11218 5352
rect 11304 5296 11360 5352
rect 11162 5154 11218 5210
rect 11304 5154 11360 5210
rect 11162 5012 11218 5068
rect 11304 5012 11360 5068
rect 11162 4870 11218 4926
rect 11304 4870 11360 4926
rect 11162 4728 11218 4784
rect 11304 4728 11360 4784
rect 11162 4586 11218 4642
rect 11304 4586 11360 4642
rect 11162 4444 11218 4500
rect 11304 4444 11360 4500
rect 11162 4302 11218 4358
rect 11304 4302 11360 4358
rect 11162 4160 11218 4216
rect 11304 4160 11360 4216
rect 11162 4018 11218 4074
rect 11304 4018 11360 4074
rect 11162 3876 11218 3932
rect 11304 3876 11360 3932
rect 11162 3734 11218 3790
rect 11304 3734 11360 3790
rect 11162 3592 11218 3648
rect 11304 3592 11360 3648
rect 11162 3450 11218 3506
rect 11304 3450 11360 3506
rect 11162 3308 11218 3364
rect 11304 3308 11360 3364
rect 11162 3166 11218 3222
rect 11304 3166 11360 3222
rect 11162 3024 11218 3080
rect 11304 3024 11360 3080
rect 11162 2882 11218 2938
rect 11304 2882 11360 2938
rect 11162 2740 11218 2796
rect 11304 2740 11360 2796
rect 11162 2598 11218 2654
rect 11304 2598 11360 2654
rect 11162 2456 11218 2512
rect 11304 2456 11360 2512
rect 11162 2314 11218 2370
rect 11304 2314 11360 2370
rect 11162 2172 11218 2228
rect 11304 2172 11360 2228
rect 11162 2030 11218 2086
rect 11304 2030 11360 2086
rect 11162 1888 11218 1944
rect 11304 1888 11360 1944
rect 11162 1746 11218 1802
rect 11304 1746 11360 1802
rect 11162 1604 11218 1660
rect 11304 1604 11360 1660
rect 11162 1462 11218 1518
rect 11304 1462 11360 1518
rect 11162 1320 11218 1376
rect 11304 1320 11360 1376
rect 11162 1178 11218 1234
rect 11304 1178 11360 1234
rect 11162 1036 11218 1092
rect 11304 1036 11360 1092
rect 11162 894 11218 950
rect 11304 894 11360 950
rect 11162 752 11218 808
rect 11304 752 11360 808
rect 11162 610 11218 666
rect 11304 610 11360 666
rect 11162 468 11218 524
rect 11304 468 11360 524
rect 11702 12254 11758 12310
rect 11844 12254 11900 12310
rect 11702 12112 11758 12168
rect 11844 12112 11900 12168
rect 11702 11970 11758 12026
rect 11844 11970 11900 12026
rect 11702 11828 11758 11884
rect 11844 11828 11900 11884
rect 11702 11686 11758 11742
rect 11844 11686 11900 11742
rect 11702 11544 11758 11600
rect 11844 11544 11900 11600
rect 11702 11402 11758 11458
rect 11844 11402 11900 11458
rect 11702 11260 11758 11316
rect 11844 11260 11900 11316
rect 11702 11118 11758 11174
rect 11844 11118 11900 11174
rect 11702 10976 11758 11032
rect 11844 10976 11900 11032
rect 11702 10834 11758 10890
rect 11844 10834 11900 10890
rect 11702 10692 11758 10748
rect 11844 10692 11900 10748
rect 11702 10550 11758 10606
rect 11844 10550 11900 10606
rect 11702 10408 11758 10464
rect 11844 10408 11900 10464
rect 11702 10266 11758 10322
rect 11844 10266 11900 10322
rect 11702 10124 11758 10180
rect 11844 10124 11900 10180
rect 11702 9982 11758 10038
rect 11844 9982 11900 10038
rect 11702 9840 11758 9896
rect 11844 9840 11900 9896
rect 11702 9698 11758 9754
rect 11844 9698 11900 9754
rect 11702 9556 11758 9612
rect 11844 9556 11900 9612
rect 11702 9414 11758 9470
rect 11844 9414 11900 9470
rect 11702 9272 11758 9328
rect 11844 9272 11900 9328
rect 11702 9130 11758 9186
rect 11844 9130 11900 9186
rect 11702 8988 11758 9044
rect 11844 8988 11900 9044
rect 11702 8846 11758 8902
rect 11844 8846 11900 8902
rect 11702 8704 11758 8760
rect 11844 8704 11900 8760
rect 11702 8562 11758 8618
rect 11844 8562 11900 8618
rect 11702 8420 11758 8476
rect 11844 8420 11900 8476
rect 11702 8278 11758 8334
rect 11844 8278 11900 8334
rect 11702 8136 11758 8192
rect 11844 8136 11900 8192
rect 11702 7994 11758 8050
rect 11844 7994 11900 8050
rect 11702 7852 11758 7908
rect 11844 7852 11900 7908
rect 11702 7710 11758 7766
rect 11844 7710 11900 7766
rect 11702 7568 11758 7624
rect 11844 7568 11900 7624
rect 11702 7426 11758 7482
rect 11844 7426 11900 7482
rect 11702 7284 11758 7340
rect 11844 7284 11900 7340
rect 11702 7142 11758 7198
rect 11844 7142 11900 7198
rect 11702 7000 11758 7056
rect 11844 7000 11900 7056
rect 11702 6858 11758 6914
rect 11844 6858 11900 6914
rect 11702 6716 11758 6772
rect 11844 6716 11900 6772
rect 11702 6574 11758 6630
rect 11844 6574 11900 6630
rect 11702 6432 11758 6488
rect 11844 6432 11900 6488
rect 11702 6290 11758 6346
rect 11844 6290 11900 6346
rect 11702 6148 11758 6204
rect 11844 6148 11900 6204
rect 11702 6006 11758 6062
rect 11844 6006 11900 6062
rect 11702 5864 11758 5920
rect 11844 5864 11900 5920
rect 11702 5722 11758 5778
rect 11844 5722 11900 5778
rect 11702 5580 11758 5636
rect 11844 5580 11900 5636
rect 11702 5438 11758 5494
rect 11844 5438 11900 5494
rect 11702 5296 11758 5352
rect 11844 5296 11900 5352
rect 11702 5154 11758 5210
rect 11844 5154 11900 5210
rect 11702 5012 11758 5068
rect 11844 5012 11900 5068
rect 11702 4870 11758 4926
rect 11844 4870 11900 4926
rect 11702 4728 11758 4784
rect 11844 4728 11900 4784
rect 11702 4586 11758 4642
rect 11844 4586 11900 4642
rect 11702 4444 11758 4500
rect 11844 4444 11900 4500
rect 11702 4302 11758 4358
rect 11844 4302 11900 4358
rect 11702 4160 11758 4216
rect 11844 4160 11900 4216
rect 11702 4018 11758 4074
rect 11844 4018 11900 4074
rect 11702 3876 11758 3932
rect 11844 3876 11900 3932
rect 11702 3734 11758 3790
rect 11844 3734 11900 3790
rect 11702 3592 11758 3648
rect 11844 3592 11900 3648
rect 11702 3450 11758 3506
rect 11844 3450 11900 3506
rect 11702 3308 11758 3364
rect 11844 3308 11900 3364
rect 11702 3166 11758 3222
rect 11844 3166 11900 3222
rect 11702 3024 11758 3080
rect 11844 3024 11900 3080
rect 11702 2882 11758 2938
rect 11844 2882 11900 2938
rect 11702 2740 11758 2796
rect 11844 2740 11900 2796
rect 11702 2598 11758 2654
rect 11844 2598 11900 2654
rect 11702 2456 11758 2512
rect 11844 2456 11900 2512
rect 11702 2314 11758 2370
rect 11844 2314 11900 2370
rect 11702 2172 11758 2228
rect 11844 2172 11900 2228
rect 11702 2030 11758 2086
rect 11844 2030 11900 2086
rect 11702 1888 11758 1944
rect 11844 1888 11900 1944
rect 11702 1746 11758 1802
rect 11844 1746 11900 1802
rect 11702 1604 11758 1660
rect 11844 1604 11900 1660
rect 11702 1462 11758 1518
rect 11844 1462 11900 1518
rect 11702 1320 11758 1376
rect 11844 1320 11900 1376
rect 11702 1178 11758 1234
rect 11844 1178 11900 1234
rect 11702 1036 11758 1092
rect 11844 1036 11900 1092
rect 11702 894 11758 950
rect 11844 894 11900 950
rect 11702 752 11758 808
rect 11844 752 11900 808
rect 11702 610 11758 666
rect 11844 610 11900 666
rect 11702 468 11758 524
rect 11844 468 11900 524
rect 12526 12302 12582 12358
rect 12650 12302 12706 12358
rect 12774 12302 12830 12358
rect 12898 12302 12954 12358
rect 13022 12302 13078 12358
rect 12526 12178 12582 12234
rect 12650 12178 12706 12234
rect 12774 12178 12830 12234
rect 12898 12178 12954 12234
rect 13022 12178 13078 12234
rect 12526 12054 12582 12110
rect 12650 12054 12706 12110
rect 12774 12054 12830 12110
rect 12898 12054 12954 12110
rect 13022 12054 13078 12110
rect 12526 11930 12582 11986
rect 12650 11930 12706 11986
rect 12774 11930 12830 11986
rect 12898 11930 12954 11986
rect 13022 11930 13078 11986
rect 12526 11806 12582 11862
rect 12650 11806 12706 11862
rect 12774 11806 12830 11862
rect 12898 11806 12954 11862
rect 13022 11806 13078 11862
rect 12526 11682 12582 11738
rect 12650 11682 12706 11738
rect 12774 11682 12830 11738
rect 12898 11682 12954 11738
rect 13022 11682 13078 11738
rect 12526 11558 12582 11614
rect 12650 11558 12706 11614
rect 12774 11558 12830 11614
rect 12898 11558 12954 11614
rect 13022 11558 13078 11614
rect 12526 11434 12582 11490
rect 12650 11434 12706 11490
rect 12774 11434 12830 11490
rect 12898 11434 12954 11490
rect 13022 11434 13078 11490
rect 12526 11310 12582 11366
rect 12650 11310 12706 11366
rect 12774 11310 12830 11366
rect 12898 11310 12954 11366
rect 13022 11310 13078 11366
rect 12526 11186 12582 11242
rect 12650 11186 12706 11242
rect 12774 11186 12830 11242
rect 12898 11186 12954 11242
rect 13022 11186 13078 11242
rect 12526 11062 12582 11118
rect 12650 11062 12706 11118
rect 12774 11062 12830 11118
rect 12898 11062 12954 11118
rect 13022 11062 13078 11118
rect 12526 10938 12582 10994
rect 12650 10938 12706 10994
rect 12774 10938 12830 10994
rect 12898 10938 12954 10994
rect 13022 10938 13078 10994
rect 12526 10814 12582 10870
rect 12650 10814 12706 10870
rect 12774 10814 12830 10870
rect 12898 10814 12954 10870
rect 13022 10814 13078 10870
rect 12526 10690 12582 10746
rect 12650 10690 12706 10746
rect 12774 10690 12830 10746
rect 12898 10690 12954 10746
rect 13022 10690 13078 10746
rect 12526 10566 12582 10622
rect 12650 10566 12706 10622
rect 12774 10566 12830 10622
rect 12898 10566 12954 10622
rect 13022 10566 13078 10622
rect 12526 10442 12582 10498
rect 12650 10442 12706 10498
rect 12774 10442 12830 10498
rect 12898 10442 12954 10498
rect 13022 10442 13078 10498
rect 12526 10318 12582 10374
rect 12650 10318 12706 10374
rect 12774 10318 12830 10374
rect 12898 10318 12954 10374
rect 13022 10318 13078 10374
rect 12526 10194 12582 10250
rect 12650 10194 12706 10250
rect 12774 10194 12830 10250
rect 12898 10194 12954 10250
rect 13022 10194 13078 10250
rect 12526 10070 12582 10126
rect 12650 10070 12706 10126
rect 12774 10070 12830 10126
rect 12898 10070 12954 10126
rect 13022 10070 13078 10126
rect 12526 9946 12582 10002
rect 12650 9946 12706 10002
rect 12774 9946 12830 10002
rect 12898 9946 12954 10002
rect 13022 9946 13078 10002
rect 12526 9822 12582 9878
rect 12650 9822 12706 9878
rect 12774 9822 12830 9878
rect 12898 9822 12954 9878
rect 13022 9822 13078 9878
rect 12526 9698 12582 9754
rect 12650 9698 12706 9754
rect 12774 9698 12830 9754
rect 12898 9698 12954 9754
rect 13022 9698 13078 9754
rect 12526 9574 12582 9630
rect 12650 9574 12706 9630
rect 12774 9574 12830 9630
rect 12898 9574 12954 9630
rect 13022 9574 13078 9630
rect 12526 9450 12582 9506
rect 12650 9450 12706 9506
rect 12774 9450 12830 9506
rect 12898 9450 12954 9506
rect 13022 9450 13078 9506
rect 12526 9326 12582 9382
rect 12650 9326 12706 9382
rect 12774 9326 12830 9382
rect 12898 9326 12954 9382
rect 13022 9326 13078 9382
rect 12526 9202 12582 9258
rect 12650 9202 12706 9258
rect 12774 9202 12830 9258
rect 12898 9202 12954 9258
rect 13022 9202 13078 9258
rect 12526 9078 12582 9134
rect 12650 9078 12706 9134
rect 12774 9078 12830 9134
rect 12898 9078 12954 9134
rect 13022 9078 13078 9134
rect 12526 8954 12582 9010
rect 12650 8954 12706 9010
rect 12774 8954 12830 9010
rect 12898 8954 12954 9010
rect 13022 8954 13078 9010
rect 12526 8830 12582 8886
rect 12650 8830 12706 8886
rect 12774 8830 12830 8886
rect 12898 8830 12954 8886
rect 13022 8830 13078 8886
rect 12526 8706 12582 8762
rect 12650 8706 12706 8762
rect 12774 8706 12830 8762
rect 12898 8706 12954 8762
rect 13022 8706 13078 8762
rect 12526 8582 12582 8638
rect 12650 8582 12706 8638
rect 12774 8582 12830 8638
rect 12898 8582 12954 8638
rect 13022 8582 13078 8638
rect 12526 8458 12582 8514
rect 12650 8458 12706 8514
rect 12774 8458 12830 8514
rect 12898 8458 12954 8514
rect 13022 8458 13078 8514
rect 12526 8334 12582 8390
rect 12650 8334 12706 8390
rect 12774 8334 12830 8390
rect 12898 8334 12954 8390
rect 13022 8334 13078 8390
rect 12526 8210 12582 8266
rect 12650 8210 12706 8266
rect 12774 8210 12830 8266
rect 12898 8210 12954 8266
rect 13022 8210 13078 8266
rect 12526 8086 12582 8142
rect 12650 8086 12706 8142
rect 12774 8086 12830 8142
rect 12898 8086 12954 8142
rect 13022 8086 13078 8142
rect 12526 7962 12582 8018
rect 12650 7962 12706 8018
rect 12774 7962 12830 8018
rect 12898 7962 12954 8018
rect 13022 7962 13078 8018
rect 12526 7838 12582 7894
rect 12650 7838 12706 7894
rect 12774 7838 12830 7894
rect 12898 7838 12954 7894
rect 13022 7838 13078 7894
rect 12526 7714 12582 7770
rect 12650 7714 12706 7770
rect 12774 7714 12830 7770
rect 12898 7714 12954 7770
rect 13022 7714 13078 7770
rect 12526 7590 12582 7646
rect 12650 7590 12706 7646
rect 12774 7590 12830 7646
rect 12898 7590 12954 7646
rect 13022 7590 13078 7646
rect 12526 7466 12582 7522
rect 12650 7466 12706 7522
rect 12774 7466 12830 7522
rect 12898 7466 12954 7522
rect 13022 7466 13078 7522
rect 12526 7342 12582 7398
rect 12650 7342 12706 7398
rect 12774 7342 12830 7398
rect 12898 7342 12954 7398
rect 13022 7342 13078 7398
rect 12526 7218 12582 7274
rect 12650 7218 12706 7274
rect 12774 7218 12830 7274
rect 12898 7218 12954 7274
rect 13022 7218 13078 7274
rect 12526 7094 12582 7150
rect 12650 7094 12706 7150
rect 12774 7094 12830 7150
rect 12898 7094 12954 7150
rect 13022 7094 13078 7150
rect 12526 6970 12582 7026
rect 12650 6970 12706 7026
rect 12774 6970 12830 7026
rect 12898 6970 12954 7026
rect 13022 6970 13078 7026
rect 12526 6846 12582 6902
rect 12650 6846 12706 6902
rect 12774 6846 12830 6902
rect 12898 6846 12954 6902
rect 13022 6846 13078 6902
rect 12526 6722 12582 6778
rect 12650 6722 12706 6778
rect 12774 6722 12830 6778
rect 12898 6722 12954 6778
rect 13022 6722 13078 6778
rect 12526 6598 12582 6654
rect 12650 6598 12706 6654
rect 12774 6598 12830 6654
rect 12898 6598 12954 6654
rect 13022 6598 13078 6654
rect 12526 6474 12582 6530
rect 12650 6474 12706 6530
rect 12774 6474 12830 6530
rect 12898 6474 12954 6530
rect 13022 6474 13078 6530
rect 12526 6350 12582 6406
rect 12650 6350 12706 6406
rect 12774 6350 12830 6406
rect 12898 6350 12954 6406
rect 13022 6350 13078 6406
rect 12526 6226 12582 6282
rect 12650 6226 12706 6282
rect 12774 6226 12830 6282
rect 12898 6226 12954 6282
rect 13022 6226 13078 6282
rect 12526 6102 12582 6158
rect 12650 6102 12706 6158
rect 12774 6102 12830 6158
rect 12898 6102 12954 6158
rect 13022 6102 13078 6158
rect 12526 5978 12582 6034
rect 12650 5978 12706 6034
rect 12774 5978 12830 6034
rect 12898 5978 12954 6034
rect 13022 5978 13078 6034
rect 12526 5854 12582 5910
rect 12650 5854 12706 5910
rect 12774 5854 12830 5910
rect 12898 5854 12954 5910
rect 13022 5854 13078 5910
rect 12526 5730 12582 5786
rect 12650 5730 12706 5786
rect 12774 5730 12830 5786
rect 12898 5730 12954 5786
rect 13022 5730 13078 5786
rect 12526 5606 12582 5662
rect 12650 5606 12706 5662
rect 12774 5606 12830 5662
rect 12898 5606 12954 5662
rect 13022 5606 13078 5662
rect 12526 5482 12582 5538
rect 12650 5482 12706 5538
rect 12774 5482 12830 5538
rect 12898 5482 12954 5538
rect 13022 5482 13078 5538
rect 12526 5358 12582 5414
rect 12650 5358 12706 5414
rect 12774 5358 12830 5414
rect 12898 5358 12954 5414
rect 13022 5358 13078 5414
rect 12526 5234 12582 5290
rect 12650 5234 12706 5290
rect 12774 5234 12830 5290
rect 12898 5234 12954 5290
rect 13022 5234 13078 5290
rect 12526 5110 12582 5166
rect 12650 5110 12706 5166
rect 12774 5110 12830 5166
rect 12898 5110 12954 5166
rect 13022 5110 13078 5166
rect 12526 4986 12582 5042
rect 12650 4986 12706 5042
rect 12774 4986 12830 5042
rect 12898 4986 12954 5042
rect 13022 4986 13078 5042
rect 12526 4862 12582 4918
rect 12650 4862 12706 4918
rect 12774 4862 12830 4918
rect 12898 4862 12954 4918
rect 13022 4862 13078 4918
rect 12526 4738 12582 4794
rect 12650 4738 12706 4794
rect 12774 4738 12830 4794
rect 12898 4738 12954 4794
rect 13022 4738 13078 4794
rect 12526 4614 12582 4670
rect 12650 4614 12706 4670
rect 12774 4614 12830 4670
rect 12898 4614 12954 4670
rect 13022 4614 13078 4670
rect 12526 4490 12582 4546
rect 12650 4490 12706 4546
rect 12774 4490 12830 4546
rect 12898 4490 12954 4546
rect 13022 4490 13078 4546
rect 12526 4366 12582 4422
rect 12650 4366 12706 4422
rect 12774 4366 12830 4422
rect 12898 4366 12954 4422
rect 13022 4366 13078 4422
rect 12526 4242 12582 4298
rect 12650 4242 12706 4298
rect 12774 4242 12830 4298
rect 12898 4242 12954 4298
rect 13022 4242 13078 4298
rect 12526 4118 12582 4174
rect 12650 4118 12706 4174
rect 12774 4118 12830 4174
rect 12898 4118 12954 4174
rect 13022 4118 13078 4174
rect 12526 3994 12582 4050
rect 12650 3994 12706 4050
rect 12774 3994 12830 4050
rect 12898 3994 12954 4050
rect 13022 3994 13078 4050
rect 12526 3870 12582 3926
rect 12650 3870 12706 3926
rect 12774 3870 12830 3926
rect 12898 3870 12954 3926
rect 13022 3870 13078 3926
rect 12526 3746 12582 3802
rect 12650 3746 12706 3802
rect 12774 3746 12830 3802
rect 12898 3746 12954 3802
rect 13022 3746 13078 3802
rect 12526 3622 12582 3678
rect 12650 3622 12706 3678
rect 12774 3622 12830 3678
rect 12898 3622 12954 3678
rect 13022 3622 13078 3678
rect 12526 3498 12582 3554
rect 12650 3498 12706 3554
rect 12774 3498 12830 3554
rect 12898 3498 12954 3554
rect 13022 3498 13078 3554
rect 12526 3374 12582 3430
rect 12650 3374 12706 3430
rect 12774 3374 12830 3430
rect 12898 3374 12954 3430
rect 13022 3374 13078 3430
rect 12526 3250 12582 3306
rect 12650 3250 12706 3306
rect 12774 3250 12830 3306
rect 12898 3250 12954 3306
rect 13022 3250 13078 3306
rect 12526 3126 12582 3182
rect 12650 3126 12706 3182
rect 12774 3126 12830 3182
rect 12898 3126 12954 3182
rect 13022 3126 13078 3182
rect 12526 3002 12582 3058
rect 12650 3002 12706 3058
rect 12774 3002 12830 3058
rect 12898 3002 12954 3058
rect 13022 3002 13078 3058
rect 12526 2878 12582 2934
rect 12650 2878 12706 2934
rect 12774 2878 12830 2934
rect 12898 2878 12954 2934
rect 13022 2878 13078 2934
rect 12526 2754 12582 2810
rect 12650 2754 12706 2810
rect 12774 2754 12830 2810
rect 12898 2754 12954 2810
rect 13022 2754 13078 2810
rect 12526 2630 12582 2686
rect 12650 2630 12706 2686
rect 12774 2630 12830 2686
rect 12898 2630 12954 2686
rect 13022 2630 13078 2686
rect 12526 2506 12582 2562
rect 12650 2506 12706 2562
rect 12774 2506 12830 2562
rect 12898 2506 12954 2562
rect 13022 2506 13078 2562
rect 12526 2382 12582 2438
rect 12650 2382 12706 2438
rect 12774 2382 12830 2438
rect 12898 2382 12954 2438
rect 13022 2382 13078 2438
rect 12526 2258 12582 2314
rect 12650 2258 12706 2314
rect 12774 2258 12830 2314
rect 12898 2258 12954 2314
rect 13022 2258 13078 2314
rect 12526 2134 12582 2190
rect 12650 2134 12706 2190
rect 12774 2134 12830 2190
rect 12898 2134 12954 2190
rect 13022 2134 13078 2190
rect 12526 2010 12582 2066
rect 12650 2010 12706 2066
rect 12774 2010 12830 2066
rect 12898 2010 12954 2066
rect 13022 2010 13078 2066
rect 12526 1886 12582 1942
rect 12650 1886 12706 1942
rect 12774 1886 12830 1942
rect 12898 1886 12954 1942
rect 13022 1886 13078 1942
rect 12526 1762 12582 1818
rect 12650 1762 12706 1818
rect 12774 1762 12830 1818
rect 12898 1762 12954 1818
rect 13022 1762 13078 1818
rect 12526 1638 12582 1694
rect 12650 1638 12706 1694
rect 12774 1638 12830 1694
rect 12898 1638 12954 1694
rect 13022 1638 13078 1694
rect 12526 1514 12582 1570
rect 12650 1514 12706 1570
rect 12774 1514 12830 1570
rect 12898 1514 12954 1570
rect 13022 1514 13078 1570
rect 12526 1390 12582 1446
rect 12650 1390 12706 1446
rect 12774 1390 12830 1446
rect 12898 1390 12954 1446
rect 13022 1390 13078 1446
rect 12526 1266 12582 1322
rect 12650 1266 12706 1322
rect 12774 1266 12830 1322
rect 12898 1266 12954 1322
rect 13022 1266 13078 1322
rect 12526 1142 12582 1198
rect 12650 1142 12706 1198
rect 12774 1142 12830 1198
rect 12898 1142 12954 1198
rect 13022 1142 13078 1198
rect 12526 1018 12582 1074
rect 12650 1018 12706 1074
rect 12774 1018 12830 1074
rect 12898 1018 12954 1074
rect 13022 1018 13078 1074
rect 12526 894 12582 950
rect 12650 894 12706 950
rect 12774 894 12830 950
rect 12898 894 12954 950
rect 13022 894 13078 950
rect 12526 770 12582 826
rect 12650 770 12706 826
rect 12774 770 12830 826
rect 12898 770 12954 826
rect 13022 770 13078 826
rect 12526 646 12582 702
rect 12650 646 12706 702
rect 12774 646 12830 702
rect 12898 646 12954 702
rect 13022 646 13078 702
rect 12526 522 12582 578
rect 12650 522 12706 578
rect 12774 522 12830 578
rect 12898 522 12954 578
rect 13022 522 13078 578
rect -286 398 -230 454
rect -162 398 -106 454
rect -38 398 18 454
rect 86 398 142 454
rect 210 398 266 454
rect 12526 398 12582 454
rect 12650 398 12706 454
rect 12774 398 12830 454
rect 12898 398 12954 454
rect 13022 398 13078 454
rect -286 274 -230 330
rect -162 274 -106 330
rect -38 274 18 330
rect 86 274 142 330
rect 210 274 266 330
rect 415 246 471 302
rect 557 246 613 302
rect 699 246 755 302
rect 841 246 897 302
rect 983 246 1039 302
rect 1125 246 1181 302
rect 1267 246 1323 302
rect 1409 246 1465 302
rect 1551 246 1607 302
rect 1693 246 1749 302
rect 1835 246 1891 302
rect 1977 246 2033 302
rect 2119 246 2175 302
rect 2261 246 2317 302
rect 2403 246 2459 302
rect 2545 246 2601 302
rect 2687 246 2743 302
rect 2829 246 2885 302
rect 2971 246 3027 302
rect 3113 246 3169 302
rect 3255 246 3311 302
rect 3397 246 3453 302
rect 3539 246 3595 302
rect 3681 246 3737 302
rect 3823 246 3879 302
rect 3965 246 4021 302
rect 4107 246 4163 302
rect 4249 246 4305 302
rect 4391 246 4447 302
rect 4533 246 4589 302
rect 4675 246 4731 302
rect 4817 246 4873 302
rect 4959 246 5015 302
rect 5101 246 5157 302
rect 5243 246 5299 302
rect 5385 246 5441 302
rect 5527 246 5583 302
rect 5669 246 5725 302
rect 5811 246 5867 302
rect 5953 246 6009 302
rect 6095 246 6151 302
rect 6237 246 6293 302
rect 6379 246 6435 302
rect 6521 246 6577 302
rect 6663 246 6719 302
rect 6805 246 6861 302
rect 6947 246 7003 302
rect 7089 246 7145 302
rect 7231 246 7287 302
rect 7373 246 7429 302
rect 7515 246 7571 302
rect 7657 246 7713 302
rect 7799 246 7855 302
rect 7941 246 7997 302
rect 8083 246 8139 302
rect 8225 246 8281 302
rect 8367 246 8423 302
rect 8509 246 8565 302
rect 8651 246 8707 302
rect 8793 246 8849 302
rect 8935 246 8991 302
rect 9077 246 9133 302
rect 9219 246 9275 302
rect 9361 246 9417 302
rect 9503 246 9559 302
rect 9645 246 9701 302
rect 9787 246 9843 302
rect 9929 246 9985 302
rect 10071 246 10127 302
rect 10213 246 10269 302
rect 10355 246 10411 302
rect 10497 246 10553 302
rect 10639 246 10695 302
rect 10781 246 10837 302
rect 10923 246 10979 302
rect 11065 246 11121 302
rect 11207 246 11263 302
rect 11349 246 11405 302
rect 11491 246 11547 302
rect 11633 246 11689 302
rect 11775 246 11831 302
rect 11917 246 11973 302
rect 12059 246 12115 302
rect 12201 246 12257 302
rect 12343 246 12399 302
rect 12526 274 12582 330
rect 12650 274 12706 330
rect 12774 274 12830 330
rect 12898 274 12954 330
rect 13022 274 13078 330
rect -286 150 -230 206
rect -162 150 -106 206
rect -38 150 18 206
rect 86 150 142 206
rect 210 150 266 206
rect 415 104 471 160
rect 557 104 613 160
rect 699 104 755 160
rect 841 104 897 160
rect 983 104 1039 160
rect 1125 104 1181 160
rect 1267 104 1323 160
rect 1409 104 1465 160
rect 1551 104 1607 160
rect 1693 104 1749 160
rect 1835 104 1891 160
rect 1977 104 2033 160
rect 2119 104 2175 160
rect 2261 104 2317 160
rect 2403 104 2459 160
rect 2545 104 2601 160
rect 2687 104 2743 160
rect 2829 104 2885 160
rect 2971 104 3027 160
rect 3113 104 3169 160
rect 3255 104 3311 160
rect 3397 104 3453 160
rect 3539 104 3595 160
rect 3681 104 3737 160
rect 3823 104 3879 160
rect 3965 104 4021 160
rect 4107 104 4163 160
rect 4249 104 4305 160
rect 4391 104 4447 160
rect 4533 104 4589 160
rect 4675 104 4731 160
rect 4817 104 4873 160
rect 4959 104 5015 160
rect 5101 104 5157 160
rect 5243 104 5299 160
rect 5385 104 5441 160
rect 5527 104 5583 160
rect 5669 104 5725 160
rect 5811 104 5867 160
rect 5953 104 6009 160
rect 6095 104 6151 160
rect 6237 104 6293 160
rect 6379 104 6435 160
rect 6521 104 6577 160
rect 6663 104 6719 160
rect 6805 104 6861 160
rect 6947 104 7003 160
rect 7089 104 7145 160
rect 7231 104 7287 160
rect 7373 104 7429 160
rect 7515 104 7571 160
rect 7657 104 7713 160
rect 7799 104 7855 160
rect 7941 104 7997 160
rect 8083 104 8139 160
rect 8225 104 8281 160
rect 8367 104 8423 160
rect 8509 104 8565 160
rect 8651 104 8707 160
rect 8793 104 8849 160
rect 8935 104 8991 160
rect 9077 104 9133 160
rect 9219 104 9275 160
rect 9361 104 9417 160
rect 9503 104 9559 160
rect 9645 104 9701 160
rect 9787 104 9843 160
rect 9929 104 9985 160
rect 10071 104 10127 160
rect 10213 104 10269 160
rect 10355 104 10411 160
rect 10497 104 10553 160
rect 10639 104 10695 160
rect 10781 104 10837 160
rect 10923 104 10979 160
rect 11065 104 11121 160
rect 11207 104 11263 160
rect 11349 104 11405 160
rect 11491 104 11547 160
rect 11633 104 11689 160
rect 11775 104 11831 160
rect 11917 104 11973 160
rect 12059 104 12115 160
rect 12201 104 12257 160
rect 12343 104 12399 160
rect 12526 150 12582 206
rect 12650 150 12706 206
rect 12774 150 12830 206
rect 12898 150 12954 206
rect 13022 150 13078 206
<< metal5 >>
rect -400 12949 13200 13065
rect -400 12893 -254 12949
rect -198 12893 -130 12949
rect -74 12893 -6 12949
rect 50 12893 118 12949
rect 174 12893 242 12949
rect 298 12893 366 12949
rect 422 12893 490 12949
rect 546 12893 614 12949
rect 670 12893 738 12949
rect 794 12893 862 12949
rect 918 12893 986 12949
rect 1042 12893 1110 12949
rect 1166 12893 1234 12949
rect 1290 12893 1358 12949
rect 1414 12893 1482 12949
rect 1538 12893 1606 12949
rect 1662 12893 1730 12949
rect 1786 12893 1854 12949
rect 1910 12893 1978 12949
rect 2034 12893 2102 12949
rect 2158 12893 2226 12949
rect 2282 12893 2350 12949
rect 2406 12893 2474 12949
rect 2530 12893 2598 12949
rect 2654 12893 2722 12949
rect 2778 12893 2846 12949
rect 2902 12893 2970 12949
rect 3026 12893 3094 12949
rect 3150 12893 3218 12949
rect 3274 12893 3342 12949
rect 3398 12893 3466 12949
rect 3522 12893 3590 12949
rect 3646 12893 3714 12949
rect 3770 12893 3838 12949
rect 3894 12893 3962 12949
rect 4018 12893 4086 12949
rect 4142 12893 4210 12949
rect 4266 12893 4334 12949
rect 4390 12893 4458 12949
rect 4514 12893 4582 12949
rect 4638 12893 4706 12949
rect 4762 12893 4830 12949
rect 4886 12893 4954 12949
rect 5010 12893 5078 12949
rect 5134 12893 5202 12949
rect 5258 12893 5326 12949
rect 5382 12893 5450 12949
rect 5506 12893 5574 12949
rect 5630 12893 5698 12949
rect 5754 12893 5822 12949
rect 5878 12893 5946 12949
rect 6002 12893 6070 12949
rect 6126 12893 6194 12949
rect 6250 12893 6318 12949
rect 6374 12893 6442 12949
rect 6498 12893 6566 12949
rect 6622 12893 6690 12949
rect 6746 12893 6814 12949
rect 6870 12893 6938 12949
rect 6994 12893 7062 12949
rect 7118 12893 7186 12949
rect 7242 12893 7310 12949
rect 7366 12893 7434 12949
rect 7490 12893 7558 12949
rect 7614 12893 7682 12949
rect 7738 12893 7806 12949
rect 7862 12893 7930 12949
rect 7986 12893 8054 12949
rect 8110 12893 8178 12949
rect 8234 12893 8302 12949
rect 8358 12893 8426 12949
rect 8482 12893 8550 12949
rect 8606 12893 8674 12949
rect 8730 12893 8798 12949
rect 8854 12893 8922 12949
rect 8978 12893 9046 12949
rect 9102 12893 9170 12949
rect 9226 12893 9294 12949
rect 9350 12893 9418 12949
rect 9474 12893 9542 12949
rect 9598 12893 9666 12949
rect 9722 12893 9790 12949
rect 9846 12893 9914 12949
rect 9970 12893 10038 12949
rect 10094 12893 10162 12949
rect 10218 12893 10286 12949
rect 10342 12893 10410 12949
rect 10466 12893 10534 12949
rect 10590 12893 10658 12949
rect 10714 12893 10782 12949
rect 10838 12893 10906 12949
rect 10962 12893 11030 12949
rect 11086 12893 11154 12949
rect 11210 12893 11278 12949
rect 11334 12893 11402 12949
rect 11458 12893 11526 12949
rect 11582 12893 11650 12949
rect 11706 12893 11774 12949
rect 11830 12893 11898 12949
rect 11954 12893 12022 12949
rect 12078 12893 12146 12949
rect 12202 12893 12270 12949
rect 12326 12893 12394 12949
rect 12450 12893 12518 12949
rect 12574 12893 12642 12949
rect 12698 12893 12766 12949
rect 12822 12893 12890 12949
rect 12946 12893 13014 12949
rect 13070 12893 13200 12949
rect -400 12825 13200 12893
rect -400 12769 -254 12825
rect -198 12769 -130 12825
rect -74 12769 -6 12825
rect 50 12769 118 12825
rect 174 12769 242 12825
rect 298 12769 366 12825
rect 422 12769 490 12825
rect 546 12769 614 12825
rect 670 12769 738 12825
rect 794 12769 862 12825
rect 918 12769 986 12825
rect 1042 12769 1110 12825
rect 1166 12769 1234 12825
rect 1290 12769 1358 12825
rect 1414 12769 1482 12825
rect 1538 12769 1606 12825
rect 1662 12769 1730 12825
rect 1786 12769 1854 12825
rect 1910 12769 1978 12825
rect 2034 12769 2102 12825
rect 2158 12769 2226 12825
rect 2282 12769 2350 12825
rect 2406 12769 2474 12825
rect 2530 12769 2598 12825
rect 2654 12769 2722 12825
rect 2778 12769 2846 12825
rect 2902 12769 2970 12825
rect 3026 12769 3094 12825
rect 3150 12769 3218 12825
rect 3274 12769 3342 12825
rect 3398 12769 3466 12825
rect 3522 12769 3590 12825
rect 3646 12769 3714 12825
rect 3770 12769 3838 12825
rect 3894 12769 3962 12825
rect 4018 12769 4086 12825
rect 4142 12769 4210 12825
rect 4266 12769 4334 12825
rect 4390 12769 4458 12825
rect 4514 12769 4582 12825
rect 4638 12769 4706 12825
rect 4762 12769 4830 12825
rect 4886 12769 4954 12825
rect 5010 12769 5078 12825
rect 5134 12769 5202 12825
rect 5258 12769 5326 12825
rect 5382 12769 5450 12825
rect 5506 12769 5574 12825
rect 5630 12769 5698 12825
rect 5754 12769 5822 12825
rect 5878 12769 5946 12825
rect 6002 12769 6070 12825
rect 6126 12769 6194 12825
rect 6250 12769 6318 12825
rect 6374 12769 6442 12825
rect 6498 12769 6566 12825
rect 6622 12769 6690 12825
rect 6746 12769 6814 12825
rect 6870 12769 6938 12825
rect 6994 12769 7062 12825
rect 7118 12769 7186 12825
rect 7242 12769 7310 12825
rect 7366 12769 7434 12825
rect 7490 12769 7558 12825
rect 7614 12769 7682 12825
rect 7738 12769 7806 12825
rect 7862 12769 7930 12825
rect 7986 12769 8054 12825
rect 8110 12769 8178 12825
rect 8234 12769 8302 12825
rect 8358 12769 8426 12825
rect 8482 12769 8550 12825
rect 8606 12769 8674 12825
rect 8730 12769 8798 12825
rect 8854 12769 8922 12825
rect 8978 12769 9046 12825
rect 9102 12769 9170 12825
rect 9226 12769 9294 12825
rect 9350 12769 9418 12825
rect 9474 12769 9542 12825
rect 9598 12769 9666 12825
rect 9722 12769 9790 12825
rect 9846 12769 9914 12825
rect 9970 12769 10038 12825
rect 10094 12769 10162 12825
rect 10218 12769 10286 12825
rect 10342 12769 10410 12825
rect 10466 12769 10534 12825
rect 10590 12769 10658 12825
rect 10714 12769 10782 12825
rect 10838 12769 10906 12825
rect 10962 12769 11030 12825
rect 11086 12769 11154 12825
rect 11210 12769 11278 12825
rect 11334 12769 11402 12825
rect 11458 12769 11526 12825
rect 11582 12769 11650 12825
rect 11706 12769 11774 12825
rect 11830 12769 11898 12825
rect 11954 12769 12022 12825
rect 12078 12769 12146 12825
rect 12202 12769 12270 12825
rect 12326 12769 12394 12825
rect 12450 12769 12518 12825
rect 12574 12769 12642 12825
rect 12698 12769 12766 12825
rect 12822 12769 12890 12825
rect 12946 12769 13014 12825
rect 13070 12769 13200 12825
rect -400 12701 13200 12769
rect -400 12645 -254 12701
rect -198 12645 -130 12701
rect -74 12645 -6 12701
rect 50 12645 118 12701
rect 174 12645 242 12701
rect 298 12645 366 12701
rect 422 12645 490 12701
rect 546 12645 614 12701
rect 670 12645 738 12701
rect 794 12645 862 12701
rect 918 12645 986 12701
rect 1042 12645 1110 12701
rect 1166 12645 1234 12701
rect 1290 12645 1358 12701
rect 1414 12645 1482 12701
rect 1538 12645 1606 12701
rect 1662 12645 1730 12701
rect 1786 12645 1854 12701
rect 1910 12645 1978 12701
rect 2034 12645 2102 12701
rect 2158 12645 2226 12701
rect 2282 12645 2350 12701
rect 2406 12645 2474 12701
rect 2530 12645 2598 12701
rect 2654 12645 2722 12701
rect 2778 12645 2846 12701
rect 2902 12645 2970 12701
rect 3026 12645 3094 12701
rect 3150 12645 3218 12701
rect 3274 12645 3342 12701
rect 3398 12645 3466 12701
rect 3522 12645 3590 12701
rect 3646 12645 3714 12701
rect 3770 12645 3838 12701
rect 3894 12645 3962 12701
rect 4018 12645 4086 12701
rect 4142 12645 4210 12701
rect 4266 12645 4334 12701
rect 4390 12645 4458 12701
rect 4514 12645 4582 12701
rect 4638 12645 4706 12701
rect 4762 12645 4830 12701
rect 4886 12645 4954 12701
rect 5010 12645 5078 12701
rect 5134 12645 5202 12701
rect 5258 12645 5326 12701
rect 5382 12645 5450 12701
rect 5506 12645 5574 12701
rect 5630 12645 5698 12701
rect 5754 12645 5822 12701
rect 5878 12645 5946 12701
rect 6002 12645 6070 12701
rect 6126 12645 6194 12701
rect 6250 12645 6318 12701
rect 6374 12645 6442 12701
rect 6498 12645 6566 12701
rect 6622 12645 6690 12701
rect 6746 12645 6814 12701
rect 6870 12645 6938 12701
rect 6994 12645 7062 12701
rect 7118 12645 7186 12701
rect 7242 12645 7310 12701
rect 7366 12645 7434 12701
rect 7490 12645 7558 12701
rect 7614 12645 7682 12701
rect 7738 12645 7806 12701
rect 7862 12645 7930 12701
rect 7986 12645 8054 12701
rect 8110 12645 8178 12701
rect 8234 12645 8302 12701
rect 8358 12645 8426 12701
rect 8482 12645 8550 12701
rect 8606 12645 8674 12701
rect 8730 12645 8798 12701
rect 8854 12645 8922 12701
rect 8978 12645 9046 12701
rect 9102 12645 9170 12701
rect 9226 12645 9294 12701
rect 9350 12645 9418 12701
rect 9474 12645 9542 12701
rect 9598 12645 9666 12701
rect 9722 12645 9790 12701
rect 9846 12645 9914 12701
rect 9970 12645 10038 12701
rect 10094 12645 10162 12701
rect 10218 12645 10286 12701
rect 10342 12645 10410 12701
rect 10466 12645 10534 12701
rect 10590 12645 10658 12701
rect 10714 12645 10782 12701
rect 10838 12645 10906 12701
rect 10962 12645 11030 12701
rect 11086 12645 11154 12701
rect 11210 12645 11278 12701
rect 11334 12645 11402 12701
rect 11458 12645 11526 12701
rect 11582 12645 11650 12701
rect 11706 12645 11774 12701
rect 11830 12645 11898 12701
rect 11954 12645 12022 12701
rect 12078 12645 12146 12701
rect 12202 12645 12270 12701
rect 12326 12645 12394 12701
rect 12450 12645 12518 12701
rect 12574 12645 12642 12701
rect 12698 12645 12766 12701
rect 12822 12645 12890 12701
rect 12946 12645 13014 12701
rect 13070 12645 13200 12701
rect -400 12577 13200 12645
rect -400 12521 -254 12577
rect -198 12521 -130 12577
rect -74 12521 -6 12577
rect 50 12521 118 12577
rect 174 12521 242 12577
rect 298 12521 366 12577
rect 422 12521 490 12577
rect 546 12521 614 12577
rect 670 12521 738 12577
rect 794 12521 862 12577
rect 918 12521 986 12577
rect 1042 12521 1110 12577
rect 1166 12521 1234 12577
rect 1290 12521 1358 12577
rect 1414 12521 1482 12577
rect 1538 12521 1606 12577
rect 1662 12521 1730 12577
rect 1786 12521 1854 12577
rect 1910 12521 1978 12577
rect 2034 12521 2102 12577
rect 2158 12521 2226 12577
rect 2282 12521 2350 12577
rect 2406 12521 2474 12577
rect 2530 12521 2598 12577
rect 2654 12521 2722 12577
rect 2778 12521 2846 12577
rect 2902 12521 2970 12577
rect 3026 12521 3094 12577
rect 3150 12521 3218 12577
rect 3274 12521 3342 12577
rect 3398 12521 3466 12577
rect 3522 12521 3590 12577
rect 3646 12521 3714 12577
rect 3770 12521 3838 12577
rect 3894 12521 3962 12577
rect 4018 12521 4086 12577
rect 4142 12521 4210 12577
rect 4266 12521 4334 12577
rect 4390 12521 4458 12577
rect 4514 12521 4582 12577
rect 4638 12521 4706 12577
rect 4762 12521 4830 12577
rect 4886 12521 4954 12577
rect 5010 12521 5078 12577
rect 5134 12521 5202 12577
rect 5258 12521 5326 12577
rect 5382 12521 5450 12577
rect 5506 12521 5574 12577
rect 5630 12521 5698 12577
rect 5754 12521 5822 12577
rect 5878 12521 5946 12577
rect 6002 12521 6070 12577
rect 6126 12521 6194 12577
rect 6250 12521 6318 12577
rect 6374 12521 6442 12577
rect 6498 12521 6566 12577
rect 6622 12521 6690 12577
rect 6746 12521 6814 12577
rect 6870 12521 6938 12577
rect 6994 12521 7062 12577
rect 7118 12521 7186 12577
rect 7242 12521 7310 12577
rect 7366 12521 7434 12577
rect 7490 12521 7558 12577
rect 7614 12521 7682 12577
rect 7738 12521 7806 12577
rect 7862 12521 7930 12577
rect 7986 12521 8054 12577
rect 8110 12521 8178 12577
rect 8234 12521 8302 12577
rect 8358 12521 8426 12577
rect 8482 12521 8550 12577
rect 8606 12521 8674 12577
rect 8730 12521 8798 12577
rect 8854 12521 8922 12577
rect 8978 12521 9046 12577
rect 9102 12521 9170 12577
rect 9226 12521 9294 12577
rect 9350 12521 9418 12577
rect 9474 12521 9542 12577
rect 9598 12521 9666 12577
rect 9722 12521 9790 12577
rect 9846 12521 9914 12577
rect 9970 12521 10038 12577
rect 10094 12521 10162 12577
rect 10218 12521 10286 12577
rect 10342 12521 10410 12577
rect 10466 12521 10534 12577
rect 10590 12521 10658 12577
rect 10714 12521 10782 12577
rect 10838 12521 10906 12577
rect 10962 12521 11030 12577
rect 11086 12521 11154 12577
rect 11210 12521 11278 12577
rect 11334 12521 11402 12577
rect 11458 12521 11526 12577
rect 11582 12521 11650 12577
rect 11706 12521 11774 12577
rect 11830 12521 11898 12577
rect 11954 12521 12022 12577
rect 12078 12521 12146 12577
rect 12202 12521 12270 12577
rect 12326 12521 12394 12577
rect 12450 12521 12518 12577
rect 12574 12521 12642 12577
rect 12698 12521 12766 12577
rect 12822 12521 12890 12577
rect 12946 12521 13014 12577
rect 13070 12521 13200 12577
rect -400 12358 13200 12521
rect -400 12302 -286 12358
rect -230 12302 -162 12358
rect -106 12302 -38 12358
rect 18 12302 86 12358
rect 142 12302 210 12358
rect 266 12310 12526 12358
rect 266 12302 903 12310
rect -400 12254 903 12302
rect 959 12254 1045 12310
rect 1101 12254 1444 12310
rect 1500 12254 1586 12310
rect 1642 12254 1984 12310
rect 2040 12254 2126 12310
rect 2182 12254 2521 12310
rect 2577 12254 2663 12310
rect 2719 12254 3058 12310
rect 3114 12254 3200 12310
rect 3256 12254 3602 12310
rect 3658 12254 3744 12310
rect 3800 12254 4138 12310
rect 4194 12254 4280 12310
rect 4336 12254 4678 12310
rect 4734 12254 4820 12310
rect 4876 12254 5215 12310
rect 5271 12254 5357 12310
rect 5413 12254 5760 12310
rect 5816 12254 5902 12310
rect 5958 12254 6300 12310
rect 6356 12254 6442 12310
rect 6498 12254 6845 12310
rect 6901 12254 6987 12310
rect 7043 12254 7382 12310
rect 7438 12254 7524 12310
rect 7580 12254 7919 12310
rect 7975 12254 8061 12310
rect 8117 12254 8462 12310
rect 8518 12254 8604 12310
rect 8660 12254 9004 12310
rect 9060 12254 9146 12310
rect 9202 12254 9547 12310
rect 9603 12254 9689 12310
rect 9745 12254 10081 12310
rect 10137 12254 10223 12310
rect 10279 12254 10622 12310
rect 10678 12254 10764 12310
rect 10820 12254 11162 12310
rect 11218 12254 11304 12310
rect 11360 12254 11702 12310
rect 11758 12254 11844 12310
rect 11900 12302 12526 12310
rect 12582 12302 12650 12358
rect 12706 12302 12774 12358
rect 12830 12302 12898 12358
rect 12954 12302 13022 12358
rect 13078 12302 13200 12358
rect 11900 12254 13200 12302
rect -400 12234 13200 12254
rect -400 12178 -286 12234
rect -230 12178 -162 12234
rect -106 12178 -38 12234
rect 18 12178 86 12234
rect 142 12178 210 12234
rect 266 12178 12526 12234
rect 12582 12178 12650 12234
rect 12706 12178 12774 12234
rect 12830 12178 12898 12234
rect 12954 12178 13022 12234
rect 13078 12178 13200 12234
rect -400 12168 13200 12178
rect -400 12112 903 12168
rect 959 12112 1045 12168
rect 1101 12112 1444 12168
rect 1500 12112 1586 12168
rect 1642 12112 1984 12168
rect 2040 12112 2126 12168
rect 2182 12112 2521 12168
rect 2577 12112 2663 12168
rect 2719 12112 3058 12168
rect 3114 12112 3200 12168
rect 3256 12112 3602 12168
rect 3658 12112 3744 12168
rect 3800 12112 4138 12168
rect 4194 12112 4280 12168
rect 4336 12112 4678 12168
rect 4734 12112 4820 12168
rect 4876 12112 5215 12168
rect 5271 12112 5357 12168
rect 5413 12112 5760 12168
rect 5816 12112 5902 12168
rect 5958 12112 6300 12168
rect 6356 12112 6442 12168
rect 6498 12112 6845 12168
rect 6901 12112 6987 12168
rect 7043 12112 7382 12168
rect 7438 12112 7524 12168
rect 7580 12112 7919 12168
rect 7975 12112 8061 12168
rect 8117 12112 8462 12168
rect 8518 12112 8604 12168
rect 8660 12112 9004 12168
rect 9060 12112 9146 12168
rect 9202 12112 9547 12168
rect 9603 12112 9689 12168
rect 9745 12112 10081 12168
rect 10137 12112 10223 12168
rect 10279 12112 10622 12168
rect 10678 12112 10764 12168
rect 10820 12112 11162 12168
rect 11218 12112 11304 12168
rect 11360 12112 11702 12168
rect 11758 12112 11844 12168
rect 11900 12112 13200 12168
rect -400 12110 13200 12112
rect -400 12054 -286 12110
rect -230 12054 -162 12110
rect -106 12054 -38 12110
rect 18 12054 86 12110
rect 142 12054 210 12110
rect 266 12054 12526 12110
rect 12582 12054 12650 12110
rect 12706 12054 12774 12110
rect 12830 12054 12898 12110
rect 12954 12054 13022 12110
rect 13078 12054 13200 12110
rect -400 12026 13200 12054
rect -400 11986 903 12026
rect -400 11930 -286 11986
rect -230 11930 -162 11986
rect -106 11930 -38 11986
rect 18 11930 86 11986
rect 142 11930 210 11986
rect 266 11970 903 11986
rect 959 11970 1045 12026
rect 1101 11970 1444 12026
rect 1500 11970 1586 12026
rect 1642 11970 1984 12026
rect 2040 11970 2126 12026
rect 2182 11970 2521 12026
rect 2577 11970 2663 12026
rect 2719 11970 3058 12026
rect 3114 11970 3200 12026
rect 3256 11970 3602 12026
rect 3658 11970 3744 12026
rect 3800 11970 4138 12026
rect 4194 11970 4280 12026
rect 4336 11970 4678 12026
rect 4734 11970 4820 12026
rect 4876 11970 5215 12026
rect 5271 11970 5357 12026
rect 5413 11970 5760 12026
rect 5816 11970 5902 12026
rect 5958 11970 6300 12026
rect 6356 11970 6442 12026
rect 6498 11970 6845 12026
rect 6901 11970 6987 12026
rect 7043 11970 7382 12026
rect 7438 11970 7524 12026
rect 7580 11970 7919 12026
rect 7975 11970 8061 12026
rect 8117 11970 8462 12026
rect 8518 11970 8604 12026
rect 8660 11970 9004 12026
rect 9060 11970 9146 12026
rect 9202 11970 9547 12026
rect 9603 11970 9689 12026
rect 9745 11970 10081 12026
rect 10137 11970 10223 12026
rect 10279 11970 10622 12026
rect 10678 11970 10764 12026
rect 10820 11970 11162 12026
rect 11218 11970 11304 12026
rect 11360 11970 11702 12026
rect 11758 11970 11844 12026
rect 11900 11986 13200 12026
rect 11900 11970 12526 11986
rect 266 11930 12526 11970
rect 12582 11930 12650 11986
rect 12706 11930 12774 11986
rect 12830 11930 12898 11986
rect 12954 11930 13022 11986
rect 13078 11930 13200 11986
rect -400 11884 13200 11930
rect -400 11862 903 11884
rect -400 11806 -286 11862
rect -230 11806 -162 11862
rect -106 11806 -38 11862
rect 18 11806 86 11862
rect 142 11806 210 11862
rect 266 11828 903 11862
rect 959 11828 1045 11884
rect 1101 11828 1444 11884
rect 1500 11828 1586 11884
rect 1642 11828 1984 11884
rect 2040 11828 2126 11884
rect 2182 11828 2521 11884
rect 2577 11828 2663 11884
rect 2719 11828 3058 11884
rect 3114 11828 3200 11884
rect 3256 11828 3602 11884
rect 3658 11828 3744 11884
rect 3800 11828 4138 11884
rect 4194 11828 4280 11884
rect 4336 11828 4678 11884
rect 4734 11828 4820 11884
rect 4876 11828 5215 11884
rect 5271 11828 5357 11884
rect 5413 11828 5760 11884
rect 5816 11828 5902 11884
rect 5958 11828 6300 11884
rect 6356 11828 6442 11884
rect 6498 11828 6845 11884
rect 6901 11828 6987 11884
rect 7043 11828 7382 11884
rect 7438 11828 7524 11884
rect 7580 11828 7919 11884
rect 7975 11828 8061 11884
rect 8117 11828 8462 11884
rect 8518 11828 8604 11884
rect 8660 11828 9004 11884
rect 9060 11828 9146 11884
rect 9202 11828 9547 11884
rect 9603 11828 9689 11884
rect 9745 11828 10081 11884
rect 10137 11828 10223 11884
rect 10279 11828 10622 11884
rect 10678 11828 10764 11884
rect 10820 11828 11162 11884
rect 11218 11828 11304 11884
rect 11360 11828 11702 11884
rect 11758 11828 11844 11884
rect 11900 11862 13200 11884
rect 11900 11828 12526 11862
rect 266 11806 12526 11828
rect 12582 11806 12650 11862
rect 12706 11806 12774 11862
rect 12830 11806 12898 11862
rect 12954 11806 13022 11862
rect 13078 11806 13200 11862
rect -400 11742 13200 11806
rect -400 11738 903 11742
rect -400 11682 -286 11738
rect -230 11682 -162 11738
rect -106 11682 -38 11738
rect 18 11682 86 11738
rect 142 11682 210 11738
rect 266 11686 903 11738
rect 959 11686 1045 11742
rect 1101 11686 1444 11742
rect 1500 11686 1586 11742
rect 1642 11686 1984 11742
rect 2040 11686 2126 11742
rect 2182 11686 2521 11742
rect 2577 11686 2663 11742
rect 2719 11686 3058 11742
rect 3114 11686 3200 11742
rect 3256 11686 3602 11742
rect 3658 11686 3744 11742
rect 3800 11686 4138 11742
rect 4194 11686 4280 11742
rect 4336 11686 4678 11742
rect 4734 11686 4820 11742
rect 4876 11686 5215 11742
rect 5271 11686 5357 11742
rect 5413 11686 5760 11742
rect 5816 11686 5902 11742
rect 5958 11686 6300 11742
rect 6356 11686 6442 11742
rect 6498 11686 6845 11742
rect 6901 11686 6987 11742
rect 7043 11686 7382 11742
rect 7438 11686 7524 11742
rect 7580 11686 7919 11742
rect 7975 11686 8061 11742
rect 8117 11686 8462 11742
rect 8518 11686 8604 11742
rect 8660 11686 9004 11742
rect 9060 11686 9146 11742
rect 9202 11686 9547 11742
rect 9603 11686 9689 11742
rect 9745 11686 10081 11742
rect 10137 11686 10223 11742
rect 10279 11686 10622 11742
rect 10678 11686 10764 11742
rect 10820 11686 11162 11742
rect 11218 11686 11304 11742
rect 11360 11686 11702 11742
rect 11758 11686 11844 11742
rect 11900 11738 13200 11742
rect 11900 11686 12526 11738
rect 266 11682 12526 11686
rect 12582 11682 12650 11738
rect 12706 11682 12774 11738
rect 12830 11682 12898 11738
rect 12954 11682 13022 11738
rect 13078 11682 13200 11738
rect -400 11614 13200 11682
rect -400 11558 -286 11614
rect -230 11558 -162 11614
rect -106 11558 -38 11614
rect 18 11558 86 11614
rect 142 11558 210 11614
rect 266 11600 12526 11614
rect 266 11558 903 11600
rect -400 11544 903 11558
rect 959 11544 1045 11600
rect 1101 11544 1444 11600
rect 1500 11544 1586 11600
rect 1642 11544 1984 11600
rect 2040 11544 2126 11600
rect 2182 11544 2521 11600
rect 2577 11544 2663 11600
rect 2719 11544 3058 11600
rect 3114 11544 3200 11600
rect 3256 11544 3602 11600
rect 3658 11544 3744 11600
rect 3800 11544 4138 11600
rect 4194 11544 4280 11600
rect 4336 11544 4678 11600
rect 4734 11544 4820 11600
rect 4876 11544 5215 11600
rect 5271 11544 5357 11600
rect 5413 11544 5760 11600
rect 5816 11544 5902 11600
rect 5958 11544 6300 11600
rect 6356 11544 6442 11600
rect 6498 11544 6845 11600
rect 6901 11544 6987 11600
rect 7043 11544 7382 11600
rect 7438 11544 7524 11600
rect 7580 11544 7919 11600
rect 7975 11544 8061 11600
rect 8117 11544 8462 11600
rect 8518 11544 8604 11600
rect 8660 11544 9004 11600
rect 9060 11544 9146 11600
rect 9202 11544 9547 11600
rect 9603 11544 9689 11600
rect 9745 11544 10081 11600
rect 10137 11544 10223 11600
rect 10279 11544 10622 11600
rect 10678 11544 10764 11600
rect 10820 11544 11162 11600
rect 11218 11544 11304 11600
rect 11360 11544 11702 11600
rect 11758 11544 11844 11600
rect 11900 11558 12526 11600
rect 12582 11558 12650 11614
rect 12706 11558 12774 11614
rect 12830 11558 12898 11614
rect 12954 11558 13022 11614
rect 13078 11558 13200 11614
rect 11900 11544 13200 11558
rect -400 11490 13200 11544
rect -400 11434 -286 11490
rect -230 11434 -162 11490
rect -106 11434 -38 11490
rect 18 11434 86 11490
rect 142 11434 210 11490
rect 266 11458 12526 11490
rect 266 11434 903 11458
rect -400 11402 903 11434
rect 959 11402 1045 11458
rect 1101 11402 1444 11458
rect 1500 11402 1586 11458
rect 1642 11402 1984 11458
rect 2040 11402 2126 11458
rect 2182 11402 2521 11458
rect 2577 11402 2663 11458
rect 2719 11402 3058 11458
rect 3114 11402 3200 11458
rect 3256 11402 3602 11458
rect 3658 11402 3744 11458
rect 3800 11402 4138 11458
rect 4194 11402 4280 11458
rect 4336 11402 4678 11458
rect 4734 11402 4820 11458
rect 4876 11402 5215 11458
rect 5271 11402 5357 11458
rect 5413 11402 5760 11458
rect 5816 11402 5902 11458
rect 5958 11402 6300 11458
rect 6356 11402 6442 11458
rect 6498 11402 6845 11458
rect 6901 11402 6987 11458
rect 7043 11402 7382 11458
rect 7438 11402 7524 11458
rect 7580 11402 7919 11458
rect 7975 11402 8061 11458
rect 8117 11402 8462 11458
rect 8518 11402 8604 11458
rect 8660 11402 9004 11458
rect 9060 11402 9146 11458
rect 9202 11402 9547 11458
rect 9603 11402 9689 11458
rect 9745 11402 10081 11458
rect 10137 11402 10223 11458
rect 10279 11402 10622 11458
rect 10678 11402 10764 11458
rect 10820 11402 11162 11458
rect 11218 11402 11304 11458
rect 11360 11402 11702 11458
rect 11758 11402 11844 11458
rect 11900 11434 12526 11458
rect 12582 11434 12650 11490
rect 12706 11434 12774 11490
rect 12830 11434 12898 11490
rect 12954 11434 13022 11490
rect 13078 11434 13200 11490
rect 11900 11402 13200 11434
rect -400 11366 13200 11402
rect -400 11310 -286 11366
rect -230 11310 -162 11366
rect -106 11310 -38 11366
rect 18 11310 86 11366
rect 142 11310 210 11366
rect 266 11316 12526 11366
rect 266 11310 903 11316
rect -400 11260 903 11310
rect 959 11260 1045 11316
rect 1101 11260 1444 11316
rect 1500 11260 1586 11316
rect 1642 11260 1984 11316
rect 2040 11260 2126 11316
rect 2182 11260 2521 11316
rect 2577 11260 2663 11316
rect 2719 11260 3058 11316
rect 3114 11260 3200 11316
rect 3256 11260 3602 11316
rect 3658 11260 3744 11316
rect 3800 11260 4138 11316
rect 4194 11260 4280 11316
rect 4336 11260 4678 11316
rect 4734 11260 4820 11316
rect 4876 11260 5215 11316
rect 5271 11260 5357 11316
rect 5413 11260 5760 11316
rect 5816 11260 5902 11316
rect 5958 11260 6300 11316
rect 6356 11260 6442 11316
rect 6498 11260 6845 11316
rect 6901 11260 6987 11316
rect 7043 11260 7382 11316
rect 7438 11260 7524 11316
rect 7580 11260 7919 11316
rect 7975 11260 8061 11316
rect 8117 11260 8462 11316
rect 8518 11260 8604 11316
rect 8660 11260 9004 11316
rect 9060 11260 9146 11316
rect 9202 11260 9547 11316
rect 9603 11260 9689 11316
rect 9745 11260 10081 11316
rect 10137 11260 10223 11316
rect 10279 11260 10622 11316
rect 10678 11260 10764 11316
rect 10820 11260 11162 11316
rect 11218 11260 11304 11316
rect 11360 11260 11702 11316
rect 11758 11260 11844 11316
rect 11900 11310 12526 11316
rect 12582 11310 12650 11366
rect 12706 11310 12774 11366
rect 12830 11310 12898 11366
rect 12954 11310 13022 11366
rect 13078 11310 13200 11366
rect 11900 11260 13200 11310
rect -400 11242 13200 11260
rect -400 11186 -286 11242
rect -230 11186 -162 11242
rect -106 11186 -38 11242
rect 18 11186 86 11242
rect 142 11186 210 11242
rect 266 11186 12526 11242
rect 12582 11186 12650 11242
rect 12706 11186 12774 11242
rect 12830 11186 12898 11242
rect 12954 11186 13022 11242
rect 13078 11186 13200 11242
rect -400 11174 13200 11186
rect -400 11118 903 11174
rect 959 11118 1045 11174
rect 1101 11118 1444 11174
rect 1500 11118 1586 11174
rect 1642 11118 1984 11174
rect 2040 11118 2126 11174
rect 2182 11118 2521 11174
rect 2577 11118 2663 11174
rect 2719 11118 3058 11174
rect 3114 11118 3200 11174
rect 3256 11118 3602 11174
rect 3658 11118 3744 11174
rect 3800 11118 4138 11174
rect 4194 11118 4280 11174
rect 4336 11118 4678 11174
rect 4734 11118 4820 11174
rect 4876 11118 5215 11174
rect 5271 11118 5357 11174
rect 5413 11118 5760 11174
rect 5816 11118 5902 11174
rect 5958 11118 6300 11174
rect 6356 11118 6442 11174
rect 6498 11118 6845 11174
rect 6901 11118 6987 11174
rect 7043 11118 7382 11174
rect 7438 11118 7524 11174
rect 7580 11118 7919 11174
rect 7975 11118 8061 11174
rect 8117 11118 8462 11174
rect 8518 11118 8604 11174
rect 8660 11118 9004 11174
rect 9060 11118 9146 11174
rect 9202 11118 9547 11174
rect 9603 11118 9689 11174
rect 9745 11118 10081 11174
rect 10137 11118 10223 11174
rect 10279 11118 10622 11174
rect 10678 11118 10764 11174
rect 10820 11118 11162 11174
rect 11218 11118 11304 11174
rect 11360 11118 11702 11174
rect 11758 11118 11844 11174
rect 11900 11118 13200 11174
rect -400 11062 -286 11118
rect -230 11062 -162 11118
rect -106 11062 -38 11118
rect 18 11062 86 11118
rect 142 11062 210 11118
rect 266 11062 12526 11118
rect 12582 11062 12650 11118
rect 12706 11062 12774 11118
rect 12830 11062 12898 11118
rect 12954 11062 13022 11118
rect 13078 11062 13200 11118
rect -400 11032 13200 11062
rect -400 10994 903 11032
rect -400 10938 -286 10994
rect -230 10938 -162 10994
rect -106 10938 -38 10994
rect 18 10938 86 10994
rect 142 10938 210 10994
rect 266 10976 903 10994
rect 959 10976 1045 11032
rect 1101 10976 1444 11032
rect 1500 10976 1586 11032
rect 1642 10976 1984 11032
rect 2040 10976 2126 11032
rect 2182 10976 2521 11032
rect 2577 10976 2663 11032
rect 2719 10976 3058 11032
rect 3114 10976 3200 11032
rect 3256 10976 3602 11032
rect 3658 10976 3744 11032
rect 3800 10976 4138 11032
rect 4194 10976 4280 11032
rect 4336 10976 4678 11032
rect 4734 10976 4820 11032
rect 4876 10976 5215 11032
rect 5271 10976 5357 11032
rect 5413 10976 5760 11032
rect 5816 10976 5902 11032
rect 5958 10976 6300 11032
rect 6356 10976 6442 11032
rect 6498 10976 6845 11032
rect 6901 10976 6987 11032
rect 7043 10976 7382 11032
rect 7438 10976 7524 11032
rect 7580 10976 7919 11032
rect 7975 10976 8061 11032
rect 8117 10976 8462 11032
rect 8518 10976 8604 11032
rect 8660 10976 9004 11032
rect 9060 10976 9146 11032
rect 9202 10976 9547 11032
rect 9603 10976 9689 11032
rect 9745 10976 10081 11032
rect 10137 10976 10223 11032
rect 10279 10976 10622 11032
rect 10678 10976 10764 11032
rect 10820 10976 11162 11032
rect 11218 10976 11304 11032
rect 11360 10976 11702 11032
rect 11758 10976 11844 11032
rect 11900 10994 13200 11032
rect 11900 10976 12526 10994
rect 266 10938 12526 10976
rect 12582 10938 12650 10994
rect 12706 10938 12774 10994
rect 12830 10938 12898 10994
rect 12954 10938 13022 10994
rect 13078 10938 13200 10994
rect -400 10890 13200 10938
rect -400 10870 903 10890
rect -400 10814 -286 10870
rect -230 10814 -162 10870
rect -106 10814 -38 10870
rect 18 10814 86 10870
rect 142 10814 210 10870
rect 266 10834 903 10870
rect 959 10834 1045 10890
rect 1101 10834 1444 10890
rect 1500 10834 1586 10890
rect 1642 10834 1984 10890
rect 2040 10834 2126 10890
rect 2182 10834 2521 10890
rect 2577 10834 2663 10890
rect 2719 10834 3058 10890
rect 3114 10834 3200 10890
rect 3256 10834 3602 10890
rect 3658 10834 3744 10890
rect 3800 10834 4138 10890
rect 4194 10834 4280 10890
rect 4336 10834 4678 10890
rect 4734 10834 4820 10890
rect 4876 10834 5215 10890
rect 5271 10834 5357 10890
rect 5413 10834 5760 10890
rect 5816 10834 5902 10890
rect 5958 10834 6300 10890
rect 6356 10834 6442 10890
rect 6498 10834 6845 10890
rect 6901 10834 6987 10890
rect 7043 10834 7382 10890
rect 7438 10834 7524 10890
rect 7580 10834 7919 10890
rect 7975 10834 8061 10890
rect 8117 10834 8462 10890
rect 8518 10834 8604 10890
rect 8660 10834 9004 10890
rect 9060 10834 9146 10890
rect 9202 10834 9547 10890
rect 9603 10834 9689 10890
rect 9745 10834 10081 10890
rect 10137 10834 10223 10890
rect 10279 10834 10622 10890
rect 10678 10834 10764 10890
rect 10820 10834 11162 10890
rect 11218 10834 11304 10890
rect 11360 10834 11702 10890
rect 11758 10834 11844 10890
rect 11900 10870 13200 10890
rect 11900 10834 12526 10870
rect 266 10814 12526 10834
rect 12582 10814 12650 10870
rect 12706 10814 12774 10870
rect 12830 10814 12898 10870
rect 12954 10814 13022 10870
rect 13078 10814 13200 10870
rect -400 10748 13200 10814
rect -400 10746 903 10748
rect -400 10690 -286 10746
rect -230 10690 -162 10746
rect -106 10690 -38 10746
rect 18 10690 86 10746
rect 142 10690 210 10746
rect 266 10692 903 10746
rect 959 10692 1045 10748
rect 1101 10692 1444 10748
rect 1500 10692 1586 10748
rect 1642 10692 1984 10748
rect 2040 10692 2126 10748
rect 2182 10692 2521 10748
rect 2577 10692 2663 10748
rect 2719 10692 3058 10748
rect 3114 10692 3200 10748
rect 3256 10692 3602 10748
rect 3658 10692 3744 10748
rect 3800 10692 4138 10748
rect 4194 10692 4280 10748
rect 4336 10692 4678 10748
rect 4734 10692 4820 10748
rect 4876 10692 5215 10748
rect 5271 10692 5357 10748
rect 5413 10692 5760 10748
rect 5816 10692 5902 10748
rect 5958 10692 6300 10748
rect 6356 10692 6442 10748
rect 6498 10692 6845 10748
rect 6901 10692 6987 10748
rect 7043 10692 7382 10748
rect 7438 10692 7524 10748
rect 7580 10692 7919 10748
rect 7975 10692 8061 10748
rect 8117 10692 8462 10748
rect 8518 10692 8604 10748
rect 8660 10692 9004 10748
rect 9060 10692 9146 10748
rect 9202 10692 9547 10748
rect 9603 10692 9689 10748
rect 9745 10692 10081 10748
rect 10137 10692 10223 10748
rect 10279 10692 10622 10748
rect 10678 10692 10764 10748
rect 10820 10692 11162 10748
rect 11218 10692 11304 10748
rect 11360 10692 11702 10748
rect 11758 10692 11844 10748
rect 11900 10746 13200 10748
rect 11900 10692 12526 10746
rect 266 10690 12526 10692
rect 12582 10690 12650 10746
rect 12706 10690 12774 10746
rect 12830 10690 12898 10746
rect 12954 10690 13022 10746
rect 13078 10690 13200 10746
rect -400 10622 13200 10690
rect -400 10566 -286 10622
rect -230 10566 -162 10622
rect -106 10566 -38 10622
rect 18 10566 86 10622
rect 142 10566 210 10622
rect 266 10606 12526 10622
rect 266 10566 903 10606
rect -400 10550 903 10566
rect 959 10550 1045 10606
rect 1101 10550 1444 10606
rect 1500 10550 1586 10606
rect 1642 10550 1984 10606
rect 2040 10550 2126 10606
rect 2182 10550 2521 10606
rect 2577 10550 2663 10606
rect 2719 10550 3058 10606
rect 3114 10550 3200 10606
rect 3256 10550 3602 10606
rect 3658 10550 3744 10606
rect 3800 10550 4138 10606
rect 4194 10550 4280 10606
rect 4336 10550 4678 10606
rect 4734 10550 4820 10606
rect 4876 10550 5215 10606
rect 5271 10550 5357 10606
rect 5413 10550 5760 10606
rect 5816 10550 5902 10606
rect 5958 10550 6300 10606
rect 6356 10550 6442 10606
rect 6498 10550 6845 10606
rect 6901 10550 6987 10606
rect 7043 10550 7382 10606
rect 7438 10550 7524 10606
rect 7580 10550 7919 10606
rect 7975 10550 8061 10606
rect 8117 10550 8462 10606
rect 8518 10550 8604 10606
rect 8660 10550 9004 10606
rect 9060 10550 9146 10606
rect 9202 10550 9547 10606
rect 9603 10550 9689 10606
rect 9745 10550 10081 10606
rect 10137 10550 10223 10606
rect 10279 10550 10622 10606
rect 10678 10550 10764 10606
rect 10820 10550 11162 10606
rect 11218 10550 11304 10606
rect 11360 10550 11702 10606
rect 11758 10550 11844 10606
rect 11900 10566 12526 10606
rect 12582 10566 12650 10622
rect 12706 10566 12774 10622
rect 12830 10566 12898 10622
rect 12954 10566 13022 10622
rect 13078 10566 13200 10622
rect 11900 10550 13200 10566
rect -400 10498 13200 10550
rect -400 10442 -286 10498
rect -230 10442 -162 10498
rect -106 10442 -38 10498
rect 18 10442 86 10498
rect 142 10442 210 10498
rect 266 10464 12526 10498
rect 266 10442 903 10464
rect -400 10408 903 10442
rect 959 10408 1045 10464
rect 1101 10408 1444 10464
rect 1500 10408 1586 10464
rect 1642 10408 1984 10464
rect 2040 10408 2126 10464
rect 2182 10408 2521 10464
rect 2577 10408 2663 10464
rect 2719 10408 3058 10464
rect 3114 10408 3200 10464
rect 3256 10408 3602 10464
rect 3658 10408 3744 10464
rect 3800 10408 4138 10464
rect 4194 10408 4280 10464
rect 4336 10408 4678 10464
rect 4734 10408 4820 10464
rect 4876 10408 5215 10464
rect 5271 10408 5357 10464
rect 5413 10408 5760 10464
rect 5816 10408 5902 10464
rect 5958 10408 6300 10464
rect 6356 10408 6442 10464
rect 6498 10408 6845 10464
rect 6901 10408 6987 10464
rect 7043 10408 7382 10464
rect 7438 10408 7524 10464
rect 7580 10408 7919 10464
rect 7975 10408 8061 10464
rect 8117 10408 8462 10464
rect 8518 10408 8604 10464
rect 8660 10408 9004 10464
rect 9060 10408 9146 10464
rect 9202 10408 9547 10464
rect 9603 10408 9689 10464
rect 9745 10408 10081 10464
rect 10137 10408 10223 10464
rect 10279 10408 10622 10464
rect 10678 10408 10764 10464
rect 10820 10408 11162 10464
rect 11218 10408 11304 10464
rect 11360 10408 11702 10464
rect 11758 10408 11844 10464
rect 11900 10442 12526 10464
rect 12582 10442 12650 10498
rect 12706 10442 12774 10498
rect 12830 10442 12898 10498
rect 12954 10442 13022 10498
rect 13078 10442 13200 10498
rect 11900 10408 13200 10442
rect -400 10374 13200 10408
rect -400 10318 -286 10374
rect -230 10318 -162 10374
rect -106 10318 -38 10374
rect 18 10318 86 10374
rect 142 10318 210 10374
rect 266 10322 12526 10374
rect 266 10318 903 10322
rect -400 10266 903 10318
rect 959 10266 1045 10322
rect 1101 10266 1444 10322
rect 1500 10266 1586 10322
rect 1642 10266 1984 10322
rect 2040 10266 2126 10322
rect 2182 10266 2521 10322
rect 2577 10266 2663 10322
rect 2719 10266 3058 10322
rect 3114 10266 3200 10322
rect 3256 10266 3602 10322
rect 3658 10266 3744 10322
rect 3800 10266 4138 10322
rect 4194 10266 4280 10322
rect 4336 10266 4678 10322
rect 4734 10266 4820 10322
rect 4876 10266 5215 10322
rect 5271 10266 5357 10322
rect 5413 10266 5760 10322
rect 5816 10266 5902 10322
rect 5958 10266 6300 10322
rect 6356 10266 6442 10322
rect 6498 10266 6845 10322
rect 6901 10266 6987 10322
rect 7043 10266 7382 10322
rect 7438 10266 7524 10322
rect 7580 10266 7919 10322
rect 7975 10266 8061 10322
rect 8117 10266 8462 10322
rect 8518 10266 8604 10322
rect 8660 10266 9004 10322
rect 9060 10266 9146 10322
rect 9202 10266 9547 10322
rect 9603 10266 9689 10322
rect 9745 10266 10081 10322
rect 10137 10266 10223 10322
rect 10279 10266 10622 10322
rect 10678 10266 10764 10322
rect 10820 10266 11162 10322
rect 11218 10266 11304 10322
rect 11360 10266 11702 10322
rect 11758 10266 11844 10322
rect 11900 10318 12526 10322
rect 12582 10318 12650 10374
rect 12706 10318 12774 10374
rect 12830 10318 12898 10374
rect 12954 10318 13022 10374
rect 13078 10318 13200 10374
rect 11900 10266 13200 10318
rect -400 10250 13200 10266
rect -400 10194 -286 10250
rect -230 10194 -162 10250
rect -106 10194 -38 10250
rect 18 10194 86 10250
rect 142 10194 210 10250
rect 266 10194 12526 10250
rect 12582 10194 12650 10250
rect 12706 10194 12774 10250
rect 12830 10194 12898 10250
rect 12954 10194 13022 10250
rect 13078 10194 13200 10250
rect -400 10180 13200 10194
rect -400 10126 903 10180
rect -400 10070 -286 10126
rect -230 10070 -162 10126
rect -106 10070 -38 10126
rect 18 10070 86 10126
rect 142 10070 210 10126
rect 266 10124 903 10126
rect 959 10124 1045 10180
rect 1101 10124 1444 10180
rect 1500 10124 1586 10180
rect 1642 10124 1984 10180
rect 2040 10124 2126 10180
rect 2182 10124 2521 10180
rect 2577 10124 2663 10180
rect 2719 10124 3058 10180
rect 3114 10124 3200 10180
rect 3256 10124 3602 10180
rect 3658 10124 3744 10180
rect 3800 10124 4138 10180
rect 4194 10124 4280 10180
rect 4336 10124 4678 10180
rect 4734 10124 4820 10180
rect 4876 10124 5215 10180
rect 5271 10124 5357 10180
rect 5413 10124 5760 10180
rect 5816 10124 5902 10180
rect 5958 10124 6300 10180
rect 6356 10124 6442 10180
rect 6498 10124 6845 10180
rect 6901 10124 6987 10180
rect 7043 10124 7382 10180
rect 7438 10124 7524 10180
rect 7580 10124 7919 10180
rect 7975 10124 8061 10180
rect 8117 10124 8462 10180
rect 8518 10124 8604 10180
rect 8660 10124 9004 10180
rect 9060 10124 9146 10180
rect 9202 10124 9547 10180
rect 9603 10124 9689 10180
rect 9745 10124 10081 10180
rect 10137 10124 10223 10180
rect 10279 10124 10622 10180
rect 10678 10124 10764 10180
rect 10820 10124 11162 10180
rect 11218 10124 11304 10180
rect 11360 10124 11702 10180
rect 11758 10124 11844 10180
rect 11900 10126 13200 10180
rect 11900 10124 12526 10126
rect 266 10070 12526 10124
rect 12582 10070 12650 10126
rect 12706 10070 12774 10126
rect 12830 10070 12898 10126
rect 12954 10070 13022 10126
rect 13078 10070 13200 10126
rect -400 10038 13200 10070
rect -400 10002 903 10038
rect -400 9946 -286 10002
rect -230 9946 -162 10002
rect -106 9946 -38 10002
rect 18 9946 86 10002
rect 142 9946 210 10002
rect 266 9982 903 10002
rect 959 9982 1045 10038
rect 1101 9982 1444 10038
rect 1500 9982 1586 10038
rect 1642 9982 1984 10038
rect 2040 9982 2126 10038
rect 2182 9982 2521 10038
rect 2577 9982 2663 10038
rect 2719 9982 3058 10038
rect 3114 9982 3200 10038
rect 3256 9982 3602 10038
rect 3658 9982 3744 10038
rect 3800 9982 4138 10038
rect 4194 9982 4280 10038
rect 4336 9982 4678 10038
rect 4734 9982 4820 10038
rect 4876 9982 5215 10038
rect 5271 9982 5357 10038
rect 5413 9982 5760 10038
rect 5816 9982 5902 10038
rect 5958 9982 6300 10038
rect 6356 9982 6442 10038
rect 6498 9982 6845 10038
rect 6901 9982 6987 10038
rect 7043 9982 7382 10038
rect 7438 9982 7524 10038
rect 7580 9982 7919 10038
rect 7975 9982 8061 10038
rect 8117 9982 8462 10038
rect 8518 9982 8604 10038
rect 8660 9982 9004 10038
rect 9060 9982 9146 10038
rect 9202 9982 9547 10038
rect 9603 9982 9689 10038
rect 9745 9982 10081 10038
rect 10137 9982 10223 10038
rect 10279 9982 10622 10038
rect 10678 9982 10764 10038
rect 10820 9982 11162 10038
rect 11218 9982 11304 10038
rect 11360 9982 11702 10038
rect 11758 9982 11844 10038
rect 11900 10002 13200 10038
rect 11900 9982 12526 10002
rect 266 9946 12526 9982
rect 12582 9946 12650 10002
rect 12706 9946 12774 10002
rect 12830 9946 12898 10002
rect 12954 9946 13022 10002
rect 13078 9946 13200 10002
rect -400 9896 13200 9946
rect -400 9878 903 9896
rect -400 9822 -286 9878
rect -230 9822 -162 9878
rect -106 9822 -38 9878
rect 18 9822 86 9878
rect 142 9822 210 9878
rect 266 9840 903 9878
rect 959 9840 1045 9896
rect 1101 9840 1444 9896
rect 1500 9840 1586 9896
rect 1642 9840 1984 9896
rect 2040 9840 2126 9896
rect 2182 9840 2521 9896
rect 2577 9840 2663 9896
rect 2719 9840 3058 9896
rect 3114 9840 3200 9896
rect 3256 9840 3602 9896
rect 3658 9840 3744 9896
rect 3800 9840 4138 9896
rect 4194 9840 4280 9896
rect 4336 9840 4678 9896
rect 4734 9840 4820 9896
rect 4876 9840 5215 9896
rect 5271 9840 5357 9896
rect 5413 9840 5760 9896
rect 5816 9840 5902 9896
rect 5958 9840 6300 9896
rect 6356 9840 6442 9896
rect 6498 9840 6845 9896
rect 6901 9840 6987 9896
rect 7043 9840 7382 9896
rect 7438 9840 7524 9896
rect 7580 9840 7919 9896
rect 7975 9840 8061 9896
rect 8117 9840 8462 9896
rect 8518 9840 8604 9896
rect 8660 9840 9004 9896
rect 9060 9840 9146 9896
rect 9202 9840 9547 9896
rect 9603 9840 9689 9896
rect 9745 9840 10081 9896
rect 10137 9840 10223 9896
rect 10279 9840 10622 9896
rect 10678 9840 10764 9896
rect 10820 9840 11162 9896
rect 11218 9840 11304 9896
rect 11360 9840 11702 9896
rect 11758 9840 11844 9896
rect 11900 9878 13200 9896
rect 11900 9840 12526 9878
rect 266 9822 12526 9840
rect 12582 9822 12650 9878
rect 12706 9822 12774 9878
rect 12830 9822 12898 9878
rect 12954 9822 13022 9878
rect 13078 9822 13200 9878
rect -400 9754 13200 9822
rect -400 9698 -286 9754
rect -230 9698 -162 9754
rect -106 9698 -38 9754
rect 18 9698 86 9754
rect 142 9698 210 9754
rect 266 9698 903 9754
rect 959 9698 1045 9754
rect 1101 9698 1444 9754
rect 1500 9698 1586 9754
rect 1642 9698 1984 9754
rect 2040 9698 2126 9754
rect 2182 9698 2521 9754
rect 2577 9698 2663 9754
rect 2719 9698 3058 9754
rect 3114 9698 3200 9754
rect 3256 9698 3602 9754
rect 3658 9698 3744 9754
rect 3800 9698 4138 9754
rect 4194 9698 4280 9754
rect 4336 9698 4678 9754
rect 4734 9698 4820 9754
rect 4876 9698 5215 9754
rect 5271 9698 5357 9754
rect 5413 9698 5760 9754
rect 5816 9698 5902 9754
rect 5958 9698 6300 9754
rect 6356 9698 6442 9754
rect 6498 9698 6845 9754
rect 6901 9698 6987 9754
rect 7043 9698 7382 9754
rect 7438 9698 7524 9754
rect 7580 9698 7919 9754
rect 7975 9698 8061 9754
rect 8117 9698 8462 9754
rect 8518 9698 8604 9754
rect 8660 9698 9004 9754
rect 9060 9698 9146 9754
rect 9202 9698 9547 9754
rect 9603 9698 9689 9754
rect 9745 9698 10081 9754
rect 10137 9698 10223 9754
rect 10279 9698 10622 9754
rect 10678 9698 10764 9754
rect 10820 9698 11162 9754
rect 11218 9698 11304 9754
rect 11360 9698 11702 9754
rect 11758 9698 11844 9754
rect 11900 9698 12526 9754
rect 12582 9698 12650 9754
rect 12706 9698 12774 9754
rect 12830 9698 12898 9754
rect 12954 9698 13022 9754
rect 13078 9698 13200 9754
rect -400 9630 13200 9698
rect -400 9574 -286 9630
rect -230 9574 -162 9630
rect -106 9574 -38 9630
rect 18 9574 86 9630
rect 142 9574 210 9630
rect 266 9612 12526 9630
rect 266 9574 903 9612
rect -400 9556 903 9574
rect 959 9556 1045 9612
rect 1101 9556 1444 9612
rect 1500 9556 1586 9612
rect 1642 9556 1984 9612
rect 2040 9556 2126 9612
rect 2182 9556 2521 9612
rect 2577 9556 2663 9612
rect 2719 9556 3058 9612
rect 3114 9556 3200 9612
rect 3256 9556 3602 9612
rect 3658 9556 3744 9612
rect 3800 9556 4138 9612
rect 4194 9556 4280 9612
rect 4336 9556 4678 9612
rect 4734 9556 4820 9612
rect 4876 9556 5215 9612
rect 5271 9556 5357 9612
rect 5413 9556 5760 9612
rect 5816 9556 5902 9612
rect 5958 9556 6300 9612
rect 6356 9556 6442 9612
rect 6498 9556 6845 9612
rect 6901 9556 6987 9612
rect 7043 9556 7382 9612
rect 7438 9556 7524 9612
rect 7580 9556 7919 9612
rect 7975 9556 8061 9612
rect 8117 9556 8462 9612
rect 8518 9556 8604 9612
rect 8660 9556 9004 9612
rect 9060 9556 9146 9612
rect 9202 9556 9547 9612
rect 9603 9556 9689 9612
rect 9745 9556 10081 9612
rect 10137 9556 10223 9612
rect 10279 9556 10622 9612
rect 10678 9556 10764 9612
rect 10820 9556 11162 9612
rect 11218 9556 11304 9612
rect 11360 9556 11702 9612
rect 11758 9556 11844 9612
rect 11900 9574 12526 9612
rect 12582 9574 12650 9630
rect 12706 9574 12774 9630
rect 12830 9574 12898 9630
rect 12954 9574 13022 9630
rect 13078 9574 13200 9630
rect 11900 9556 13200 9574
rect -400 9506 13200 9556
rect -400 9450 -286 9506
rect -230 9450 -162 9506
rect -106 9450 -38 9506
rect 18 9450 86 9506
rect 142 9450 210 9506
rect 266 9470 12526 9506
rect 266 9450 903 9470
rect -400 9414 903 9450
rect 959 9414 1045 9470
rect 1101 9414 1444 9470
rect 1500 9414 1586 9470
rect 1642 9414 1984 9470
rect 2040 9414 2126 9470
rect 2182 9414 2521 9470
rect 2577 9414 2663 9470
rect 2719 9414 3058 9470
rect 3114 9414 3200 9470
rect 3256 9414 3602 9470
rect 3658 9414 3744 9470
rect 3800 9414 4138 9470
rect 4194 9414 4280 9470
rect 4336 9414 4678 9470
rect 4734 9414 4820 9470
rect 4876 9414 5215 9470
rect 5271 9414 5357 9470
rect 5413 9414 5760 9470
rect 5816 9414 5902 9470
rect 5958 9414 6300 9470
rect 6356 9414 6442 9470
rect 6498 9414 6845 9470
rect 6901 9414 6987 9470
rect 7043 9414 7382 9470
rect 7438 9414 7524 9470
rect 7580 9414 7919 9470
rect 7975 9414 8061 9470
rect 8117 9414 8462 9470
rect 8518 9414 8604 9470
rect 8660 9414 9004 9470
rect 9060 9414 9146 9470
rect 9202 9414 9547 9470
rect 9603 9414 9689 9470
rect 9745 9414 10081 9470
rect 10137 9414 10223 9470
rect 10279 9414 10622 9470
rect 10678 9414 10764 9470
rect 10820 9414 11162 9470
rect 11218 9414 11304 9470
rect 11360 9414 11702 9470
rect 11758 9414 11844 9470
rect 11900 9450 12526 9470
rect 12582 9450 12650 9506
rect 12706 9450 12774 9506
rect 12830 9450 12898 9506
rect 12954 9450 13022 9506
rect 13078 9450 13200 9506
rect 11900 9414 13200 9450
rect -400 9382 13200 9414
rect -400 9326 -286 9382
rect -230 9326 -162 9382
rect -106 9326 -38 9382
rect 18 9326 86 9382
rect 142 9326 210 9382
rect 266 9328 12526 9382
rect 266 9326 903 9328
rect -400 9272 903 9326
rect 959 9272 1045 9328
rect 1101 9272 1444 9328
rect 1500 9272 1586 9328
rect 1642 9272 1984 9328
rect 2040 9272 2126 9328
rect 2182 9272 2521 9328
rect 2577 9272 2663 9328
rect 2719 9272 3058 9328
rect 3114 9272 3200 9328
rect 3256 9272 3602 9328
rect 3658 9272 3744 9328
rect 3800 9272 4138 9328
rect 4194 9272 4280 9328
rect 4336 9272 4678 9328
rect 4734 9272 4820 9328
rect 4876 9272 5215 9328
rect 5271 9272 5357 9328
rect 5413 9272 5760 9328
rect 5816 9272 5902 9328
rect 5958 9272 6300 9328
rect 6356 9272 6442 9328
rect 6498 9272 6845 9328
rect 6901 9272 6987 9328
rect 7043 9272 7382 9328
rect 7438 9272 7524 9328
rect 7580 9272 7919 9328
rect 7975 9272 8061 9328
rect 8117 9272 8462 9328
rect 8518 9272 8604 9328
rect 8660 9272 9004 9328
rect 9060 9272 9146 9328
rect 9202 9272 9547 9328
rect 9603 9272 9689 9328
rect 9745 9272 10081 9328
rect 10137 9272 10223 9328
rect 10279 9272 10622 9328
rect 10678 9272 10764 9328
rect 10820 9272 11162 9328
rect 11218 9272 11304 9328
rect 11360 9272 11702 9328
rect 11758 9272 11844 9328
rect 11900 9326 12526 9328
rect 12582 9326 12650 9382
rect 12706 9326 12774 9382
rect 12830 9326 12898 9382
rect 12954 9326 13022 9382
rect 13078 9326 13200 9382
rect 11900 9272 13200 9326
rect -400 9258 13200 9272
rect -400 9202 -286 9258
rect -230 9202 -162 9258
rect -106 9202 -38 9258
rect 18 9202 86 9258
rect 142 9202 210 9258
rect 266 9202 12526 9258
rect 12582 9202 12650 9258
rect 12706 9202 12774 9258
rect 12830 9202 12898 9258
rect 12954 9202 13022 9258
rect 13078 9202 13200 9258
rect -400 9186 13200 9202
rect -400 9134 903 9186
rect -400 9078 -286 9134
rect -230 9078 -162 9134
rect -106 9078 -38 9134
rect 18 9078 86 9134
rect 142 9078 210 9134
rect 266 9130 903 9134
rect 959 9130 1045 9186
rect 1101 9130 1444 9186
rect 1500 9130 1586 9186
rect 1642 9130 1984 9186
rect 2040 9130 2126 9186
rect 2182 9130 2521 9186
rect 2577 9130 2663 9186
rect 2719 9130 3058 9186
rect 3114 9130 3200 9186
rect 3256 9130 3602 9186
rect 3658 9130 3744 9186
rect 3800 9130 4138 9186
rect 4194 9130 4280 9186
rect 4336 9130 4678 9186
rect 4734 9130 4820 9186
rect 4876 9130 5215 9186
rect 5271 9130 5357 9186
rect 5413 9130 5760 9186
rect 5816 9130 5902 9186
rect 5958 9130 6300 9186
rect 6356 9130 6442 9186
rect 6498 9130 6845 9186
rect 6901 9130 6987 9186
rect 7043 9130 7382 9186
rect 7438 9130 7524 9186
rect 7580 9130 7919 9186
rect 7975 9130 8061 9186
rect 8117 9130 8462 9186
rect 8518 9130 8604 9186
rect 8660 9130 9004 9186
rect 9060 9130 9146 9186
rect 9202 9130 9547 9186
rect 9603 9130 9689 9186
rect 9745 9130 10081 9186
rect 10137 9130 10223 9186
rect 10279 9130 10622 9186
rect 10678 9130 10764 9186
rect 10820 9130 11162 9186
rect 11218 9130 11304 9186
rect 11360 9130 11702 9186
rect 11758 9130 11844 9186
rect 11900 9134 13200 9186
rect 11900 9130 12526 9134
rect 266 9078 12526 9130
rect 12582 9078 12650 9134
rect 12706 9078 12774 9134
rect 12830 9078 12898 9134
rect 12954 9078 13022 9134
rect 13078 9078 13200 9134
rect -400 9044 13200 9078
rect -400 9010 903 9044
rect -400 8954 -286 9010
rect -230 8954 -162 9010
rect -106 8954 -38 9010
rect 18 8954 86 9010
rect 142 8954 210 9010
rect 266 8988 903 9010
rect 959 8988 1045 9044
rect 1101 8988 1444 9044
rect 1500 8988 1586 9044
rect 1642 8988 1984 9044
rect 2040 8988 2126 9044
rect 2182 8988 2521 9044
rect 2577 8988 2663 9044
rect 2719 8988 3058 9044
rect 3114 8988 3200 9044
rect 3256 8988 3602 9044
rect 3658 8988 3744 9044
rect 3800 8988 4138 9044
rect 4194 8988 4280 9044
rect 4336 8988 4678 9044
rect 4734 8988 4820 9044
rect 4876 8988 5215 9044
rect 5271 8988 5357 9044
rect 5413 8988 5760 9044
rect 5816 8988 5902 9044
rect 5958 8988 6300 9044
rect 6356 8988 6442 9044
rect 6498 8988 6845 9044
rect 6901 8988 6987 9044
rect 7043 8988 7382 9044
rect 7438 8988 7524 9044
rect 7580 8988 7919 9044
rect 7975 8988 8061 9044
rect 8117 8988 8462 9044
rect 8518 8988 8604 9044
rect 8660 8988 9004 9044
rect 9060 8988 9146 9044
rect 9202 8988 9547 9044
rect 9603 8988 9689 9044
rect 9745 8988 10081 9044
rect 10137 8988 10223 9044
rect 10279 8988 10622 9044
rect 10678 8988 10764 9044
rect 10820 8988 11162 9044
rect 11218 8988 11304 9044
rect 11360 8988 11702 9044
rect 11758 8988 11844 9044
rect 11900 9010 13200 9044
rect 11900 8988 12526 9010
rect 266 8954 12526 8988
rect 12582 8954 12650 9010
rect 12706 8954 12774 9010
rect 12830 8954 12898 9010
rect 12954 8954 13022 9010
rect 13078 8954 13200 9010
rect -400 8902 13200 8954
rect -400 8886 903 8902
rect -400 8830 -286 8886
rect -230 8830 -162 8886
rect -106 8830 -38 8886
rect 18 8830 86 8886
rect 142 8830 210 8886
rect 266 8846 903 8886
rect 959 8846 1045 8902
rect 1101 8846 1444 8902
rect 1500 8846 1586 8902
rect 1642 8846 1984 8902
rect 2040 8846 2126 8902
rect 2182 8846 2521 8902
rect 2577 8846 2663 8902
rect 2719 8846 3058 8902
rect 3114 8846 3200 8902
rect 3256 8846 3602 8902
rect 3658 8846 3744 8902
rect 3800 8846 4138 8902
rect 4194 8846 4280 8902
rect 4336 8846 4678 8902
rect 4734 8846 4820 8902
rect 4876 8846 5215 8902
rect 5271 8846 5357 8902
rect 5413 8846 5760 8902
rect 5816 8846 5902 8902
rect 5958 8846 6300 8902
rect 6356 8846 6442 8902
rect 6498 8846 6845 8902
rect 6901 8846 6987 8902
rect 7043 8846 7382 8902
rect 7438 8846 7524 8902
rect 7580 8846 7919 8902
rect 7975 8846 8061 8902
rect 8117 8846 8462 8902
rect 8518 8846 8604 8902
rect 8660 8846 9004 8902
rect 9060 8846 9146 8902
rect 9202 8846 9547 8902
rect 9603 8846 9689 8902
rect 9745 8846 10081 8902
rect 10137 8846 10223 8902
rect 10279 8846 10622 8902
rect 10678 8846 10764 8902
rect 10820 8846 11162 8902
rect 11218 8846 11304 8902
rect 11360 8846 11702 8902
rect 11758 8846 11844 8902
rect 11900 8886 13200 8902
rect 11900 8846 12526 8886
rect 266 8830 12526 8846
rect 12582 8830 12650 8886
rect 12706 8830 12774 8886
rect 12830 8830 12898 8886
rect 12954 8830 13022 8886
rect 13078 8830 13200 8886
rect -400 8762 13200 8830
rect -400 8706 -286 8762
rect -230 8706 -162 8762
rect -106 8706 -38 8762
rect 18 8706 86 8762
rect 142 8706 210 8762
rect 266 8760 12526 8762
rect 266 8706 903 8760
rect -400 8704 903 8706
rect 959 8704 1045 8760
rect 1101 8704 1444 8760
rect 1500 8704 1586 8760
rect 1642 8704 1984 8760
rect 2040 8704 2126 8760
rect 2182 8704 2521 8760
rect 2577 8704 2663 8760
rect 2719 8704 3058 8760
rect 3114 8704 3200 8760
rect 3256 8704 3602 8760
rect 3658 8704 3744 8760
rect 3800 8704 4138 8760
rect 4194 8704 4280 8760
rect 4336 8704 4678 8760
rect 4734 8704 4820 8760
rect 4876 8704 5215 8760
rect 5271 8704 5357 8760
rect 5413 8704 5760 8760
rect 5816 8704 5902 8760
rect 5958 8704 6300 8760
rect 6356 8704 6442 8760
rect 6498 8704 6845 8760
rect 6901 8704 6987 8760
rect 7043 8704 7382 8760
rect 7438 8704 7524 8760
rect 7580 8704 7919 8760
rect 7975 8704 8061 8760
rect 8117 8704 8462 8760
rect 8518 8704 8604 8760
rect 8660 8704 9004 8760
rect 9060 8704 9146 8760
rect 9202 8704 9547 8760
rect 9603 8704 9689 8760
rect 9745 8704 10081 8760
rect 10137 8704 10223 8760
rect 10279 8704 10622 8760
rect 10678 8704 10764 8760
rect 10820 8704 11162 8760
rect 11218 8704 11304 8760
rect 11360 8704 11702 8760
rect 11758 8704 11844 8760
rect 11900 8706 12526 8760
rect 12582 8706 12650 8762
rect 12706 8706 12774 8762
rect 12830 8706 12898 8762
rect 12954 8706 13022 8762
rect 13078 8706 13200 8762
rect 11900 8704 13200 8706
rect -400 8638 13200 8704
rect -400 8582 -286 8638
rect -230 8582 -162 8638
rect -106 8582 -38 8638
rect 18 8582 86 8638
rect 142 8582 210 8638
rect 266 8618 12526 8638
rect 266 8582 903 8618
rect -400 8562 903 8582
rect 959 8562 1045 8618
rect 1101 8562 1444 8618
rect 1500 8562 1586 8618
rect 1642 8562 1984 8618
rect 2040 8562 2126 8618
rect 2182 8562 2521 8618
rect 2577 8562 2663 8618
rect 2719 8562 3058 8618
rect 3114 8562 3200 8618
rect 3256 8562 3602 8618
rect 3658 8562 3744 8618
rect 3800 8562 4138 8618
rect 4194 8562 4280 8618
rect 4336 8562 4678 8618
rect 4734 8562 4820 8618
rect 4876 8562 5215 8618
rect 5271 8562 5357 8618
rect 5413 8562 5760 8618
rect 5816 8562 5902 8618
rect 5958 8562 6300 8618
rect 6356 8562 6442 8618
rect 6498 8562 6845 8618
rect 6901 8562 6987 8618
rect 7043 8562 7382 8618
rect 7438 8562 7524 8618
rect 7580 8562 7919 8618
rect 7975 8562 8061 8618
rect 8117 8562 8462 8618
rect 8518 8562 8604 8618
rect 8660 8562 9004 8618
rect 9060 8562 9146 8618
rect 9202 8562 9547 8618
rect 9603 8562 9689 8618
rect 9745 8562 10081 8618
rect 10137 8562 10223 8618
rect 10279 8562 10622 8618
rect 10678 8562 10764 8618
rect 10820 8562 11162 8618
rect 11218 8562 11304 8618
rect 11360 8562 11702 8618
rect 11758 8562 11844 8618
rect 11900 8582 12526 8618
rect 12582 8582 12650 8638
rect 12706 8582 12774 8638
rect 12830 8582 12898 8638
rect 12954 8582 13022 8638
rect 13078 8582 13200 8638
rect 11900 8562 13200 8582
rect -400 8514 13200 8562
rect -400 8458 -286 8514
rect -230 8458 -162 8514
rect -106 8458 -38 8514
rect 18 8458 86 8514
rect 142 8458 210 8514
rect 266 8476 12526 8514
rect 266 8458 903 8476
rect -400 8420 903 8458
rect 959 8420 1045 8476
rect 1101 8420 1444 8476
rect 1500 8420 1586 8476
rect 1642 8420 1984 8476
rect 2040 8420 2126 8476
rect 2182 8420 2521 8476
rect 2577 8420 2663 8476
rect 2719 8420 3058 8476
rect 3114 8420 3200 8476
rect 3256 8420 3602 8476
rect 3658 8420 3744 8476
rect 3800 8420 4138 8476
rect 4194 8420 4280 8476
rect 4336 8420 4678 8476
rect 4734 8420 4820 8476
rect 4876 8420 5215 8476
rect 5271 8420 5357 8476
rect 5413 8420 5760 8476
rect 5816 8420 5902 8476
rect 5958 8420 6300 8476
rect 6356 8420 6442 8476
rect 6498 8420 6845 8476
rect 6901 8420 6987 8476
rect 7043 8420 7382 8476
rect 7438 8420 7524 8476
rect 7580 8420 7919 8476
rect 7975 8420 8061 8476
rect 8117 8420 8462 8476
rect 8518 8420 8604 8476
rect 8660 8420 9004 8476
rect 9060 8420 9146 8476
rect 9202 8420 9547 8476
rect 9603 8420 9689 8476
rect 9745 8420 10081 8476
rect 10137 8420 10223 8476
rect 10279 8420 10622 8476
rect 10678 8420 10764 8476
rect 10820 8420 11162 8476
rect 11218 8420 11304 8476
rect 11360 8420 11702 8476
rect 11758 8420 11844 8476
rect 11900 8458 12526 8476
rect 12582 8458 12650 8514
rect 12706 8458 12774 8514
rect 12830 8458 12898 8514
rect 12954 8458 13022 8514
rect 13078 8458 13200 8514
rect 11900 8420 13200 8458
rect -400 8390 13200 8420
rect -400 8334 -286 8390
rect -230 8334 -162 8390
rect -106 8334 -38 8390
rect 18 8334 86 8390
rect 142 8334 210 8390
rect 266 8334 12526 8390
rect 12582 8334 12650 8390
rect 12706 8334 12774 8390
rect 12830 8334 12898 8390
rect 12954 8334 13022 8390
rect 13078 8334 13200 8390
rect -400 8278 903 8334
rect 959 8278 1045 8334
rect 1101 8278 1444 8334
rect 1500 8278 1586 8334
rect 1642 8278 1984 8334
rect 2040 8278 2126 8334
rect 2182 8278 2521 8334
rect 2577 8278 2663 8334
rect 2719 8278 3058 8334
rect 3114 8278 3200 8334
rect 3256 8278 3602 8334
rect 3658 8278 3744 8334
rect 3800 8278 4138 8334
rect 4194 8278 4280 8334
rect 4336 8278 4678 8334
rect 4734 8278 4820 8334
rect 4876 8278 5215 8334
rect 5271 8278 5357 8334
rect 5413 8278 5760 8334
rect 5816 8278 5902 8334
rect 5958 8278 6300 8334
rect 6356 8278 6442 8334
rect 6498 8278 6845 8334
rect 6901 8278 6987 8334
rect 7043 8278 7382 8334
rect 7438 8278 7524 8334
rect 7580 8278 7919 8334
rect 7975 8278 8061 8334
rect 8117 8278 8462 8334
rect 8518 8278 8604 8334
rect 8660 8278 9004 8334
rect 9060 8278 9146 8334
rect 9202 8278 9547 8334
rect 9603 8278 9689 8334
rect 9745 8278 10081 8334
rect 10137 8278 10223 8334
rect 10279 8278 10622 8334
rect 10678 8278 10764 8334
rect 10820 8278 11162 8334
rect 11218 8278 11304 8334
rect 11360 8278 11702 8334
rect 11758 8278 11844 8334
rect 11900 8278 13200 8334
rect -400 8266 13200 8278
rect -400 8210 -286 8266
rect -230 8210 -162 8266
rect -106 8210 -38 8266
rect 18 8210 86 8266
rect 142 8210 210 8266
rect 266 8210 12526 8266
rect 12582 8210 12650 8266
rect 12706 8210 12774 8266
rect 12830 8210 12898 8266
rect 12954 8210 13022 8266
rect 13078 8210 13200 8266
rect -400 8192 13200 8210
rect -400 8142 903 8192
rect -400 8086 -286 8142
rect -230 8086 -162 8142
rect -106 8086 -38 8142
rect 18 8086 86 8142
rect 142 8086 210 8142
rect 266 8136 903 8142
rect 959 8136 1045 8192
rect 1101 8136 1444 8192
rect 1500 8136 1586 8192
rect 1642 8136 1984 8192
rect 2040 8136 2126 8192
rect 2182 8136 2521 8192
rect 2577 8136 2663 8192
rect 2719 8136 3058 8192
rect 3114 8136 3200 8192
rect 3256 8136 3602 8192
rect 3658 8136 3744 8192
rect 3800 8136 4138 8192
rect 4194 8136 4280 8192
rect 4336 8136 4678 8192
rect 4734 8136 4820 8192
rect 4876 8136 5215 8192
rect 5271 8136 5357 8192
rect 5413 8136 5760 8192
rect 5816 8136 5902 8192
rect 5958 8136 6300 8192
rect 6356 8136 6442 8192
rect 6498 8136 6845 8192
rect 6901 8136 6987 8192
rect 7043 8136 7382 8192
rect 7438 8136 7524 8192
rect 7580 8136 7919 8192
rect 7975 8136 8061 8192
rect 8117 8136 8462 8192
rect 8518 8136 8604 8192
rect 8660 8136 9004 8192
rect 9060 8136 9146 8192
rect 9202 8136 9547 8192
rect 9603 8136 9689 8192
rect 9745 8136 10081 8192
rect 10137 8136 10223 8192
rect 10279 8136 10622 8192
rect 10678 8136 10764 8192
rect 10820 8136 11162 8192
rect 11218 8136 11304 8192
rect 11360 8136 11702 8192
rect 11758 8136 11844 8192
rect 11900 8142 13200 8192
rect 11900 8136 12526 8142
rect 266 8086 12526 8136
rect 12582 8086 12650 8142
rect 12706 8086 12774 8142
rect 12830 8086 12898 8142
rect 12954 8086 13022 8142
rect 13078 8086 13200 8142
rect -400 8050 13200 8086
rect -400 8018 903 8050
rect -400 7962 -286 8018
rect -230 7962 -162 8018
rect -106 7962 -38 8018
rect 18 7962 86 8018
rect 142 7962 210 8018
rect 266 7994 903 8018
rect 959 7994 1045 8050
rect 1101 7994 1444 8050
rect 1500 7994 1586 8050
rect 1642 7994 1984 8050
rect 2040 7994 2126 8050
rect 2182 7994 2521 8050
rect 2577 7994 2663 8050
rect 2719 7994 3058 8050
rect 3114 7994 3200 8050
rect 3256 7994 3602 8050
rect 3658 7994 3744 8050
rect 3800 7994 4138 8050
rect 4194 7994 4280 8050
rect 4336 7994 4678 8050
rect 4734 7994 4820 8050
rect 4876 7994 5215 8050
rect 5271 7994 5357 8050
rect 5413 7994 5760 8050
rect 5816 7994 5902 8050
rect 5958 7994 6300 8050
rect 6356 7994 6442 8050
rect 6498 7994 6845 8050
rect 6901 7994 6987 8050
rect 7043 7994 7382 8050
rect 7438 7994 7524 8050
rect 7580 7994 7919 8050
rect 7975 7994 8061 8050
rect 8117 7994 8462 8050
rect 8518 7994 8604 8050
rect 8660 7994 9004 8050
rect 9060 7994 9146 8050
rect 9202 7994 9547 8050
rect 9603 7994 9689 8050
rect 9745 7994 10081 8050
rect 10137 7994 10223 8050
rect 10279 7994 10622 8050
rect 10678 7994 10764 8050
rect 10820 7994 11162 8050
rect 11218 7994 11304 8050
rect 11360 7994 11702 8050
rect 11758 7994 11844 8050
rect 11900 8018 13200 8050
rect 11900 7994 12526 8018
rect 266 7962 12526 7994
rect 12582 7962 12650 8018
rect 12706 7962 12774 8018
rect 12830 7962 12898 8018
rect 12954 7962 13022 8018
rect 13078 7962 13200 8018
rect -400 7908 13200 7962
rect -400 7894 903 7908
rect -400 7838 -286 7894
rect -230 7838 -162 7894
rect -106 7838 -38 7894
rect 18 7838 86 7894
rect 142 7838 210 7894
rect 266 7852 903 7894
rect 959 7852 1045 7908
rect 1101 7852 1444 7908
rect 1500 7852 1586 7908
rect 1642 7852 1984 7908
rect 2040 7852 2126 7908
rect 2182 7852 2521 7908
rect 2577 7852 2663 7908
rect 2719 7852 3058 7908
rect 3114 7852 3200 7908
rect 3256 7852 3602 7908
rect 3658 7852 3744 7908
rect 3800 7852 4138 7908
rect 4194 7852 4280 7908
rect 4336 7852 4678 7908
rect 4734 7852 4820 7908
rect 4876 7852 5215 7908
rect 5271 7852 5357 7908
rect 5413 7852 5760 7908
rect 5816 7852 5902 7908
rect 5958 7852 6300 7908
rect 6356 7852 6442 7908
rect 6498 7852 6845 7908
rect 6901 7852 6987 7908
rect 7043 7852 7382 7908
rect 7438 7852 7524 7908
rect 7580 7852 7919 7908
rect 7975 7852 8061 7908
rect 8117 7852 8462 7908
rect 8518 7852 8604 7908
rect 8660 7852 9004 7908
rect 9060 7852 9146 7908
rect 9202 7852 9547 7908
rect 9603 7852 9689 7908
rect 9745 7852 10081 7908
rect 10137 7852 10223 7908
rect 10279 7852 10622 7908
rect 10678 7852 10764 7908
rect 10820 7852 11162 7908
rect 11218 7852 11304 7908
rect 11360 7852 11702 7908
rect 11758 7852 11844 7908
rect 11900 7894 13200 7908
rect 11900 7852 12526 7894
rect 266 7838 12526 7852
rect 12582 7838 12650 7894
rect 12706 7838 12774 7894
rect 12830 7838 12898 7894
rect 12954 7838 13022 7894
rect 13078 7838 13200 7894
rect -400 7770 13200 7838
rect -400 7714 -286 7770
rect -230 7714 -162 7770
rect -106 7714 -38 7770
rect 18 7714 86 7770
rect 142 7714 210 7770
rect 266 7766 12526 7770
rect 266 7714 903 7766
rect -400 7710 903 7714
rect 959 7710 1045 7766
rect 1101 7710 1444 7766
rect 1500 7710 1586 7766
rect 1642 7710 1984 7766
rect 2040 7710 2126 7766
rect 2182 7710 2521 7766
rect 2577 7710 2663 7766
rect 2719 7710 3058 7766
rect 3114 7710 3200 7766
rect 3256 7710 3602 7766
rect 3658 7710 3744 7766
rect 3800 7710 4138 7766
rect 4194 7710 4280 7766
rect 4336 7710 4678 7766
rect 4734 7710 4820 7766
rect 4876 7710 5215 7766
rect 5271 7710 5357 7766
rect 5413 7710 5760 7766
rect 5816 7710 5902 7766
rect 5958 7710 6300 7766
rect 6356 7710 6442 7766
rect 6498 7710 6845 7766
rect 6901 7710 6987 7766
rect 7043 7710 7382 7766
rect 7438 7710 7524 7766
rect 7580 7710 7919 7766
rect 7975 7710 8061 7766
rect 8117 7710 8462 7766
rect 8518 7710 8604 7766
rect 8660 7710 9004 7766
rect 9060 7710 9146 7766
rect 9202 7710 9547 7766
rect 9603 7710 9689 7766
rect 9745 7710 10081 7766
rect 10137 7710 10223 7766
rect 10279 7710 10622 7766
rect 10678 7710 10764 7766
rect 10820 7710 11162 7766
rect 11218 7710 11304 7766
rect 11360 7710 11702 7766
rect 11758 7710 11844 7766
rect 11900 7714 12526 7766
rect 12582 7714 12650 7770
rect 12706 7714 12774 7770
rect 12830 7714 12898 7770
rect 12954 7714 13022 7770
rect 13078 7714 13200 7770
rect 11900 7710 13200 7714
rect -400 7646 13200 7710
rect -400 7590 -286 7646
rect -230 7590 -162 7646
rect -106 7590 -38 7646
rect 18 7590 86 7646
rect 142 7590 210 7646
rect 266 7624 12526 7646
rect 266 7590 903 7624
rect -400 7568 903 7590
rect 959 7568 1045 7624
rect 1101 7568 1444 7624
rect 1500 7568 1586 7624
rect 1642 7568 1984 7624
rect 2040 7568 2126 7624
rect 2182 7568 2521 7624
rect 2577 7568 2663 7624
rect 2719 7568 3058 7624
rect 3114 7568 3200 7624
rect 3256 7568 3602 7624
rect 3658 7568 3744 7624
rect 3800 7568 4138 7624
rect 4194 7568 4280 7624
rect 4336 7568 4678 7624
rect 4734 7568 4820 7624
rect 4876 7568 5215 7624
rect 5271 7568 5357 7624
rect 5413 7568 5760 7624
rect 5816 7568 5902 7624
rect 5958 7568 6300 7624
rect 6356 7568 6442 7624
rect 6498 7568 6845 7624
rect 6901 7568 6987 7624
rect 7043 7568 7382 7624
rect 7438 7568 7524 7624
rect 7580 7568 7919 7624
rect 7975 7568 8061 7624
rect 8117 7568 8462 7624
rect 8518 7568 8604 7624
rect 8660 7568 9004 7624
rect 9060 7568 9146 7624
rect 9202 7568 9547 7624
rect 9603 7568 9689 7624
rect 9745 7568 10081 7624
rect 10137 7568 10223 7624
rect 10279 7568 10622 7624
rect 10678 7568 10764 7624
rect 10820 7568 11162 7624
rect 11218 7568 11304 7624
rect 11360 7568 11702 7624
rect 11758 7568 11844 7624
rect 11900 7590 12526 7624
rect 12582 7590 12650 7646
rect 12706 7590 12774 7646
rect 12830 7590 12898 7646
rect 12954 7590 13022 7646
rect 13078 7590 13200 7646
rect 11900 7568 13200 7590
rect -400 7522 13200 7568
rect -400 7466 -286 7522
rect -230 7466 -162 7522
rect -106 7466 -38 7522
rect 18 7466 86 7522
rect 142 7466 210 7522
rect 266 7482 12526 7522
rect 266 7466 903 7482
rect -400 7426 903 7466
rect 959 7426 1045 7482
rect 1101 7426 1444 7482
rect 1500 7426 1586 7482
rect 1642 7426 1984 7482
rect 2040 7426 2126 7482
rect 2182 7426 2521 7482
rect 2577 7426 2663 7482
rect 2719 7426 3058 7482
rect 3114 7426 3200 7482
rect 3256 7426 3602 7482
rect 3658 7426 3744 7482
rect 3800 7426 4138 7482
rect 4194 7426 4280 7482
rect 4336 7426 4678 7482
rect 4734 7426 4820 7482
rect 4876 7426 5215 7482
rect 5271 7426 5357 7482
rect 5413 7426 5760 7482
rect 5816 7426 5902 7482
rect 5958 7426 6300 7482
rect 6356 7426 6442 7482
rect 6498 7426 6845 7482
rect 6901 7426 6987 7482
rect 7043 7426 7382 7482
rect 7438 7426 7524 7482
rect 7580 7426 7919 7482
rect 7975 7426 8061 7482
rect 8117 7426 8462 7482
rect 8518 7426 8604 7482
rect 8660 7426 9004 7482
rect 9060 7426 9146 7482
rect 9202 7426 9547 7482
rect 9603 7426 9689 7482
rect 9745 7426 10081 7482
rect 10137 7426 10223 7482
rect 10279 7426 10622 7482
rect 10678 7426 10764 7482
rect 10820 7426 11162 7482
rect 11218 7426 11304 7482
rect 11360 7426 11702 7482
rect 11758 7426 11844 7482
rect 11900 7466 12526 7482
rect 12582 7466 12650 7522
rect 12706 7466 12774 7522
rect 12830 7466 12898 7522
rect 12954 7466 13022 7522
rect 13078 7466 13200 7522
rect 11900 7426 13200 7466
rect -400 7398 13200 7426
rect -400 7342 -286 7398
rect -230 7342 -162 7398
rect -106 7342 -38 7398
rect 18 7342 86 7398
rect 142 7342 210 7398
rect 266 7342 12526 7398
rect 12582 7342 12650 7398
rect 12706 7342 12774 7398
rect 12830 7342 12898 7398
rect 12954 7342 13022 7398
rect 13078 7342 13200 7398
rect -400 7340 13200 7342
rect -400 7284 903 7340
rect 959 7284 1045 7340
rect 1101 7284 1444 7340
rect 1500 7284 1586 7340
rect 1642 7284 1984 7340
rect 2040 7284 2126 7340
rect 2182 7284 2521 7340
rect 2577 7284 2663 7340
rect 2719 7284 3058 7340
rect 3114 7284 3200 7340
rect 3256 7284 3602 7340
rect 3658 7284 3744 7340
rect 3800 7284 4138 7340
rect 4194 7284 4280 7340
rect 4336 7284 4678 7340
rect 4734 7284 4820 7340
rect 4876 7284 5215 7340
rect 5271 7284 5357 7340
rect 5413 7284 5760 7340
rect 5816 7284 5902 7340
rect 5958 7284 6300 7340
rect 6356 7284 6442 7340
rect 6498 7284 6845 7340
rect 6901 7284 6987 7340
rect 7043 7284 7382 7340
rect 7438 7284 7524 7340
rect 7580 7284 7919 7340
rect 7975 7284 8061 7340
rect 8117 7284 8462 7340
rect 8518 7284 8604 7340
rect 8660 7284 9004 7340
rect 9060 7284 9146 7340
rect 9202 7284 9547 7340
rect 9603 7284 9689 7340
rect 9745 7284 10081 7340
rect 10137 7284 10223 7340
rect 10279 7284 10622 7340
rect 10678 7284 10764 7340
rect 10820 7284 11162 7340
rect 11218 7284 11304 7340
rect 11360 7284 11702 7340
rect 11758 7284 11844 7340
rect 11900 7284 13200 7340
rect -400 7274 13200 7284
rect -400 7218 -286 7274
rect -230 7218 -162 7274
rect -106 7218 -38 7274
rect 18 7218 86 7274
rect 142 7218 210 7274
rect 266 7218 12526 7274
rect 12582 7218 12650 7274
rect 12706 7218 12774 7274
rect 12830 7218 12898 7274
rect 12954 7218 13022 7274
rect 13078 7218 13200 7274
rect -400 7198 13200 7218
rect -400 7150 903 7198
rect -400 7094 -286 7150
rect -230 7094 -162 7150
rect -106 7094 -38 7150
rect 18 7094 86 7150
rect 142 7094 210 7150
rect 266 7142 903 7150
rect 959 7142 1045 7198
rect 1101 7142 1444 7198
rect 1500 7142 1586 7198
rect 1642 7142 1984 7198
rect 2040 7142 2126 7198
rect 2182 7142 2521 7198
rect 2577 7142 2663 7198
rect 2719 7142 3058 7198
rect 3114 7142 3200 7198
rect 3256 7142 3602 7198
rect 3658 7142 3744 7198
rect 3800 7142 4138 7198
rect 4194 7142 4280 7198
rect 4336 7142 4678 7198
rect 4734 7142 4820 7198
rect 4876 7142 5215 7198
rect 5271 7142 5357 7198
rect 5413 7142 5760 7198
rect 5816 7142 5902 7198
rect 5958 7142 6300 7198
rect 6356 7142 6442 7198
rect 6498 7142 6845 7198
rect 6901 7142 6987 7198
rect 7043 7142 7382 7198
rect 7438 7142 7524 7198
rect 7580 7142 7919 7198
rect 7975 7142 8061 7198
rect 8117 7142 8462 7198
rect 8518 7142 8604 7198
rect 8660 7142 9004 7198
rect 9060 7142 9146 7198
rect 9202 7142 9547 7198
rect 9603 7142 9689 7198
rect 9745 7142 10081 7198
rect 10137 7142 10223 7198
rect 10279 7142 10622 7198
rect 10678 7142 10764 7198
rect 10820 7142 11162 7198
rect 11218 7142 11304 7198
rect 11360 7142 11702 7198
rect 11758 7142 11844 7198
rect 11900 7150 13200 7198
rect 11900 7142 12526 7150
rect 266 7094 12526 7142
rect 12582 7094 12650 7150
rect 12706 7094 12774 7150
rect 12830 7094 12898 7150
rect 12954 7094 13022 7150
rect 13078 7094 13200 7150
rect -400 7056 13200 7094
rect -400 7026 903 7056
rect -400 6970 -286 7026
rect -230 6970 -162 7026
rect -106 6970 -38 7026
rect 18 6970 86 7026
rect 142 6970 210 7026
rect 266 7000 903 7026
rect 959 7000 1045 7056
rect 1101 7000 1444 7056
rect 1500 7000 1586 7056
rect 1642 7000 1984 7056
rect 2040 7000 2126 7056
rect 2182 7000 2521 7056
rect 2577 7000 2663 7056
rect 2719 7000 3058 7056
rect 3114 7000 3200 7056
rect 3256 7000 3602 7056
rect 3658 7000 3744 7056
rect 3800 7000 4138 7056
rect 4194 7000 4280 7056
rect 4336 7000 4678 7056
rect 4734 7000 4820 7056
rect 4876 7000 5215 7056
rect 5271 7000 5357 7056
rect 5413 7000 5760 7056
rect 5816 7000 5902 7056
rect 5958 7000 6300 7056
rect 6356 7000 6442 7056
rect 6498 7000 6845 7056
rect 6901 7000 6987 7056
rect 7043 7000 7382 7056
rect 7438 7000 7524 7056
rect 7580 7000 7919 7056
rect 7975 7000 8061 7056
rect 8117 7000 8462 7056
rect 8518 7000 8604 7056
rect 8660 7000 9004 7056
rect 9060 7000 9146 7056
rect 9202 7000 9547 7056
rect 9603 7000 9689 7056
rect 9745 7000 10081 7056
rect 10137 7000 10223 7056
rect 10279 7000 10622 7056
rect 10678 7000 10764 7056
rect 10820 7000 11162 7056
rect 11218 7000 11304 7056
rect 11360 7000 11702 7056
rect 11758 7000 11844 7056
rect 11900 7026 13200 7056
rect 11900 7000 12526 7026
rect 266 6970 12526 7000
rect 12582 6970 12650 7026
rect 12706 6970 12774 7026
rect 12830 6970 12898 7026
rect 12954 6970 13022 7026
rect 13078 6970 13200 7026
rect -400 6914 13200 6970
rect -400 6902 903 6914
rect -400 6846 -286 6902
rect -230 6846 -162 6902
rect -106 6846 -38 6902
rect 18 6846 86 6902
rect 142 6846 210 6902
rect 266 6858 903 6902
rect 959 6858 1045 6914
rect 1101 6858 1444 6914
rect 1500 6858 1586 6914
rect 1642 6858 1984 6914
rect 2040 6858 2126 6914
rect 2182 6858 2521 6914
rect 2577 6858 2663 6914
rect 2719 6858 3058 6914
rect 3114 6858 3200 6914
rect 3256 6858 3602 6914
rect 3658 6858 3744 6914
rect 3800 6858 4138 6914
rect 4194 6858 4280 6914
rect 4336 6858 4678 6914
rect 4734 6858 4820 6914
rect 4876 6858 5215 6914
rect 5271 6858 5357 6914
rect 5413 6858 5760 6914
rect 5816 6858 5902 6914
rect 5958 6858 6300 6914
rect 6356 6858 6442 6914
rect 6498 6858 6845 6914
rect 6901 6858 6987 6914
rect 7043 6858 7382 6914
rect 7438 6858 7524 6914
rect 7580 6858 7919 6914
rect 7975 6858 8061 6914
rect 8117 6858 8462 6914
rect 8518 6858 8604 6914
rect 8660 6858 9004 6914
rect 9060 6858 9146 6914
rect 9202 6858 9547 6914
rect 9603 6858 9689 6914
rect 9745 6858 10081 6914
rect 10137 6858 10223 6914
rect 10279 6858 10622 6914
rect 10678 6858 10764 6914
rect 10820 6858 11162 6914
rect 11218 6858 11304 6914
rect 11360 6858 11702 6914
rect 11758 6858 11844 6914
rect 11900 6902 13200 6914
rect 11900 6858 12526 6902
rect 266 6846 12526 6858
rect 12582 6846 12650 6902
rect 12706 6846 12774 6902
rect 12830 6846 12898 6902
rect 12954 6846 13022 6902
rect 13078 6846 13200 6902
rect -400 6778 13200 6846
rect -400 6722 -286 6778
rect -230 6722 -162 6778
rect -106 6722 -38 6778
rect 18 6722 86 6778
rect 142 6722 210 6778
rect 266 6772 12526 6778
rect 266 6722 903 6772
rect -400 6716 903 6722
rect 959 6716 1045 6772
rect 1101 6716 1444 6772
rect 1500 6716 1586 6772
rect 1642 6716 1984 6772
rect 2040 6716 2126 6772
rect 2182 6716 2521 6772
rect 2577 6716 2663 6772
rect 2719 6716 3058 6772
rect 3114 6716 3200 6772
rect 3256 6716 3602 6772
rect 3658 6716 3744 6772
rect 3800 6716 4138 6772
rect 4194 6716 4280 6772
rect 4336 6716 4678 6772
rect 4734 6716 4820 6772
rect 4876 6716 5215 6772
rect 5271 6716 5357 6772
rect 5413 6716 5760 6772
rect 5816 6716 5902 6772
rect 5958 6716 6300 6772
rect 6356 6716 6442 6772
rect 6498 6716 6845 6772
rect 6901 6716 6987 6772
rect 7043 6716 7382 6772
rect 7438 6716 7524 6772
rect 7580 6716 7919 6772
rect 7975 6716 8061 6772
rect 8117 6716 8462 6772
rect 8518 6716 8604 6772
rect 8660 6716 9004 6772
rect 9060 6716 9146 6772
rect 9202 6716 9547 6772
rect 9603 6716 9689 6772
rect 9745 6716 10081 6772
rect 10137 6716 10223 6772
rect 10279 6716 10622 6772
rect 10678 6716 10764 6772
rect 10820 6716 11162 6772
rect 11218 6716 11304 6772
rect 11360 6716 11702 6772
rect 11758 6716 11844 6772
rect 11900 6722 12526 6772
rect 12582 6722 12650 6778
rect 12706 6722 12774 6778
rect 12830 6722 12898 6778
rect 12954 6722 13022 6778
rect 13078 6722 13200 6778
rect 11900 6716 13200 6722
rect -400 6654 13200 6716
rect -400 6598 -286 6654
rect -230 6598 -162 6654
rect -106 6598 -38 6654
rect 18 6598 86 6654
rect 142 6598 210 6654
rect 266 6630 12526 6654
rect 266 6598 903 6630
rect -400 6574 903 6598
rect 959 6574 1045 6630
rect 1101 6574 1444 6630
rect 1500 6574 1586 6630
rect 1642 6574 1984 6630
rect 2040 6574 2126 6630
rect 2182 6574 2521 6630
rect 2577 6574 2663 6630
rect 2719 6574 3058 6630
rect 3114 6574 3200 6630
rect 3256 6574 3602 6630
rect 3658 6574 3744 6630
rect 3800 6574 4138 6630
rect 4194 6574 4280 6630
rect 4336 6574 4678 6630
rect 4734 6574 4820 6630
rect 4876 6574 5215 6630
rect 5271 6574 5357 6630
rect 5413 6574 5760 6630
rect 5816 6574 5902 6630
rect 5958 6574 6300 6630
rect 6356 6574 6442 6630
rect 6498 6574 6845 6630
rect 6901 6574 6987 6630
rect 7043 6574 7382 6630
rect 7438 6574 7524 6630
rect 7580 6574 7919 6630
rect 7975 6574 8061 6630
rect 8117 6574 8462 6630
rect 8518 6574 8604 6630
rect 8660 6574 9004 6630
rect 9060 6574 9146 6630
rect 9202 6574 9547 6630
rect 9603 6574 9689 6630
rect 9745 6574 10081 6630
rect 10137 6574 10223 6630
rect 10279 6574 10622 6630
rect 10678 6574 10764 6630
rect 10820 6574 11162 6630
rect 11218 6574 11304 6630
rect 11360 6574 11702 6630
rect 11758 6574 11844 6630
rect 11900 6598 12526 6630
rect 12582 6598 12650 6654
rect 12706 6598 12774 6654
rect 12830 6598 12898 6654
rect 12954 6598 13022 6654
rect 13078 6598 13200 6654
rect 11900 6574 13200 6598
rect -400 6530 13200 6574
rect -400 6474 -286 6530
rect -230 6474 -162 6530
rect -106 6474 -38 6530
rect 18 6474 86 6530
rect 142 6474 210 6530
rect 266 6488 12526 6530
rect 266 6474 903 6488
rect -400 6432 903 6474
rect 959 6432 1045 6488
rect 1101 6432 1444 6488
rect 1500 6432 1586 6488
rect 1642 6432 1984 6488
rect 2040 6432 2126 6488
rect 2182 6432 2521 6488
rect 2577 6432 2663 6488
rect 2719 6432 3058 6488
rect 3114 6432 3200 6488
rect 3256 6432 3602 6488
rect 3658 6432 3744 6488
rect 3800 6432 4138 6488
rect 4194 6432 4280 6488
rect 4336 6432 4678 6488
rect 4734 6432 4820 6488
rect 4876 6432 5215 6488
rect 5271 6432 5357 6488
rect 5413 6432 5760 6488
rect 5816 6432 5902 6488
rect 5958 6432 6300 6488
rect 6356 6432 6442 6488
rect 6498 6432 6845 6488
rect 6901 6432 6987 6488
rect 7043 6432 7382 6488
rect 7438 6432 7524 6488
rect 7580 6432 7919 6488
rect 7975 6432 8061 6488
rect 8117 6432 8462 6488
rect 8518 6432 8604 6488
rect 8660 6432 9004 6488
rect 9060 6432 9146 6488
rect 9202 6432 9547 6488
rect 9603 6432 9689 6488
rect 9745 6432 10081 6488
rect 10137 6432 10223 6488
rect 10279 6432 10622 6488
rect 10678 6432 10764 6488
rect 10820 6432 11162 6488
rect 11218 6432 11304 6488
rect 11360 6432 11702 6488
rect 11758 6432 11844 6488
rect 11900 6474 12526 6488
rect 12582 6474 12650 6530
rect 12706 6474 12774 6530
rect 12830 6474 12898 6530
rect 12954 6474 13022 6530
rect 13078 6474 13200 6530
rect 11900 6432 13200 6474
rect -400 6406 13200 6432
rect -400 6350 -286 6406
rect -230 6350 -162 6406
rect -106 6350 -38 6406
rect 18 6350 86 6406
rect 142 6350 210 6406
rect 266 6350 12526 6406
rect 12582 6350 12650 6406
rect 12706 6350 12774 6406
rect 12830 6350 12898 6406
rect 12954 6350 13022 6406
rect 13078 6350 13200 6406
rect -400 6346 13200 6350
rect -400 6290 903 6346
rect 959 6290 1045 6346
rect 1101 6290 1444 6346
rect 1500 6290 1586 6346
rect 1642 6290 1984 6346
rect 2040 6290 2126 6346
rect 2182 6290 2521 6346
rect 2577 6290 2663 6346
rect 2719 6290 3058 6346
rect 3114 6290 3200 6346
rect 3256 6290 3602 6346
rect 3658 6290 3744 6346
rect 3800 6290 4138 6346
rect 4194 6290 4280 6346
rect 4336 6290 4678 6346
rect 4734 6290 4820 6346
rect 4876 6290 5215 6346
rect 5271 6290 5357 6346
rect 5413 6290 5760 6346
rect 5816 6290 5902 6346
rect 5958 6290 6300 6346
rect 6356 6290 6442 6346
rect 6498 6290 6845 6346
rect 6901 6290 6987 6346
rect 7043 6290 7382 6346
rect 7438 6290 7524 6346
rect 7580 6290 7919 6346
rect 7975 6290 8061 6346
rect 8117 6290 8462 6346
rect 8518 6290 8604 6346
rect 8660 6290 9004 6346
rect 9060 6290 9146 6346
rect 9202 6290 9547 6346
rect 9603 6290 9689 6346
rect 9745 6290 10081 6346
rect 10137 6290 10223 6346
rect 10279 6290 10622 6346
rect 10678 6290 10764 6346
rect 10820 6290 11162 6346
rect 11218 6290 11304 6346
rect 11360 6290 11702 6346
rect 11758 6290 11844 6346
rect 11900 6290 13200 6346
rect -400 6282 13200 6290
rect -400 6226 -286 6282
rect -230 6226 -162 6282
rect -106 6226 -38 6282
rect 18 6226 86 6282
rect 142 6226 210 6282
rect 266 6226 12526 6282
rect 12582 6226 12650 6282
rect 12706 6226 12774 6282
rect 12830 6226 12898 6282
rect 12954 6226 13022 6282
rect 13078 6226 13200 6282
rect -400 6204 13200 6226
rect -400 6158 903 6204
rect -400 6102 -286 6158
rect -230 6102 -162 6158
rect -106 6102 -38 6158
rect 18 6102 86 6158
rect 142 6102 210 6158
rect 266 6148 903 6158
rect 959 6148 1045 6204
rect 1101 6148 1444 6204
rect 1500 6148 1586 6204
rect 1642 6148 1984 6204
rect 2040 6148 2126 6204
rect 2182 6148 2521 6204
rect 2577 6148 2663 6204
rect 2719 6148 3058 6204
rect 3114 6148 3200 6204
rect 3256 6148 3602 6204
rect 3658 6148 3744 6204
rect 3800 6148 4138 6204
rect 4194 6148 4280 6204
rect 4336 6148 4678 6204
rect 4734 6148 4820 6204
rect 4876 6148 5215 6204
rect 5271 6148 5357 6204
rect 5413 6148 5760 6204
rect 5816 6148 5902 6204
rect 5958 6148 6300 6204
rect 6356 6148 6442 6204
rect 6498 6148 6845 6204
rect 6901 6148 6987 6204
rect 7043 6148 7382 6204
rect 7438 6148 7524 6204
rect 7580 6148 7919 6204
rect 7975 6148 8061 6204
rect 8117 6148 8462 6204
rect 8518 6148 8604 6204
rect 8660 6148 9004 6204
rect 9060 6148 9146 6204
rect 9202 6148 9547 6204
rect 9603 6148 9689 6204
rect 9745 6148 10081 6204
rect 10137 6148 10223 6204
rect 10279 6148 10622 6204
rect 10678 6148 10764 6204
rect 10820 6148 11162 6204
rect 11218 6148 11304 6204
rect 11360 6148 11702 6204
rect 11758 6148 11844 6204
rect 11900 6158 13200 6204
rect 11900 6148 12526 6158
rect 266 6102 12526 6148
rect 12582 6102 12650 6158
rect 12706 6102 12774 6158
rect 12830 6102 12898 6158
rect 12954 6102 13022 6158
rect 13078 6102 13200 6158
rect -400 6062 13200 6102
rect -400 6034 903 6062
rect -400 5978 -286 6034
rect -230 5978 -162 6034
rect -106 5978 -38 6034
rect 18 5978 86 6034
rect 142 5978 210 6034
rect 266 6006 903 6034
rect 959 6006 1045 6062
rect 1101 6006 1444 6062
rect 1500 6006 1586 6062
rect 1642 6006 1984 6062
rect 2040 6006 2126 6062
rect 2182 6006 2521 6062
rect 2577 6006 2663 6062
rect 2719 6006 3058 6062
rect 3114 6006 3200 6062
rect 3256 6006 3602 6062
rect 3658 6006 3744 6062
rect 3800 6006 4138 6062
rect 4194 6006 4280 6062
rect 4336 6006 4678 6062
rect 4734 6006 4820 6062
rect 4876 6006 5215 6062
rect 5271 6006 5357 6062
rect 5413 6006 5760 6062
rect 5816 6006 5902 6062
rect 5958 6006 6300 6062
rect 6356 6006 6442 6062
rect 6498 6006 6845 6062
rect 6901 6006 6987 6062
rect 7043 6006 7382 6062
rect 7438 6006 7524 6062
rect 7580 6006 7919 6062
rect 7975 6006 8061 6062
rect 8117 6006 8462 6062
rect 8518 6006 8604 6062
rect 8660 6006 9004 6062
rect 9060 6006 9146 6062
rect 9202 6006 9547 6062
rect 9603 6006 9689 6062
rect 9745 6006 10081 6062
rect 10137 6006 10223 6062
rect 10279 6006 10622 6062
rect 10678 6006 10764 6062
rect 10820 6006 11162 6062
rect 11218 6006 11304 6062
rect 11360 6006 11702 6062
rect 11758 6006 11844 6062
rect 11900 6034 13200 6062
rect 11900 6006 12526 6034
rect 266 5978 12526 6006
rect 12582 5978 12650 6034
rect 12706 5978 12774 6034
rect 12830 5978 12898 6034
rect 12954 5978 13022 6034
rect 13078 5978 13200 6034
rect -400 5920 13200 5978
rect -400 5910 903 5920
rect -400 5854 -286 5910
rect -230 5854 -162 5910
rect -106 5854 -38 5910
rect 18 5854 86 5910
rect 142 5854 210 5910
rect 266 5864 903 5910
rect 959 5864 1045 5920
rect 1101 5864 1444 5920
rect 1500 5864 1586 5920
rect 1642 5864 1984 5920
rect 2040 5864 2126 5920
rect 2182 5864 2521 5920
rect 2577 5864 2663 5920
rect 2719 5864 3058 5920
rect 3114 5864 3200 5920
rect 3256 5864 3602 5920
rect 3658 5864 3744 5920
rect 3800 5864 4138 5920
rect 4194 5864 4280 5920
rect 4336 5864 4678 5920
rect 4734 5864 4820 5920
rect 4876 5864 5215 5920
rect 5271 5864 5357 5920
rect 5413 5864 5760 5920
rect 5816 5864 5902 5920
rect 5958 5864 6300 5920
rect 6356 5864 6442 5920
rect 6498 5864 6845 5920
rect 6901 5864 6987 5920
rect 7043 5864 7382 5920
rect 7438 5864 7524 5920
rect 7580 5864 7919 5920
rect 7975 5864 8061 5920
rect 8117 5864 8462 5920
rect 8518 5864 8604 5920
rect 8660 5864 9004 5920
rect 9060 5864 9146 5920
rect 9202 5864 9547 5920
rect 9603 5864 9689 5920
rect 9745 5864 10081 5920
rect 10137 5864 10223 5920
rect 10279 5864 10622 5920
rect 10678 5864 10764 5920
rect 10820 5864 11162 5920
rect 11218 5864 11304 5920
rect 11360 5864 11702 5920
rect 11758 5864 11844 5920
rect 11900 5910 13200 5920
rect 11900 5864 12526 5910
rect 266 5854 12526 5864
rect 12582 5854 12650 5910
rect 12706 5854 12774 5910
rect 12830 5854 12898 5910
rect 12954 5854 13022 5910
rect 13078 5854 13200 5910
rect -400 5786 13200 5854
rect -400 5730 -286 5786
rect -230 5730 -162 5786
rect -106 5730 -38 5786
rect 18 5730 86 5786
rect 142 5730 210 5786
rect 266 5778 12526 5786
rect 266 5730 903 5778
rect -400 5722 903 5730
rect 959 5722 1045 5778
rect 1101 5722 1444 5778
rect 1500 5722 1586 5778
rect 1642 5722 1984 5778
rect 2040 5722 2126 5778
rect 2182 5722 2521 5778
rect 2577 5722 2663 5778
rect 2719 5722 3058 5778
rect 3114 5722 3200 5778
rect 3256 5722 3602 5778
rect 3658 5722 3744 5778
rect 3800 5722 4138 5778
rect 4194 5722 4280 5778
rect 4336 5722 4678 5778
rect 4734 5722 4820 5778
rect 4876 5722 5215 5778
rect 5271 5722 5357 5778
rect 5413 5722 5760 5778
rect 5816 5722 5902 5778
rect 5958 5722 6300 5778
rect 6356 5722 6442 5778
rect 6498 5722 6845 5778
rect 6901 5722 6987 5778
rect 7043 5722 7382 5778
rect 7438 5722 7524 5778
rect 7580 5722 7919 5778
rect 7975 5722 8061 5778
rect 8117 5722 8462 5778
rect 8518 5722 8604 5778
rect 8660 5722 9004 5778
rect 9060 5722 9146 5778
rect 9202 5722 9547 5778
rect 9603 5722 9689 5778
rect 9745 5722 10081 5778
rect 10137 5722 10223 5778
rect 10279 5722 10622 5778
rect 10678 5722 10764 5778
rect 10820 5722 11162 5778
rect 11218 5722 11304 5778
rect 11360 5722 11702 5778
rect 11758 5722 11844 5778
rect 11900 5730 12526 5778
rect 12582 5730 12650 5786
rect 12706 5730 12774 5786
rect 12830 5730 12898 5786
rect 12954 5730 13022 5786
rect 13078 5730 13200 5786
rect 11900 5722 13200 5730
rect -400 5662 13200 5722
rect -400 5606 -286 5662
rect -230 5606 -162 5662
rect -106 5606 -38 5662
rect 18 5606 86 5662
rect 142 5606 210 5662
rect 266 5636 12526 5662
rect 266 5606 903 5636
rect -400 5580 903 5606
rect 959 5580 1045 5636
rect 1101 5580 1444 5636
rect 1500 5580 1586 5636
rect 1642 5580 1984 5636
rect 2040 5580 2126 5636
rect 2182 5580 2521 5636
rect 2577 5580 2663 5636
rect 2719 5580 3058 5636
rect 3114 5580 3200 5636
rect 3256 5580 3602 5636
rect 3658 5580 3744 5636
rect 3800 5580 4138 5636
rect 4194 5580 4280 5636
rect 4336 5580 4678 5636
rect 4734 5580 4820 5636
rect 4876 5580 5215 5636
rect 5271 5580 5357 5636
rect 5413 5580 5760 5636
rect 5816 5580 5902 5636
rect 5958 5580 6300 5636
rect 6356 5580 6442 5636
rect 6498 5580 6845 5636
rect 6901 5580 6987 5636
rect 7043 5580 7382 5636
rect 7438 5580 7524 5636
rect 7580 5580 7919 5636
rect 7975 5580 8061 5636
rect 8117 5580 8462 5636
rect 8518 5580 8604 5636
rect 8660 5580 9004 5636
rect 9060 5580 9146 5636
rect 9202 5580 9547 5636
rect 9603 5580 9689 5636
rect 9745 5580 10081 5636
rect 10137 5580 10223 5636
rect 10279 5580 10622 5636
rect 10678 5580 10764 5636
rect 10820 5580 11162 5636
rect 11218 5580 11304 5636
rect 11360 5580 11702 5636
rect 11758 5580 11844 5636
rect 11900 5606 12526 5636
rect 12582 5606 12650 5662
rect 12706 5606 12774 5662
rect 12830 5606 12898 5662
rect 12954 5606 13022 5662
rect 13078 5606 13200 5662
rect 11900 5580 13200 5606
rect -400 5538 13200 5580
rect -400 5482 -286 5538
rect -230 5482 -162 5538
rect -106 5482 -38 5538
rect 18 5482 86 5538
rect 142 5482 210 5538
rect 266 5494 12526 5538
rect 266 5482 903 5494
rect -400 5438 903 5482
rect 959 5438 1045 5494
rect 1101 5438 1444 5494
rect 1500 5438 1586 5494
rect 1642 5438 1984 5494
rect 2040 5438 2126 5494
rect 2182 5438 2521 5494
rect 2577 5438 2663 5494
rect 2719 5438 3058 5494
rect 3114 5438 3200 5494
rect 3256 5438 3602 5494
rect 3658 5438 3744 5494
rect 3800 5438 4138 5494
rect 4194 5438 4280 5494
rect 4336 5438 4678 5494
rect 4734 5438 4820 5494
rect 4876 5438 5215 5494
rect 5271 5438 5357 5494
rect 5413 5438 5760 5494
rect 5816 5438 5902 5494
rect 5958 5438 6300 5494
rect 6356 5438 6442 5494
rect 6498 5438 6845 5494
rect 6901 5438 6987 5494
rect 7043 5438 7382 5494
rect 7438 5438 7524 5494
rect 7580 5438 7919 5494
rect 7975 5438 8061 5494
rect 8117 5438 8462 5494
rect 8518 5438 8604 5494
rect 8660 5438 9004 5494
rect 9060 5438 9146 5494
rect 9202 5438 9547 5494
rect 9603 5438 9689 5494
rect 9745 5438 10081 5494
rect 10137 5438 10223 5494
rect 10279 5438 10622 5494
rect 10678 5438 10764 5494
rect 10820 5438 11162 5494
rect 11218 5438 11304 5494
rect 11360 5438 11702 5494
rect 11758 5438 11844 5494
rect 11900 5482 12526 5494
rect 12582 5482 12650 5538
rect 12706 5482 12774 5538
rect 12830 5482 12898 5538
rect 12954 5482 13022 5538
rect 13078 5482 13200 5538
rect 11900 5438 13200 5482
rect -400 5414 13200 5438
rect -400 5358 -286 5414
rect -230 5358 -162 5414
rect -106 5358 -38 5414
rect 18 5358 86 5414
rect 142 5358 210 5414
rect 266 5358 12526 5414
rect 12582 5358 12650 5414
rect 12706 5358 12774 5414
rect 12830 5358 12898 5414
rect 12954 5358 13022 5414
rect 13078 5358 13200 5414
rect -400 5352 13200 5358
rect -400 5296 903 5352
rect 959 5296 1045 5352
rect 1101 5296 1444 5352
rect 1500 5296 1586 5352
rect 1642 5296 1984 5352
rect 2040 5296 2126 5352
rect 2182 5296 2521 5352
rect 2577 5296 2663 5352
rect 2719 5296 3058 5352
rect 3114 5296 3200 5352
rect 3256 5296 3602 5352
rect 3658 5296 3744 5352
rect 3800 5296 4138 5352
rect 4194 5296 4280 5352
rect 4336 5296 4678 5352
rect 4734 5296 4820 5352
rect 4876 5296 5215 5352
rect 5271 5296 5357 5352
rect 5413 5296 5760 5352
rect 5816 5296 5902 5352
rect 5958 5296 6300 5352
rect 6356 5296 6442 5352
rect 6498 5296 6845 5352
rect 6901 5296 6987 5352
rect 7043 5296 7382 5352
rect 7438 5296 7524 5352
rect 7580 5296 7919 5352
rect 7975 5296 8061 5352
rect 8117 5296 8462 5352
rect 8518 5296 8604 5352
rect 8660 5296 9004 5352
rect 9060 5296 9146 5352
rect 9202 5296 9547 5352
rect 9603 5296 9689 5352
rect 9745 5296 10081 5352
rect 10137 5296 10223 5352
rect 10279 5296 10622 5352
rect 10678 5296 10764 5352
rect 10820 5296 11162 5352
rect 11218 5296 11304 5352
rect 11360 5296 11702 5352
rect 11758 5296 11844 5352
rect 11900 5296 13200 5352
rect -400 5290 13200 5296
rect -400 5234 -286 5290
rect -230 5234 -162 5290
rect -106 5234 -38 5290
rect 18 5234 86 5290
rect 142 5234 210 5290
rect 266 5234 12526 5290
rect 12582 5234 12650 5290
rect 12706 5234 12774 5290
rect 12830 5234 12898 5290
rect 12954 5234 13022 5290
rect 13078 5234 13200 5290
rect -400 5210 13200 5234
rect -400 5166 903 5210
rect -400 5110 -286 5166
rect -230 5110 -162 5166
rect -106 5110 -38 5166
rect 18 5110 86 5166
rect 142 5110 210 5166
rect 266 5154 903 5166
rect 959 5154 1045 5210
rect 1101 5154 1444 5210
rect 1500 5154 1586 5210
rect 1642 5154 1984 5210
rect 2040 5154 2126 5210
rect 2182 5154 2521 5210
rect 2577 5154 2663 5210
rect 2719 5154 3058 5210
rect 3114 5154 3200 5210
rect 3256 5154 3602 5210
rect 3658 5154 3744 5210
rect 3800 5154 4138 5210
rect 4194 5154 4280 5210
rect 4336 5154 4678 5210
rect 4734 5154 4820 5210
rect 4876 5154 5215 5210
rect 5271 5154 5357 5210
rect 5413 5154 5760 5210
rect 5816 5154 5902 5210
rect 5958 5154 6300 5210
rect 6356 5154 6442 5210
rect 6498 5154 6845 5210
rect 6901 5154 6987 5210
rect 7043 5154 7382 5210
rect 7438 5154 7524 5210
rect 7580 5154 7919 5210
rect 7975 5154 8061 5210
rect 8117 5154 8462 5210
rect 8518 5154 8604 5210
rect 8660 5154 9004 5210
rect 9060 5154 9146 5210
rect 9202 5154 9547 5210
rect 9603 5154 9689 5210
rect 9745 5154 10081 5210
rect 10137 5154 10223 5210
rect 10279 5154 10622 5210
rect 10678 5154 10764 5210
rect 10820 5154 11162 5210
rect 11218 5154 11304 5210
rect 11360 5154 11702 5210
rect 11758 5154 11844 5210
rect 11900 5166 13200 5210
rect 11900 5154 12526 5166
rect 266 5110 12526 5154
rect 12582 5110 12650 5166
rect 12706 5110 12774 5166
rect 12830 5110 12898 5166
rect 12954 5110 13022 5166
rect 13078 5110 13200 5166
rect -400 5068 13200 5110
rect -400 5042 903 5068
rect -400 4986 -286 5042
rect -230 4986 -162 5042
rect -106 4986 -38 5042
rect 18 4986 86 5042
rect 142 4986 210 5042
rect 266 5012 903 5042
rect 959 5012 1045 5068
rect 1101 5012 1444 5068
rect 1500 5012 1586 5068
rect 1642 5012 1984 5068
rect 2040 5012 2126 5068
rect 2182 5012 2521 5068
rect 2577 5012 2663 5068
rect 2719 5012 3058 5068
rect 3114 5012 3200 5068
rect 3256 5012 3602 5068
rect 3658 5012 3744 5068
rect 3800 5012 4138 5068
rect 4194 5012 4280 5068
rect 4336 5012 4678 5068
rect 4734 5012 4820 5068
rect 4876 5012 5215 5068
rect 5271 5012 5357 5068
rect 5413 5012 5760 5068
rect 5816 5012 5902 5068
rect 5958 5012 6300 5068
rect 6356 5012 6442 5068
rect 6498 5012 6845 5068
rect 6901 5012 6987 5068
rect 7043 5012 7382 5068
rect 7438 5012 7524 5068
rect 7580 5012 7919 5068
rect 7975 5012 8061 5068
rect 8117 5012 8462 5068
rect 8518 5012 8604 5068
rect 8660 5012 9004 5068
rect 9060 5012 9146 5068
rect 9202 5012 9547 5068
rect 9603 5012 9689 5068
rect 9745 5012 10081 5068
rect 10137 5012 10223 5068
rect 10279 5012 10622 5068
rect 10678 5012 10764 5068
rect 10820 5012 11162 5068
rect 11218 5012 11304 5068
rect 11360 5012 11702 5068
rect 11758 5012 11844 5068
rect 11900 5042 13200 5068
rect 11900 5012 12526 5042
rect 266 4986 12526 5012
rect 12582 4986 12650 5042
rect 12706 4986 12774 5042
rect 12830 4986 12898 5042
rect 12954 4986 13022 5042
rect 13078 4986 13200 5042
rect -400 4926 13200 4986
rect -400 4918 903 4926
rect -400 4862 -286 4918
rect -230 4862 -162 4918
rect -106 4862 -38 4918
rect 18 4862 86 4918
rect 142 4862 210 4918
rect 266 4870 903 4918
rect 959 4870 1045 4926
rect 1101 4870 1444 4926
rect 1500 4870 1586 4926
rect 1642 4870 1984 4926
rect 2040 4870 2126 4926
rect 2182 4870 2521 4926
rect 2577 4870 2663 4926
rect 2719 4870 3058 4926
rect 3114 4870 3200 4926
rect 3256 4870 3602 4926
rect 3658 4870 3744 4926
rect 3800 4870 4138 4926
rect 4194 4870 4280 4926
rect 4336 4870 4678 4926
rect 4734 4870 4820 4926
rect 4876 4870 5215 4926
rect 5271 4870 5357 4926
rect 5413 4870 5760 4926
rect 5816 4870 5902 4926
rect 5958 4870 6300 4926
rect 6356 4870 6442 4926
rect 6498 4870 6845 4926
rect 6901 4870 6987 4926
rect 7043 4870 7382 4926
rect 7438 4870 7524 4926
rect 7580 4870 7919 4926
rect 7975 4870 8061 4926
rect 8117 4870 8462 4926
rect 8518 4870 8604 4926
rect 8660 4870 9004 4926
rect 9060 4870 9146 4926
rect 9202 4870 9547 4926
rect 9603 4870 9689 4926
rect 9745 4870 10081 4926
rect 10137 4870 10223 4926
rect 10279 4870 10622 4926
rect 10678 4870 10764 4926
rect 10820 4870 11162 4926
rect 11218 4870 11304 4926
rect 11360 4870 11702 4926
rect 11758 4870 11844 4926
rect 11900 4918 13200 4926
rect 11900 4870 12526 4918
rect 266 4862 12526 4870
rect 12582 4862 12650 4918
rect 12706 4862 12774 4918
rect 12830 4862 12898 4918
rect 12954 4862 13022 4918
rect 13078 4862 13200 4918
rect -400 4794 13200 4862
rect -400 4738 -286 4794
rect -230 4738 -162 4794
rect -106 4738 -38 4794
rect 18 4738 86 4794
rect 142 4738 210 4794
rect 266 4784 12526 4794
rect 266 4738 903 4784
rect -400 4728 903 4738
rect 959 4728 1045 4784
rect 1101 4728 1444 4784
rect 1500 4728 1586 4784
rect 1642 4728 1984 4784
rect 2040 4728 2126 4784
rect 2182 4728 2521 4784
rect 2577 4728 2663 4784
rect 2719 4728 3058 4784
rect 3114 4728 3200 4784
rect 3256 4728 3602 4784
rect 3658 4728 3744 4784
rect 3800 4728 4138 4784
rect 4194 4728 4280 4784
rect 4336 4728 4678 4784
rect 4734 4728 4820 4784
rect 4876 4728 5215 4784
rect 5271 4728 5357 4784
rect 5413 4728 5760 4784
rect 5816 4728 5902 4784
rect 5958 4728 6300 4784
rect 6356 4728 6442 4784
rect 6498 4728 6845 4784
rect 6901 4728 6987 4784
rect 7043 4728 7382 4784
rect 7438 4728 7524 4784
rect 7580 4728 7919 4784
rect 7975 4728 8061 4784
rect 8117 4728 8462 4784
rect 8518 4728 8604 4784
rect 8660 4728 9004 4784
rect 9060 4728 9146 4784
rect 9202 4728 9547 4784
rect 9603 4728 9689 4784
rect 9745 4728 10081 4784
rect 10137 4728 10223 4784
rect 10279 4728 10622 4784
rect 10678 4728 10764 4784
rect 10820 4728 11162 4784
rect 11218 4728 11304 4784
rect 11360 4728 11702 4784
rect 11758 4728 11844 4784
rect 11900 4738 12526 4784
rect 12582 4738 12650 4794
rect 12706 4738 12774 4794
rect 12830 4738 12898 4794
rect 12954 4738 13022 4794
rect 13078 4738 13200 4794
rect 11900 4728 13200 4738
rect -400 4670 13200 4728
rect -400 4614 -286 4670
rect -230 4614 -162 4670
rect -106 4614 -38 4670
rect 18 4614 86 4670
rect 142 4614 210 4670
rect 266 4642 12526 4670
rect 266 4614 903 4642
rect -400 4586 903 4614
rect 959 4586 1045 4642
rect 1101 4586 1444 4642
rect 1500 4586 1586 4642
rect 1642 4586 1984 4642
rect 2040 4586 2126 4642
rect 2182 4586 2521 4642
rect 2577 4586 2663 4642
rect 2719 4586 3058 4642
rect 3114 4586 3200 4642
rect 3256 4586 3602 4642
rect 3658 4586 3744 4642
rect 3800 4586 4138 4642
rect 4194 4586 4280 4642
rect 4336 4586 4678 4642
rect 4734 4586 4820 4642
rect 4876 4586 5215 4642
rect 5271 4586 5357 4642
rect 5413 4586 5760 4642
rect 5816 4586 5902 4642
rect 5958 4586 6300 4642
rect 6356 4586 6442 4642
rect 6498 4586 6845 4642
rect 6901 4586 6987 4642
rect 7043 4586 7382 4642
rect 7438 4586 7524 4642
rect 7580 4586 7919 4642
rect 7975 4586 8061 4642
rect 8117 4586 8462 4642
rect 8518 4586 8604 4642
rect 8660 4586 9004 4642
rect 9060 4586 9146 4642
rect 9202 4586 9547 4642
rect 9603 4586 9689 4642
rect 9745 4586 10081 4642
rect 10137 4586 10223 4642
rect 10279 4586 10622 4642
rect 10678 4586 10764 4642
rect 10820 4586 11162 4642
rect 11218 4586 11304 4642
rect 11360 4586 11702 4642
rect 11758 4586 11844 4642
rect 11900 4614 12526 4642
rect 12582 4614 12650 4670
rect 12706 4614 12774 4670
rect 12830 4614 12898 4670
rect 12954 4614 13022 4670
rect 13078 4614 13200 4670
rect 11900 4586 13200 4614
rect -400 4546 13200 4586
rect -400 4490 -286 4546
rect -230 4490 -162 4546
rect -106 4490 -38 4546
rect 18 4490 86 4546
rect 142 4490 210 4546
rect 266 4500 12526 4546
rect 266 4490 903 4500
rect -400 4444 903 4490
rect 959 4444 1045 4500
rect 1101 4444 1444 4500
rect 1500 4444 1586 4500
rect 1642 4444 1984 4500
rect 2040 4444 2126 4500
rect 2182 4444 2521 4500
rect 2577 4444 2663 4500
rect 2719 4444 3058 4500
rect 3114 4444 3200 4500
rect 3256 4444 3602 4500
rect 3658 4444 3744 4500
rect 3800 4444 4138 4500
rect 4194 4444 4280 4500
rect 4336 4444 4678 4500
rect 4734 4444 4820 4500
rect 4876 4444 5215 4500
rect 5271 4444 5357 4500
rect 5413 4444 5760 4500
rect 5816 4444 5902 4500
rect 5958 4444 6300 4500
rect 6356 4444 6442 4500
rect 6498 4444 6845 4500
rect 6901 4444 6987 4500
rect 7043 4444 7382 4500
rect 7438 4444 7524 4500
rect 7580 4444 7919 4500
rect 7975 4444 8061 4500
rect 8117 4444 8462 4500
rect 8518 4444 8604 4500
rect 8660 4444 9004 4500
rect 9060 4444 9146 4500
rect 9202 4444 9547 4500
rect 9603 4444 9689 4500
rect 9745 4444 10081 4500
rect 10137 4444 10223 4500
rect 10279 4444 10622 4500
rect 10678 4444 10764 4500
rect 10820 4444 11162 4500
rect 11218 4444 11304 4500
rect 11360 4444 11702 4500
rect 11758 4444 11844 4500
rect 11900 4490 12526 4500
rect 12582 4490 12650 4546
rect 12706 4490 12774 4546
rect 12830 4490 12898 4546
rect 12954 4490 13022 4546
rect 13078 4490 13200 4546
rect 11900 4444 13200 4490
rect -400 4422 13200 4444
rect -400 4366 -286 4422
rect -230 4366 -162 4422
rect -106 4366 -38 4422
rect 18 4366 86 4422
rect 142 4366 210 4422
rect 266 4366 12526 4422
rect 12582 4366 12650 4422
rect 12706 4366 12774 4422
rect 12830 4366 12898 4422
rect 12954 4366 13022 4422
rect 13078 4366 13200 4422
rect -400 4358 13200 4366
rect -400 4302 903 4358
rect 959 4302 1045 4358
rect 1101 4302 1444 4358
rect 1500 4302 1586 4358
rect 1642 4302 1984 4358
rect 2040 4302 2126 4358
rect 2182 4302 2521 4358
rect 2577 4302 2663 4358
rect 2719 4302 3058 4358
rect 3114 4302 3200 4358
rect 3256 4302 3602 4358
rect 3658 4302 3744 4358
rect 3800 4302 4138 4358
rect 4194 4302 4280 4358
rect 4336 4302 4678 4358
rect 4734 4302 4820 4358
rect 4876 4302 5215 4358
rect 5271 4302 5357 4358
rect 5413 4302 5760 4358
rect 5816 4302 5902 4358
rect 5958 4302 6300 4358
rect 6356 4302 6442 4358
rect 6498 4302 6845 4358
rect 6901 4302 6987 4358
rect 7043 4302 7382 4358
rect 7438 4302 7524 4358
rect 7580 4302 7919 4358
rect 7975 4302 8061 4358
rect 8117 4302 8462 4358
rect 8518 4302 8604 4358
rect 8660 4302 9004 4358
rect 9060 4302 9146 4358
rect 9202 4302 9547 4358
rect 9603 4302 9689 4358
rect 9745 4302 10081 4358
rect 10137 4302 10223 4358
rect 10279 4302 10622 4358
rect 10678 4302 10764 4358
rect 10820 4302 11162 4358
rect 11218 4302 11304 4358
rect 11360 4302 11702 4358
rect 11758 4302 11844 4358
rect 11900 4302 13200 4358
rect -400 4298 13200 4302
rect -400 4242 -286 4298
rect -230 4242 -162 4298
rect -106 4242 -38 4298
rect 18 4242 86 4298
rect 142 4242 210 4298
rect 266 4242 12526 4298
rect 12582 4242 12650 4298
rect 12706 4242 12774 4298
rect 12830 4242 12898 4298
rect 12954 4242 13022 4298
rect 13078 4242 13200 4298
rect -400 4216 13200 4242
rect -400 4174 903 4216
rect -400 4118 -286 4174
rect -230 4118 -162 4174
rect -106 4118 -38 4174
rect 18 4118 86 4174
rect 142 4118 210 4174
rect 266 4160 903 4174
rect 959 4160 1045 4216
rect 1101 4160 1444 4216
rect 1500 4160 1586 4216
rect 1642 4160 1984 4216
rect 2040 4160 2126 4216
rect 2182 4160 2521 4216
rect 2577 4160 2663 4216
rect 2719 4160 3058 4216
rect 3114 4160 3200 4216
rect 3256 4160 3602 4216
rect 3658 4160 3744 4216
rect 3800 4160 4138 4216
rect 4194 4160 4280 4216
rect 4336 4160 4678 4216
rect 4734 4160 4820 4216
rect 4876 4160 5215 4216
rect 5271 4160 5357 4216
rect 5413 4160 5760 4216
rect 5816 4160 5902 4216
rect 5958 4160 6300 4216
rect 6356 4160 6442 4216
rect 6498 4160 6845 4216
rect 6901 4160 6987 4216
rect 7043 4160 7382 4216
rect 7438 4160 7524 4216
rect 7580 4160 7919 4216
rect 7975 4160 8061 4216
rect 8117 4160 8462 4216
rect 8518 4160 8604 4216
rect 8660 4160 9004 4216
rect 9060 4160 9146 4216
rect 9202 4160 9547 4216
rect 9603 4160 9689 4216
rect 9745 4160 10081 4216
rect 10137 4160 10223 4216
rect 10279 4160 10622 4216
rect 10678 4160 10764 4216
rect 10820 4160 11162 4216
rect 11218 4160 11304 4216
rect 11360 4160 11702 4216
rect 11758 4160 11844 4216
rect 11900 4174 13200 4216
rect 11900 4160 12526 4174
rect 266 4118 12526 4160
rect 12582 4118 12650 4174
rect 12706 4118 12774 4174
rect 12830 4118 12898 4174
rect 12954 4118 13022 4174
rect 13078 4118 13200 4174
rect -400 4074 13200 4118
rect -400 4050 903 4074
rect -400 3994 -286 4050
rect -230 3994 -162 4050
rect -106 3994 -38 4050
rect 18 3994 86 4050
rect 142 3994 210 4050
rect 266 4018 903 4050
rect 959 4018 1045 4074
rect 1101 4018 1444 4074
rect 1500 4018 1586 4074
rect 1642 4018 1984 4074
rect 2040 4018 2126 4074
rect 2182 4018 2521 4074
rect 2577 4018 2663 4074
rect 2719 4018 3058 4074
rect 3114 4018 3200 4074
rect 3256 4018 3602 4074
rect 3658 4018 3744 4074
rect 3800 4018 4138 4074
rect 4194 4018 4280 4074
rect 4336 4018 4678 4074
rect 4734 4018 4820 4074
rect 4876 4018 5215 4074
rect 5271 4018 5357 4074
rect 5413 4018 5760 4074
rect 5816 4018 5902 4074
rect 5958 4018 6300 4074
rect 6356 4018 6442 4074
rect 6498 4018 6845 4074
rect 6901 4018 6987 4074
rect 7043 4018 7382 4074
rect 7438 4018 7524 4074
rect 7580 4018 7919 4074
rect 7975 4018 8061 4074
rect 8117 4018 8462 4074
rect 8518 4018 8604 4074
rect 8660 4018 9004 4074
rect 9060 4018 9146 4074
rect 9202 4018 9547 4074
rect 9603 4018 9689 4074
rect 9745 4018 10081 4074
rect 10137 4018 10223 4074
rect 10279 4018 10622 4074
rect 10678 4018 10764 4074
rect 10820 4018 11162 4074
rect 11218 4018 11304 4074
rect 11360 4018 11702 4074
rect 11758 4018 11844 4074
rect 11900 4050 13200 4074
rect 11900 4018 12526 4050
rect 266 3994 12526 4018
rect 12582 3994 12650 4050
rect 12706 3994 12774 4050
rect 12830 3994 12898 4050
rect 12954 3994 13022 4050
rect 13078 3994 13200 4050
rect -400 3932 13200 3994
rect -400 3926 903 3932
rect -400 3870 -286 3926
rect -230 3870 -162 3926
rect -106 3870 -38 3926
rect 18 3870 86 3926
rect 142 3870 210 3926
rect 266 3876 903 3926
rect 959 3876 1045 3932
rect 1101 3876 1444 3932
rect 1500 3876 1586 3932
rect 1642 3876 1984 3932
rect 2040 3876 2126 3932
rect 2182 3876 2521 3932
rect 2577 3876 2663 3932
rect 2719 3876 3058 3932
rect 3114 3876 3200 3932
rect 3256 3876 3602 3932
rect 3658 3876 3744 3932
rect 3800 3876 4138 3932
rect 4194 3876 4280 3932
rect 4336 3876 4678 3932
rect 4734 3876 4820 3932
rect 4876 3876 5215 3932
rect 5271 3876 5357 3932
rect 5413 3876 5760 3932
rect 5816 3876 5902 3932
rect 5958 3876 6300 3932
rect 6356 3876 6442 3932
rect 6498 3876 6845 3932
rect 6901 3876 6987 3932
rect 7043 3876 7382 3932
rect 7438 3876 7524 3932
rect 7580 3876 7919 3932
rect 7975 3876 8061 3932
rect 8117 3876 8462 3932
rect 8518 3876 8604 3932
rect 8660 3876 9004 3932
rect 9060 3876 9146 3932
rect 9202 3876 9547 3932
rect 9603 3876 9689 3932
rect 9745 3876 10081 3932
rect 10137 3876 10223 3932
rect 10279 3876 10622 3932
rect 10678 3876 10764 3932
rect 10820 3876 11162 3932
rect 11218 3876 11304 3932
rect 11360 3876 11702 3932
rect 11758 3876 11844 3932
rect 11900 3926 13200 3932
rect 11900 3876 12526 3926
rect 266 3870 12526 3876
rect 12582 3870 12650 3926
rect 12706 3870 12774 3926
rect 12830 3870 12898 3926
rect 12954 3870 13022 3926
rect 13078 3870 13200 3926
rect -400 3802 13200 3870
rect -400 3746 -286 3802
rect -230 3746 -162 3802
rect -106 3746 -38 3802
rect 18 3746 86 3802
rect 142 3746 210 3802
rect 266 3790 12526 3802
rect 266 3746 903 3790
rect -400 3734 903 3746
rect 959 3734 1045 3790
rect 1101 3734 1444 3790
rect 1500 3734 1586 3790
rect 1642 3734 1984 3790
rect 2040 3734 2126 3790
rect 2182 3734 2521 3790
rect 2577 3734 2663 3790
rect 2719 3734 3058 3790
rect 3114 3734 3200 3790
rect 3256 3734 3602 3790
rect 3658 3734 3744 3790
rect 3800 3734 4138 3790
rect 4194 3734 4280 3790
rect 4336 3734 4678 3790
rect 4734 3734 4820 3790
rect 4876 3734 5215 3790
rect 5271 3734 5357 3790
rect 5413 3734 5760 3790
rect 5816 3734 5902 3790
rect 5958 3734 6300 3790
rect 6356 3734 6442 3790
rect 6498 3734 6845 3790
rect 6901 3734 6987 3790
rect 7043 3734 7382 3790
rect 7438 3734 7524 3790
rect 7580 3734 7919 3790
rect 7975 3734 8061 3790
rect 8117 3734 8462 3790
rect 8518 3734 8604 3790
rect 8660 3734 9004 3790
rect 9060 3734 9146 3790
rect 9202 3734 9547 3790
rect 9603 3734 9689 3790
rect 9745 3734 10081 3790
rect 10137 3734 10223 3790
rect 10279 3734 10622 3790
rect 10678 3734 10764 3790
rect 10820 3734 11162 3790
rect 11218 3734 11304 3790
rect 11360 3734 11702 3790
rect 11758 3734 11844 3790
rect 11900 3746 12526 3790
rect 12582 3746 12650 3802
rect 12706 3746 12774 3802
rect 12830 3746 12898 3802
rect 12954 3746 13022 3802
rect 13078 3746 13200 3802
rect 11900 3734 13200 3746
rect -400 3678 13200 3734
rect -400 3622 -286 3678
rect -230 3622 -162 3678
rect -106 3622 -38 3678
rect 18 3622 86 3678
rect 142 3622 210 3678
rect 266 3648 12526 3678
rect 266 3622 903 3648
rect -400 3592 903 3622
rect 959 3592 1045 3648
rect 1101 3592 1444 3648
rect 1500 3592 1586 3648
rect 1642 3592 1984 3648
rect 2040 3592 2126 3648
rect 2182 3592 2521 3648
rect 2577 3592 2663 3648
rect 2719 3592 3058 3648
rect 3114 3592 3200 3648
rect 3256 3592 3602 3648
rect 3658 3592 3744 3648
rect 3800 3592 4138 3648
rect 4194 3592 4280 3648
rect 4336 3592 4678 3648
rect 4734 3592 4820 3648
rect 4876 3592 5215 3648
rect 5271 3592 5357 3648
rect 5413 3592 5760 3648
rect 5816 3592 5902 3648
rect 5958 3592 6300 3648
rect 6356 3592 6442 3648
rect 6498 3592 6845 3648
rect 6901 3592 6987 3648
rect 7043 3592 7382 3648
rect 7438 3592 7524 3648
rect 7580 3592 7919 3648
rect 7975 3592 8061 3648
rect 8117 3592 8462 3648
rect 8518 3592 8604 3648
rect 8660 3592 9004 3648
rect 9060 3592 9146 3648
rect 9202 3592 9547 3648
rect 9603 3592 9689 3648
rect 9745 3592 10081 3648
rect 10137 3592 10223 3648
rect 10279 3592 10622 3648
rect 10678 3592 10764 3648
rect 10820 3592 11162 3648
rect 11218 3592 11304 3648
rect 11360 3592 11702 3648
rect 11758 3592 11844 3648
rect 11900 3622 12526 3648
rect 12582 3622 12650 3678
rect 12706 3622 12774 3678
rect 12830 3622 12898 3678
rect 12954 3622 13022 3678
rect 13078 3622 13200 3678
rect 11900 3592 13200 3622
rect -400 3554 13200 3592
rect -400 3498 -286 3554
rect -230 3498 -162 3554
rect -106 3498 -38 3554
rect 18 3498 86 3554
rect 142 3498 210 3554
rect 266 3506 12526 3554
rect 266 3498 903 3506
rect -400 3450 903 3498
rect 959 3450 1045 3506
rect 1101 3450 1444 3506
rect 1500 3450 1586 3506
rect 1642 3450 1984 3506
rect 2040 3450 2126 3506
rect 2182 3450 2521 3506
rect 2577 3450 2663 3506
rect 2719 3450 3058 3506
rect 3114 3450 3200 3506
rect 3256 3450 3602 3506
rect 3658 3450 3744 3506
rect 3800 3450 4138 3506
rect 4194 3450 4280 3506
rect 4336 3450 4678 3506
rect 4734 3450 4820 3506
rect 4876 3450 5215 3506
rect 5271 3450 5357 3506
rect 5413 3450 5760 3506
rect 5816 3450 5902 3506
rect 5958 3450 6300 3506
rect 6356 3450 6442 3506
rect 6498 3450 6845 3506
rect 6901 3450 6987 3506
rect 7043 3450 7382 3506
rect 7438 3450 7524 3506
rect 7580 3450 7919 3506
rect 7975 3450 8061 3506
rect 8117 3450 8462 3506
rect 8518 3450 8604 3506
rect 8660 3450 9004 3506
rect 9060 3450 9146 3506
rect 9202 3450 9547 3506
rect 9603 3450 9689 3506
rect 9745 3450 10081 3506
rect 10137 3450 10223 3506
rect 10279 3450 10622 3506
rect 10678 3450 10764 3506
rect 10820 3450 11162 3506
rect 11218 3450 11304 3506
rect 11360 3450 11702 3506
rect 11758 3450 11844 3506
rect 11900 3498 12526 3506
rect 12582 3498 12650 3554
rect 12706 3498 12774 3554
rect 12830 3498 12898 3554
rect 12954 3498 13022 3554
rect 13078 3498 13200 3554
rect 11900 3450 13200 3498
rect -400 3430 13200 3450
rect -400 3374 -286 3430
rect -230 3374 -162 3430
rect -106 3374 -38 3430
rect 18 3374 86 3430
rect 142 3374 210 3430
rect 266 3374 12526 3430
rect 12582 3374 12650 3430
rect 12706 3374 12774 3430
rect 12830 3374 12898 3430
rect 12954 3374 13022 3430
rect 13078 3374 13200 3430
rect -400 3364 13200 3374
rect -400 3308 903 3364
rect 959 3308 1045 3364
rect 1101 3308 1444 3364
rect 1500 3308 1586 3364
rect 1642 3308 1984 3364
rect 2040 3308 2126 3364
rect 2182 3308 2521 3364
rect 2577 3308 2663 3364
rect 2719 3308 3058 3364
rect 3114 3308 3200 3364
rect 3256 3308 3602 3364
rect 3658 3308 3744 3364
rect 3800 3308 4138 3364
rect 4194 3308 4280 3364
rect 4336 3308 4678 3364
rect 4734 3308 4820 3364
rect 4876 3308 5215 3364
rect 5271 3308 5357 3364
rect 5413 3308 5760 3364
rect 5816 3308 5902 3364
rect 5958 3308 6300 3364
rect 6356 3308 6442 3364
rect 6498 3308 6845 3364
rect 6901 3308 6987 3364
rect 7043 3308 7382 3364
rect 7438 3308 7524 3364
rect 7580 3308 7919 3364
rect 7975 3308 8061 3364
rect 8117 3308 8462 3364
rect 8518 3308 8604 3364
rect 8660 3308 9004 3364
rect 9060 3308 9146 3364
rect 9202 3308 9547 3364
rect 9603 3308 9689 3364
rect 9745 3308 10081 3364
rect 10137 3308 10223 3364
rect 10279 3308 10622 3364
rect 10678 3308 10764 3364
rect 10820 3308 11162 3364
rect 11218 3308 11304 3364
rect 11360 3308 11702 3364
rect 11758 3308 11844 3364
rect 11900 3308 13200 3364
rect -400 3306 13200 3308
rect -400 3250 -286 3306
rect -230 3250 -162 3306
rect -106 3250 -38 3306
rect 18 3250 86 3306
rect 142 3250 210 3306
rect 266 3250 12526 3306
rect 12582 3250 12650 3306
rect 12706 3250 12774 3306
rect 12830 3250 12898 3306
rect 12954 3250 13022 3306
rect 13078 3250 13200 3306
rect -400 3222 13200 3250
rect -400 3182 903 3222
rect -400 3126 -286 3182
rect -230 3126 -162 3182
rect -106 3126 -38 3182
rect 18 3126 86 3182
rect 142 3126 210 3182
rect 266 3166 903 3182
rect 959 3166 1045 3222
rect 1101 3166 1444 3222
rect 1500 3166 1586 3222
rect 1642 3166 1984 3222
rect 2040 3166 2126 3222
rect 2182 3166 2521 3222
rect 2577 3166 2663 3222
rect 2719 3166 3058 3222
rect 3114 3166 3200 3222
rect 3256 3166 3602 3222
rect 3658 3166 3744 3222
rect 3800 3166 4138 3222
rect 4194 3166 4280 3222
rect 4336 3166 4678 3222
rect 4734 3166 4820 3222
rect 4876 3166 5215 3222
rect 5271 3166 5357 3222
rect 5413 3166 5760 3222
rect 5816 3166 5902 3222
rect 5958 3166 6300 3222
rect 6356 3166 6442 3222
rect 6498 3166 6845 3222
rect 6901 3166 6987 3222
rect 7043 3166 7382 3222
rect 7438 3166 7524 3222
rect 7580 3166 7919 3222
rect 7975 3166 8061 3222
rect 8117 3166 8462 3222
rect 8518 3166 8604 3222
rect 8660 3166 9004 3222
rect 9060 3166 9146 3222
rect 9202 3166 9547 3222
rect 9603 3166 9689 3222
rect 9745 3166 10081 3222
rect 10137 3166 10223 3222
rect 10279 3166 10622 3222
rect 10678 3166 10764 3222
rect 10820 3166 11162 3222
rect 11218 3166 11304 3222
rect 11360 3166 11702 3222
rect 11758 3166 11844 3222
rect 11900 3182 13200 3222
rect 11900 3166 12526 3182
rect 266 3126 12526 3166
rect 12582 3126 12650 3182
rect 12706 3126 12774 3182
rect 12830 3126 12898 3182
rect 12954 3126 13022 3182
rect 13078 3126 13200 3182
rect -400 3080 13200 3126
rect -400 3058 903 3080
rect -400 3002 -286 3058
rect -230 3002 -162 3058
rect -106 3002 -38 3058
rect 18 3002 86 3058
rect 142 3002 210 3058
rect 266 3024 903 3058
rect 959 3024 1045 3080
rect 1101 3024 1444 3080
rect 1500 3024 1586 3080
rect 1642 3024 1984 3080
rect 2040 3024 2126 3080
rect 2182 3024 2521 3080
rect 2577 3024 2663 3080
rect 2719 3024 3058 3080
rect 3114 3024 3200 3080
rect 3256 3024 3602 3080
rect 3658 3024 3744 3080
rect 3800 3024 4138 3080
rect 4194 3024 4280 3080
rect 4336 3024 4678 3080
rect 4734 3024 4820 3080
rect 4876 3024 5215 3080
rect 5271 3024 5357 3080
rect 5413 3024 5760 3080
rect 5816 3024 5902 3080
rect 5958 3024 6300 3080
rect 6356 3024 6442 3080
rect 6498 3024 6845 3080
rect 6901 3024 6987 3080
rect 7043 3024 7382 3080
rect 7438 3024 7524 3080
rect 7580 3024 7919 3080
rect 7975 3024 8061 3080
rect 8117 3024 8462 3080
rect 8518 3024 8604 3080
rect 8660 3024 9004 3080
rect 9060 3024 9146 3080
rect 9202 3024 9547 3080
rect 9603 3024 9689 3080
rect 9745 3024 10081 3080
rect 10137 3024 10223 3080
rect 10279 3024 10622 3080
rect 10678 3024 10764 3080
rect 10820 3024 11162 3080
rect 11218 3024 11304 3080
rect 11360 3024 11702 3080
rect 11758 3024 11844 3080
rect 11900 3058 13200 3080
rect 11900 3024 12526 3058
rect 266 3002 12526 3024
rect 12582 3002 12650 3058
rect 12706 3002 12774 3058
rect 12830 3002 12898 3058
rect 12954 3002 13022 3058
rect 13078 3002 13200 3058
rect -400 2938 13200 3002
rect -400 2934 903 2938
rect -400 2878 -286 2934
rect -230 2878 -162 2934
rect -106 2878 -38 2934
rect 18 2878 86 2934
rect 142 2878 210 2934
rect 266 2882 903 2934
rect 959 2882 1045 2938
rect 1101 2882 1444 2938
rect 1500 2882 1586 2938
rect 1642 2882 1984 2938
rect 2040 2882 2126 2938
rect 2182 2882 2521 2938
rect 2577 2882 2663 2938
rect 2719 2882 3058 2938
rect 3114 2882 3200 2938
rect 3256 2882 3602 2938
rect 3658 2882 3744 2938
rect 3800 2882 4138 2938
rect 4194 2882 4280 2938
rect 4336 2882 4678 2938
rect 4734 2882 4820 2938
rect 4876 2882 5215 2938
rect 5271 2882 5357 2938
rect 5413 2882 5760 2938
rect 5816 2882 5902 2938
rect 5958 2882 6300 2938
rect 6356 2882 6442 2938
rect 6498 2882 6845 2938
rect 6901 2882 6987 2938
rect 7043 2882 7382 2938
rect 7438 2882 7524 2938
rect 7580 2882 7919 2938
rect 7975 2882 8061 2938
rect 8117 2882 8462 2938
rect 8518 2882 8604 2938
rect 8660 2882 9004 2938
rect 9060 2882 9146 2938
rect 9202 2882 9547 2938
rect 9603 2882 9689 2938
rect 9745 2882 10081 2938
rect 10137 2882 10223 2938
rect 10279 2882 10622 2938
rect 10678 2882 10764 2938
rect 10820 2882 11162 2938
rect 11218 2882 11304 2938
rect 11360 2882 11702 2938
rect 11758 2882 11844 2938
rect 11900 2934 13200 2938
rect 11900 2882 12526 2934
rect 266 2878 12526 2882
rect 12582 2878 12650 2934
rect 12706 2878 12774 2934
rect 12830 2878 12898 2934
rect 12954 2878 13022 2934
rect 13078 2878 13200 2934
rect -400 2810 13200 2878
rect -400 2754 -286 2810
rect -230 2754 -162 2810
rect -106 2754 -38 2810
rect 18 2754 86 2810
rect 142 2754 210 2810
rect 266 2796 12526 2810
rect 266 2754 903 2796
rect -400 2740 903 2754
rect 959 2740 1045 2796
rect 1101 2740 1444 2796
rect 1500 2740 1586 2796
rect 1642 2740 1984 2796
rect 2040 2740 2126 2796
rect 2182 2740 2521 2796
rect 2577 2740 2663 2796
rect 2719 2740 3058 2796
rect 3114 2740 3200 2796
rect 3256 2740 3602 2796
rect 3658 2740 3744 2796
rect 3800 2740 4138 2796
rect 4194 2740 4280 2796
rect 4336 2740 4678 2796
rect 4734 2740 4820 2796
rect 4876 2740 5215 2796
rect 5271 2740 5357 2796
rect 5413 2740 5760 2796
rect 5816 2740 5902 2796
rect 5958 2740 6300 2796
rect 6356 2740 6442 2796
rect 6498 2740 6845 2796
rect 6901 2740 6987 2796
rect 7043 2740 7382 2796
rect 7438 2740 7524 2796
rect 7580 2740 7919 2796
rect 7975 2740 8061 2796
rect 8117 2740 8462 2796
rect 8518 2740 8604 2796
rect 8660 2740 9004 2796
rect 9060 2740 9146 2796
rect 9202 2740 9547 2796
rect 9603 2740 9689 2796
rect 9745 2740 10081 2796
rect 10137 2740 10223 2796
rect 10279 2740 10622 2796
rect 10678 2740 10764 2796
rect 10820 2740 11162 2796
rect 11218 2740 11304 2796
rect 11360 2740 11702 2796
rect 11758 2740 11844 2796
rect 11900 2754 12526 2796
rect 12582 2754 12650 2810
rect 12706 2754 12774 2810
rect 12830 2754 12898 2810
rect 12954 2754 13022 2810
rect 13078 2754 13200 2810
rect 11900 2740 13200 2754
rect -400 2686 13200 2740
rect -400 2630 -286 2686
rect -230 2630 -162 2686
rect -106 2630 -38 2686
rect 18 2630 86 2686
rect 142 2630 210 2686
rect 266 2654 12526 2686
rect 266 2630 903 2654
rect -400 2598 903 2630
rect 959 2598 1045 2654
rect 1101 2598 1444 2654
rect 1500 2598 1586 2654
rect 1642 2598 1984 2654
rect 2040 2598 2126 2654
rect 2182 2598 2521 2654
rect 2577 2598 2663 2654
rect 2719 2598 3058 2654
rect 3114 2598 3200 2654
rect 3256 2598 3602 2654
rect 3658 2598 3744 2654
rect 3800 2598 4138 2654
rect 4194 2598 4280 2654
rect 4336 2598 4678 2654
rect 4734 2598 4820 2654
rect 4876 2598 5215 2654
rect 5271 2598 5357 2654
rect 5413 2598 5760 2654
rect 5816 2598 5902 2654
rect 5958 2598 6300 2654
rect 6356 2598 6442 2654
rect 6498 2598 6845 2654
rect 6901 2598 6987 2654
rect 7043 2598 7382 2654
rect 7438 2598 7524 2654
rect 7580 2598 7919 2654
rect 7975 2598 8061 2654
rect 8117 2598 8462 2654
rect 8518 2598 8604 2654
rect 8660 2598 9004 2654
rect 9060 2598 9146 2654
rect 9202 2598 9547 2654
rect 9603 2598 9689 2654
rect 9745 2598 10081 2654
rect 10137 2598 10223 2654
rect 10279 2598 10622 2654
rect 10678 2598 10764 2654
rect 10820 2598 11162 2654
rect 11218 2598 11304 2654
rect 11360 2598 11702 2654
rect 11758 2598 11844 2654
rect 11900 2630 12526 2654
rect 12582 2630 12650 2686
rect 12706 2630 12774 2686
rect 12830 2630 12898 2686
rect 12954 2630 13022 2686
rect 13078 2630 13200 2686
rect 11900 2598 13200 2630
rect -400 2562 13200 2598
rect -400 2506 -286 2562
rect -230 2506 -162 2562
rect -106 2506 -38 2562
rect 18 2506 86 2562
rect 142 2506 210 2562
rect 266 2512 12526 2562
rect 266 2506 903 2512
rect -400 2456 903 2506
rect 959 2456 1045 2512
rect 1101 2456 1444 2512
rect 1500 2456 1586 2512
rect 1642 2456 1984 2512
rect 2040 2456 2126 2512
rect 2182 2456 2521 2512
rect 2577 2456 2663 2512
rect 2719 2456 3058 2512
rect 3114 2456 3200 2512
rect 3256 2456 3602 2512
rect 3658 2456 3744 2512
rect 3800 2456 4138 2512
rect 4194 2456 4280 2512
rect 4336 2456 4678 2512
rect 4734 2456 4820 2512
rect 4876 2456 5215 2512
rect 5271 2456 5357 2512
rect 5413 2456 5760 2512
rect 5816 2456 5902 2512
rect 5958 2456 6300 2512
rect 6356 2456 6442 2512
rect 6498 2456 6845 2512
rect 6901 2456 6987 2512
rect 7043 2456 7382 2512
rect 7438 2456 7524 2512
rect 7580 2456 7919 2512
rect 7975 2456 8061 2512
rect 8117 2456 8462 2512
rect 8518 2456 8604 2512
rect 8660 2456 9004 2512
rect 9060 2456 9146 2512
rect 9202 2456 9547 2512
rect 9603 2456 9689 2512
rect 9745 2456 10081 2512
rect 10137 2456 10223 2512
rect 10279 2456 10622 2512
rect 10678 2456 10764 2512
rect 10820 2456 11162 2512
rect 11218 2456 11304 2512
rect 11360 2456 11702 2512
rect 11758 2456 11844 2512
rect 11900 2506 12526 2512
rect 12582 2506 12650 2562
rect 12706 2506 12774 2562
rect 12830 2506 12898 2562
rect 12954 2506 13022 2562
rect 13078 2506 13200 2562
rect 11900 2456 13200 2506
rect -400 2438 13200 2456
rect -400 2382 -286 2438
rect -230 2382 -162 2438
rect -106 2382 -38 2438
rect 18 2382 86 2438
rect 142 2382 210 2438
rect 266 2382 12526 2438
rect 12582 2382 12650 2438
rect 12706 2382 12774 2438
rect 12830 2382 12898 2438
rect 12954 2382 13022 2438
rect 13078 2382 13200 2438
rect -400 2370 13200 2382
rect -400 2314 903 2370
rect 959 2314 1045 2370
rect 1101 2314 1444 2370
rect 1500 2314 1586 2370
rect 1642 2314 1984 2370
rect 2040 2314 2126 2370
rect 2182 2314 2521 2370
rect 2577 2314 2663 2370
rect 2719 2314 3058 2370
rect 3114 2314 3200 2370
rect 3256 2314 3602 2370
rect 3658 2314 3744 2370
rect 3800 2314 4138 2370
rect 4194 2314 4280 2370
rect 4336 2314 4678 2370
rect 4734 2314 4820 2370
rect 4876 2314 5215 2370
rect 5271 2314 5357 2370
rect 5413 2314 5760 2370
rect 5816 2314 5902 2370
rect 5958 2314 6300 2370
rect 6356 2314 6442 2370
rect 6498 2314 6845 2370
rect 6901 2314 6987 2370
rect 7043 2314 7382 2370
rect 7438 2314 7524 2370
rect 7580 2314 7919 2370
rect 7975 2314 8061 2370
rect 8117 2314 8462 2370
rect 8518 2314 8604 2370
rect 8660 2314 9004 2370
rect 9060 2314 9146 2370
rect 9202 2314 9547 2370
rect 9603 2314 9689 2370
rect 9745 2314 10081 2370
rect 10137 2314 10223 2370
rect 10279 2314 10622 2370
rect 10678 2314 10764 2370
rect 10820 2314 11162 2370
rect 11218 2314 11304 2370
rect 11360 2314 11702 2370
rect 11758 2314 11844 2370
rect 11900 2314 13200 2370
rect -400 2258 -286 2314
rect -230 2258 -162 2314
rect -106 2258 -38 2314
rect 18 2258 86 2314
rect 142 2258 210 2314
rect 266 2258 12526 2314
rect 12582 2258 12650 2314
rect 12706 2258 12774 2314
rect 12830 2258 12898 2314
rect 12954 2258 13022 2314
rect 13078 2258 13200 2314
rect -400 2228 13200 2258
rect -400 2190 903 2228
rect -400 2134 -286 2190
rect -230 2134 -162 2190
rect -106 2134 -38 2190
rect 18 2134 86 2190
rect 142 2134 210 2190
rect 266 2172 903 2190
rect 959 2172 1045 2228
rect 1101 2172 1444 2228
rect 1500 2172 1586 2228
rect 1642 2172 1984 2228
rect 2040 2172 2126 2228
rect 2182 2172 2521 2228
rect 2577 2172 2663 2228
rect 2719 2172 3058 2228
rect 3114 2172 3200 2228
rect 3256 2172 3602 2228
rect 3658 2172 3744 2228
rect 3800 2172 4138 2228
rect 4194 2172 4280 2228
rect 4336 2172 4678 2228
rect 4734 2172 4820 2228
rect 4876 2172 5215 2228
rect 5271 2172 5357 2228
rect 5413 2172 5760 2228
rect 5816 2172 5902 2228
rect 5958 2172 6300 2228
rect 6356 2172 6442 2228
rect 6498 2172 6845 2228
rect 6901 2172 6987 2228
rect 7043 2172 7382 2228
rect 7438 2172 7524 2228
rect 7580 2172 7919 2228
rect 7975 2172 8061 2228
rect 8117 2172 8462 2228
rect 8518 2172 8604 2228
rect 8660 2172 9004 2228
rect 9060 2172 9146 2228
rect 9202 2172 9547 2228
rect 9603 2172 9689 2228
rect 9745 2172 10081 2228
rect 10137 2172 10223 2228
rect 10279 2172 10622 2228
rect 10678 2172 10764 2228
rect 10820 2172 11162 2228
rect 11218 2172 11304 2228
rect 11360 2172 11702 2228
rect 11758 2172 11844 2228
rect 11900 2190 13200 2228
rect 11900 2172 12526 2190
rect 266 2134 12526 2172
rect 12582 2134 12650 2190
rect 12706 2134 12774 2190
rect 12830 2134 12898 2190
rect 12954 2134 13022 2190
rect 13078 2134 13200 2190
rect -400 2086 13200 2134
rect -400 2066 903 2086
rect -400 2010 -286 2066
rect -230 2010 -162 2066
rect -106 2010 -38 2066
rect 18 2010 86 2066
rect 142 2010 210 2066
rect 266 2030 903 2066
rect 959 2030 1045 2086
rect 1101 2030 1444 2086
rect 1500 2030 1586 2086
rect 1642 2030 1984 2086
rect 2040 2030 2126 2086
rect 2182 2030 2521 2086
rect 2577 2030 2663 2086
rect 2719 2030 3058 2086
rect 3114 2030 3200 2086
rect 3256 2030 3602 2086
rect 3658 2030 3744 2086
rect 3800 2030 4138 2086
rect 4194 2030 4280 2086
rect 4336 2030 4678 2086
rect 4734 2030 4820 2086
rect 4876 2030 5215 2086
rect 5271 2030 5357 2086
rect 5413 2030 5760 2086
rect 5816 2030 5902 2086
rect 5958 2030 6300 2086
rect 6356 2030 6442 2086
rect 6498 2030 6845 2086
rect 6901 2030 6987 2086
rect 7043 2030 7382 2086
rect 7438 2030 7524 2086
rect 7580 2030 7919 2086
rect 7975 2030 8061 2086
rect 8117 2030 8462 2086
rect 8518 2030 8604 2086
rect 8660 2030 9004 2086
rect 9060 2030 9146 2086
rect 9202 2030 9547 2086
rect 9603 2030 9689 2086
rect 9745 2030 10081 2086
rect 10137 2030 10223 2086
rect 10279 2030 10622 2086
rect 10678 2030 10764 2086
rect 10820 2030 11162 2086
rect 11218 2030 11304 2086
rect 11360 2030 11702 2086
rect 11758 2030 11844 2086
rect 11900 2066 13200 2086
rect 11900 2030 12526 2066
rect 266 2010 12526 2030
rect 12582 2010 12650 2066
rect 12706 2010 12774 2066
rect 12830 2010 12898 2066
rect 12954 2010 13022 2066
rect 13078 2010 13200 2066
rect -400 1944 13200 2010
rect -400 1942 903 1944
rect -400 1886 -286 1942
rect -230 1886 -162 1942
rect -106 1886 -38 1942
rect 18 1886 86 1942
rect 142 1886 210 1942
rect 266 1888 903 1942
rect 959 1888 1045 1944
rect 1101 1888 1444 1944
rect 1500 1888 1586 1944
rect 1642 1888 1984 1944
rect 2040 1888 2126 1944
rect 2182 1888 2521 1944
rect 2577 1888 2663 1944
rect 2719 1888 3058 1944
rect 3114 1888 3200 1944
rect 3256 1888 3602 1944
rect 3658 1888 3744 1944
rect 3800 1888 4138 1944
rect 4194 1888 4280 1944
rect 4336 1888 4678 1944
rect 4734 1888 4820 1944
rect 4876 1888 5215 1944
rect 5271 1888 5357 1944
rect 5413 1888 5760 1944
rect 5816 1888 5902 1944
rect 5958 1888 6300 1944
rect 6356 1888 6442 1944
rect 6498 1888 6845 1944
rect 6901 1888 6987 1944
rect 7043 1888 7382 1944
rect 7438 1888 7524 1944
rect 7580 1888 7919 1944
rect 7975 1888 8061 1944
rect 8117 1888 8462 1944
rect 8518 1888 8604 1944
rect 8660 1888 9004 1944
rect 9060 1888 9146 1944
rect 9202 1888 9547 1944
rect 9603 1888 9689 1944
rect 9745 1888 10081 1944
rect 10137 1888 10223 1944
rect 10279 1888 10622 1944
rect 10678 1888 10764 1944
rect 10820 1888 11162 1944
rect 11218 1888 11304 1944
rect 11360 1888 11702 1944
rect 11758 1888 11844 1944
rect 11900 1942 13200 1944
rect 11900 1888 12526 1942
rect 266 1886 12526 1888
rect 12582 1886 12650 1942
rect 12706 1886 12774 1942
rect 12830 1886 12898 1942
rect 12954 1886 13022 1942
rect 13078 1886 13200 1942
rect -400 1818 13200 1886
rect -400 1762 -286 1818
rect -230 1762 -162 1818
rect -106 1762 -38 1818
rect 18 1762 86 1818
rect 142 1762 210 1818
rect 266 1802 12526 1818
rect 266 1762 903 1802
rect -400 1746 903 1762
rect 959 1746 1045 1802
rect 1101 1746 1444 1802
rect 1500 1746 1586 1802
rect 1642 1746 1984 1802
rect 2040 1746 2126 1802
rect 2182 1746 2521 1802
rect 2577 1746 2663 1802
rect 2719 1746 3058 1802
rect 3114 1746 3200 1802
rect 3256 1746 3602 1802
rect 3658 1746 3744 1802
rect 3800 1746 4138 1802
rect 4194 1746 4280 1802
rect 4336 1746 4678 1802
rect 4734 1746 4820 1802
rect 4876 1746 5215 1802
rect 5271 1746 5357 1802
rect 5413 1746 5760 1802
rect 5816 1746 5902 1802
rect 5958 1746 6300 1802
rect 6356 1746 6442 1802
rect 6498 1746 6845 1802
rect 6901 1746 6987 1802
rect 7043 1746 7382 1802
rect 7438 1746 7524 1802
rect 7580 1746 7919 1802
rect 7975 1746 8061 1802
rect 8117 1746 8462 1802
rect 8518 1746 8604 1802
rect 8660 1746 9004 1802
rect 9060 1746 9146 1802
rect 9202 1746 9547 1802
rect 9603 1746 9689 1802
rect 9745 1746 10081 1802
rect 10137 1746 10223 1802
rect 10279 1746 10622 1802
rect 10678 1746 10764 1802
rect 10820 1746 11162 1802
rect 11218 1746 11304 1802
rect 11360 1746 11702 1802
rect 11758 1746 11844 1802
rect 11900 1762 12526 1802
rect 12582 1762 12650 1818
rect 12706 1762 12774 1818
rect 12830 1762 12898 1818
rect 12954 1762 13022 1818
rect 13078 1762 13200 1818
rect 11900 1746 13200 1762
rect -400 1694 13200 1746
rect -400 1638 -286 1694
rect -230 1638 -162 1694
rect -106 1638 -38 1694
rect 18 1638 86 1694
rect 142 1638 210 1694
rect 266 1660 12526 1694
rect 266 1638 903 1660
rect -400 1604 903 1638
rect 959 1604 1045 1660
rect 1101 1604 1444 1660
rect 1500 1604 1586 1660
rect 1642 1604 1984 1660
rect 2040 1604 2126 1660
rect 2182 1604 2521 1660
rect 2577 1604 2663 1660
rect 2719 1604 3058 1660
rect 3114 1604 3200 1660
rect 3256 1604 3602 1660
rect 3658 1604 3744 1660
rect 3800 1604 4138 1660
rect 4194 1604 4280 1660
rect 4336 1604 4678 1660
rect 4734 1604 4820 1660
rect 4876 1604 5215 1660
rect 5271 1604 5357 1660
rect 5413 1604 5760 1660
rect 5816 1604 5902 1660
rect 5958 1604 6300 1660
rect 6356 1604 6442 1660
rect 6498 1604 6845 1660
rect 6901 1604 6987 1660
rect 7043 1604 7382 1660
rect 7438 1604 7524 1660
rect 7580 1604 7919 1660
rect 7975 1604 8061 1660
rect 8117 1604 8462 1660
rect 8518 1604 8604 1660
rect 8660 1604 9004 1660
rect 9060 1604 9146 1660
rect 9202 1604 9547 1660
rect 9603 1604 9689 1660
rect 9745 1604 10081 1660
rect 10137 1604 10223 1660
rect 10279 1604 10622 1660
rect 10678 1604 10764 1660
rect 10820 1604 11162 1660
rect 11218 1604 11304 1660
rect 11360 1604 11702 1660
rect 11758 1604 11844 1660
rect 11900 1638 12526 1660
rect 12582 1638 12650 1694
rect 12706 1638 12774 1694
rect 12830 1638 12898 1694
rect 12954 1638 13022 1694
rect 13078 1638 13200 1694
rect 11900 1604 13200 1638
rect -400 1570 13200 1604
rect -400 1514 -286 1570
rect -230 1514 -162 1570
rect -106 1514 -38 1570
rect 18 1514 86 1570
rect 142 1514 210 1570
rect 266 1518 12526 1570
rect 266 1514 903 1518
rect -400 1462 903 1514
rect 959 1462 1045 1518
rect 1101 1462 1444 1518
rect 1500 1462 1586 1518
rect 1642 1462 1984 1518
rect 2040 1462 2126 1518
rect 2182 1462 2521 1518
rect 2577 1462 2663 1518
rect 2719 1462 3058 1518
rect 3114 1462 3200 1518
rect 3256 1462 3602 1518
rect 3658 1462 3744 1518
rect 3800 1462 4138 1518
rect 4194 1462 4280 1518
rect 4336 1462 4678 1518
rect 4734 1462 4820 1518
rect 4876 1462 5215 1518
rect 5271 1462 5357 1518
rect 5413 1462 5760 1518
rect 5816 1462 5902 1518
rect 5958 1462 6300 1518
rect 6356 1462 6442 1518
rect 6498 1462 6845 1518
rect 6901 1462 6987 1518
rect 7043 1462 7382 1518
rect 7438 1462 7524 1518
rect 7580 1462 7919 1518
rect 7975 1462 8061 1518
rect 8117 1462 8462 1518
rect 8518 1462 8604 1518
rect 8660 1462 9004 1518
rect 9060 1462 9146 1518
rect 9202 1462 9547 1518
rect 9603 1462 9689 1518
rect 9745 1462 10081 1518
rect 10137 1462 10223 1518
rect 10279 1462 10622 1518
rect 10678 1462 10764 1518
rect 10820 1462 11162 1518
rect 11218 1462 11304 1518
rect 11360 1462 11702 1518
rect 11758 1462 11844 1518
rect 11900 1514 12526 1518
rect 12582 1514 12650 1570
rect 12706 1514 12774 1570
rect 12830 1514 12898 1570
rect 12954 1514 13022 1570
rect 13078 1514 13200 1570
rect 11900 1462 13200 1514
rect -400 1446 13200 1462
rect -400 1390 -286 1446
rect -230 1390 -162 1446
rect -106 1390 -38 1446
rect 18 1390 86 1446
rect 142 1390 210 1446
rect 266 1390 12526 1446
rect 12582 1390 12650 1446
rect 12706 1390 12774 1446
rect 12830 1390 12898 1446
rect 12954 1390 13022 1446
rect 13078 1390 13200 1446
rect -400 1376 13200 1390
rect -400 1322 903 1376
rect -400 1266 -286 1322
rect -230 1266 -162 1322
rect -106 1266 -38 1322
rect 18 1266 86 1322
rect 142 1266 210 1322
rect 266 1320 903 1322
rect 959 1320 1045 1376
rect 1101 1320 1444 1376
rect 1500 1320 1586 1376
rect 1642 1320 1984 1376
rect 2040 1320 2126 1376
rect 2182 1320 2521 1376
rect 2577 1320 2663 1376
rect 2719 1320 3058 1376
rect 3114 1320 3200 1376
rect 3256 1320 3602 1376
rect 3658 1320 3744 1376
rect 3800 1320 4138 1376
rect 4194 1320 4280 1376
rect 4336 1320 4678 1376
rect 4734 1320 4820 1376
rect 4876 1320 5215 1376
rect 5271 1320 5357 1376
rect 5413 1320 5760 1376
rect 5816 1320 5902 1376
rect 5958 1320 6300 1376
rect 6356 1320 6442 1376
rect 6498 1320 6845 1376
rect 6901 1320 6987 1376
rect 7043 1320 7382 1376
rect 7438 1320 7524 1376
rect 7580 1320 7919 1376
rect 7975 1320 8061 1376
rect 8117 1320 8462 1376
rect 8518 1320 8604 1376
rect 8660 1320 9004 1376
rect 9060 1320 9146 1376
rect 9202 1320 9547 1376
rect 9603 1320 9689 1376
rect 9745 1320 10081 1376
rect 10137 1320 10223 1376
rect 10279 1320 10622 1376
rect 10678 1320 10764 1376
rect 10820 1320 11162 1376
rect 11218 1320 11304 1376
rect 11360 1320 11702 1376
rect 11758 1320 11844 1376
rect 11900 1322 13200 1376
rect 11900 1320 12526 1322
rect 266 1266 12526 1320
rect 12582 1266 12650 1322
rect 12706 1266 12774 1322
rect 12830 1266 12898 1322
rect 12954 1266 13022 1322
rect 13078 1266 13200 1322
rect -400 1234 13200 1266
rect -400 1198 903 1234
rect -400 1142 -286 1198
rect -230 1142 -162 1198
rect -106 1142 -38 1198
rect 18 1142 86 1198
rect 142 1142 210 1198
rect 266 1178 903 1198
rect 959 1178 1045 1234
rect 1101 1178 1444 1234
rect 1500 1178 1586 1234
rect 1642 1178 1984 1234
rect 2040 1178 2126 1234
rect 2182 1178 2521 1234
rect 2577 1178 2663 1234
rect 2719 1178 3058 1234
rect 3114 1178 3200 1234
rect 3256 1178 3602 1234
rect 3658 1178 3744 1234
rect 3800 1178 4138 1234
rect 4194 1178 4280 1234
rect 4336 1178 4678 1234
rect 4734 1178 4820 1234
rect 4876 1178 5215 1234
rect 5271 1178 5357 1234
rect 5413 1178 5760 1234
rect 5816 1178 5902 1234
rect 5958 1178 6300 1234
rect 6356 1178 6442 1234
rect 6498 1178 6845 1234
rect 6901 1178 6987 1234
rect 7043 1178 7382 1234
rect 7438 1178 7524 1234
rect 7580 1178 7919 1234
rect 7975 1178 8061 1234
rect 8117 1178 8462 1234
rect 8518 1178 8604 1234
rect 8660 1178 9004 1234
rect 9060 1178 9146 1234
rect 9202 1178 9547 1234
rect 9603 1178 9689 1234
rect 9745 1178 10081 1234
rect 10137 1178 10223 1234
rect 10279 1178 10622 1234
rect 10678 1178 10764 1234
rect 10820 1178 11162 1234
rect 11218 1178 11304 1234
rect 11360 1178 11702 1234
rect 11758 1178 11844 1234
rect 11900 1198 13200 1234
rect 11900 1178 12526 1198
rect 266 1142 12526 1178
rect 12582 1142 12650 1198
rect 12706 1142 12774 1198
rect 12830 1142 12898 1198
rect 12954 1142 13022 1198
rect 13078 1142 13200 1198
rect -400 1092 13200 1142
rect -400 1074 903 1092
rect -400 1018 -286 1074
rect -230 1018 -162 1074
rect -106 1018 -38 1074
rect 18 1018 86 1074
rect 142 1018 210 1074
rect 266 1036 903 1074
rect 959 1036 1045 1092
rect 1101 1036 1444 1092
rect 1500 1036 1586 1092
rect 1642 1036 1984 1092
rect 2040 1036 2126 1092
rect 2182 1036 2521 1092
rect 2577 1036 2663 1092
rect 2719 1036 3058 1092
rect 3114 1036 3200 1092
rect 3256 1036 3602 1092
rect 3658 1036 3744 1092
rect 3800 1036 4138 1092
rect 4194 1036 4280 1092
rect 4336 1036 4678 1092
rect 4734 1036 4820 1092
rect 4876 1036 5215 1092
rect 5271 1036 5357 1092
rect 5413 1036 5760 1092
rect 5816 1036 5902 1092
rect 5958 1036 6300 1092
rect 6356 1036 6442 1092
rect 6498 1036 6845 1092
rect 6901 1036 6987 1092
rect 7043 1036 7382 1092
rect 7438 1036 7524 1092
rect 7580 1036 7919 1092
rect 7975 1036 8061 1092
rect 8117 1036 8462 1092
rect 8518 1036 8604 1092
rect 8660 1036 9004 1092
rect 9060 1036 9146 1092
rect 9202 1036 9547 1092
rect 9603 1036 9689 1092
rect 9745 1036 10081 1092
rect 10137 1036 10223 1092
rect 10279 1036 10622 1092
rect 10678 1036 10764 1092
rect 10820 1036 11162 1092
rect 11218 1036 11304 1092
rect 11360 1036 11702 1092
rect 11758 1036 11844 1092
rect 11900 1074 13200 1092
rect 11900 1036 12526 1074
rect 266 1018 12526 1036
rect 12582 1018 12650 1074
rect 12706 1018 12774 1074
rect 12830 1018 12898 1074
rect 12954 1018 13022 1074
rect 13078 1018 13200 1074
rect -400 950 13200 1018
rect -400 894 -286 950
rect -230 894 -162 950
rect -106 894 -38 950
rect 18 894 86 950
rect 142 894 210 950
rect 266 894 903 950
rect 959 894 1045 950
rect 1101 894 1444 950
rect 1500 894 1586 950
rect 1642 894 1984 950
rect 2040 894 2126 950
rect 2182 894 2521 950
rect 2577 894 2663 950
rect 2719 894 3058 950
rect 3114 894 3200 950
rect 3256 894 3602 950
rect 3658 894 3744 950
rect 3800 894 4138 950
rect 4194 894 4280 950
rect 4336 894 4678 950
rect 4734 894 4820 950
rect 4876 894 5215 950
rect 5271 894 5357 950
rect 5413 894 5760 950
rect 5816 894 5902 950
rect 5958 894 6300 950
rect 6356 894 6442 950
rect 6498 894 6845 950
rect 6901 894 6987 950
rect 7043 894 7382 950
rect 7438 894 7524 950
rect 7580 894 7919 950
rect 7975 894 8061 950
rect 8117 894 8462 950
rect 8518 894 8604 950
rect 8660 894 9004 950
rect 9060 894 9146 950
rect 9202 894 9547 950
rect 9603 894 9689 950
rect 9745 894 10081 950
rect 10137 894 10223 950
rect 10279 894 10622 950
rect 10678 894 10764 950
rect 10820 894 11162 950
rect 11218 894 11304 950
rect 11360 894 11702 950
rect 11758 894 11844 950
rect 11900 894 12526 950
rect 12582 894 12650 950
rect 12706 894 12774 950
rect 12830 894 12898 950
rect 12954 894 13022 950
rect 13078 894 13200 950
rect -400 826 13200 894
rect -400 770 -286 826
rect -230 770 -162 826
rect -106 770 -38 826
rect 18 770 86 826
rect 142 770 210 826
rect 266 808 12526 826
rect 266 770 903 808
rect -400 752 903 770
rect 959 752 1045 808
rect 1101 752 1444 808
rect 1500 752 1586 808
rect 1642 752 1984 808
rect 2040 752 2126 808
rect 2182 752 2521 808
rect 2577 752 2663 808
rect 2719 752 3058 808
rect 3114 752 3200 808
rect 3256 752 3602 808
rect 3658 752 3744 808
rect 3800 752 4138 808
rect 4194 752 4280 808
rect 4336 752 4678 808
rect 4734 752 4820 808
rect 4876 752 5215 808
rect 5271 752 5357 808
rect 5413 752 5760 808
rect 5816 752 5902 808
rect 5958 752 6300 808
rect 6356 752 6442 808
rect 6498 752 6845 808
rect 6901 752 6987 808
rect 7043 752 7382 808
rect 7438 752 7524 808
rect 7580 752 7919 808
rect 7975 752 8061 808
rect 8117 752 8462 808
rect 8518 752 8604 808
rect 8660 752 9004 808
rect 9060 752 9146 808
rect 9202 752 9547 808
rect 9603 752 9689 808
rect 9745 752 10081 808
rect 10137 752 10223 808
rect 10279 752 10622 808
rect 10678 752 10764 808
rect 10820 752 11162 808
rect 11218 752 11304 808
rect 11360 752 11702 808
rect 11758 752 11844 808
rect 11900 770 12526 808
rect 12582 770 12650 826
rect 12706 770 12774 826
rect 12830 770 12898 826
rect 12954 770 13022 826
rect 13078 770 13200 826
rect 11900 752 13200 770
rect -400 702 13200 752
rect -400 646 -286 702
rect -230 646 -162 702
rect -106 646 -38 702
rect 18 646 86 702
rect 142 646 210 702
rect 266 666 12526 702
rect 266 646 903 666
rect -400 610 903 646
rect 959 610 1045 666
rect 1101 610 1444 666
rect 1500 610 1586 666
rect 1642 610 1984 666
rect 2040 610 2126 666
rect 2182 610 2521 666
rect 2577 610 2663 666
rect 2719 610 3058 666
rect 3114 610 3200 666
rect 3256 610 3602 666
rect 3658 610 3744 666
rect 3800 610 4138 666
rect 4194 610 4280 666
rect 4336 610 4678 666
rect 4734 610 4820 666
rect 4876 610 5215 666
rect 5271 610 5357 666
rect 5413 610 5760 666
rect 5816 610 5902 666
rect 5958 610 6300 666
rect 6356 610 6442 666
rect 6498 610 6845 666
rect 6901 610 6987 666
rect 7043 610 7382 666
rect 7438 610 7524 666
rect 7580 610 7919 666
rect 7975 610 8061 666
rect 8117 610 8462 666
rect 8518 610 8604 666
rect 8660 610 9004 666
rect 9060 610 9146 666
rect 9202 610 9547 666
rect 9603 610 9689 666
rect 9745 610 10081 666
rect 10137 610 10223 666
rect 10279 610 10622 666
rect 10678 610 10764 666
rect 10820 610 11162 666
rect 11218 610 11304 666
rect 11360 610 11702 666
rect 11758 610 11844 666
rect 11900 646 12526 666
rect 12582 646 12650 702
rect 12706 646 12774 702
rect 12830 646 12898 702
rect 12954 646 13022 702
rect 13078 646 13200 702
rect 11900 610 13200 646
rect -400 578 13200 610
rect -400 522 -286 578
rect -230 522 -162 578
rect -106 522 -38 578
rect 18 522 86 578
rect 142 522 210 578
rect 266 524 12526 578
rect 266 522 903 524
rect -400 468 903 522
rect 959 468 1045 524
rect 1101 468 1444 524
rect 1500 468 1586 524
rect 1642 468 1984 524
rect 2040 468 2126 524
rect 2182 468 2521 524
rect 2577 468 2663 524
rect 2719 468 3058 524
rect 3114 468 3200 524
rect 3256 468 3602 524
rect 3658 468 3744 524
rect 3800 468 4138 524
rect 4194 468 4280 524
rect 4336 468 4678 524
rect 4734 468 4820 524
rect 4876 468 5215 524
rect 5271 468 5357 524
rect 5413 468 5760 524
rect 5816 468 5902 524
rect 5958 468 6300 524
rect 6356 468 6442 524
rect 6498 468 6845 524
rect 6901 468 6987 524
rect 7043 468 7382 524
rect 7438 468 7524 524
rect 7580 468 7919 524
rect 7975 468 8061 524
rect 8117 468 8462 524
rect 8518 468 8604 524
rect 8660 468 9004 524
rect 9060 468 9146 524
rect 9202 468 9547 524
rect 9603 468 9689 524
rect 9745 468 10081 524
rect 10137 468 10223 524
rect 10279 468 10622 524
rect 10678 468 10764 524
rect 10820 468 11162 524
rect 11218 468 11304 524
rect 11360 468 11702 524
rect 11758 468 11844 524
rect 11900 522 12526 524
rect 12582 522 12650 578
rect 12706 522 12774 578
rect 12830 522 12898 578
rect 12954 522 13022 578
rect 13078 522 13200 578
rect 11900 468 13200 522
rect -400 454 13200 468
rect -400 398 -286 454
rect -230 398 -162 454
rect -106 398 -38 454
rect 18 398 86 454
rect 142 398 210 454
rect 266 398 12526 454
rect 12582 398 12650 454
rect 12706 398 12774 454
rect 12830 398 12898 454
rect 12954 398 13022 454
rect 13078 398 13200 454
rect -400 330 13200 398
rect -400 274 -286 330
rect -230 274 -162 330
rect -106 274 -38 330
rect 18 274 86 330
rect 142 274 210 330
rect 266 302 12526 330
rect 266 274 415 302
rect -400 246 415 274
rect 471 246 557 302
rect 613 246 699 302
rect 755 246 841 302
rect 897 246 983 302
rect 1039 246 1125 302
rect 1181 246 1267 302
rect 1323 246 1409 302
rect 1465 246 1551 302
rect 1607 246 1693 302
rect 1749 246 1835 302
rect 1891 246 1977 302
rect 2033 246 2119 302
rect 2175 246 2261 302
rect 2317 246 2403 302
rect 2459 246 2545 302
rect 2601 246 2687 302
rect 2743 246 2829 302
rect 2885 246 2971 302
rect 3027 246 3113 302
rect 3169 246 3255 302
rect 3311 246 3397 302
rect 3453 246 3539 302
rect 3595 246 3681 302
rect 3737 246 3823 302
rect 3879 246 3965 302
rect 4021 246 4107 302
rect 4163 246 4249 302
rect 4305 246 4391 302
rect 4447 246 4533 302
rect 4589 246 4675 302
rect 4731 246 4817 302
rect 4873 246 4959 302
rect 5015 246 5101 302
rect 5157 246 5243 302
rect 5299 246 5385 302
rect 5441 246 5527 302
rect 5583 246 5669 302
rect 5725 246 5811 302
rect 5867 246 5953 302
rect 6009 246 6095 302
rect 6151 246 6237 302
rect 6293 246 6379 302
rect 6435 246 6521 302
rect 6577 246 6663 302
rect 6719 246 6805 302
rect 6861 246 6947 302
rect 7003 246 7089 302
rect 7145 246 7231 302
rect 7287 246 7373 302
rect 7429 246 7515 302
rect 7571 246 7657 302
rect 7713 246 7799 302
rect 7855 246 7941 302
rect 7997 246 8083 302
rect 8139 246 8225 302
rect 8281 246 8367 302
rect 8423 246 8509 302
rect 8565 246 8651 302
rect 8707 246 8793 302
rect 8849 246 8935 302
rect 8991 246 9077 302
rect 9133 246 9219 302
rect 9275 246 9361 302
rect 9417 246 9503 302
rect 9559 246 9645 302
rect 9701 246 9787 302
rect 9843 246 9929 302
rect 9985 246 10071 302
rect 10127 246 10213 302
rect 10269 246 10355 302
rect 10411 246 10497 302
rect 10553 246 10639 302
rect 10695 246 10781 302
rect 10837 246 10923 302
rect 10979 246 11065 302
rect 11121 246 11207 302
rect 11263 246 11349 302
rect 11405 246 11491 302
rect 11547 246 11633 302
rect 11689 246 11775 302
rect 11831 246 11917 302
rect 11973 246 12059 302
rect 12115 246 12201 302
rect 12257 246 12343 302
rect 12399 274 12526 302
rect 12582 274 12650 330
rect 12706 274 12774 330
rect 12830 274 12898 330
rect 12954 274 13022 330
rect 13078 274 13200 330
rect 12399 246 13200 274
rect -400 206 13200 246
rect -400 150 -286 206
rect -230 150 -162 206
rect -106 150 -38 206
rect 18 150 86 206
rect 142 150 210 206
rect 266 160 12526 206
rect 266 150 415 160
rect -400 104 415 150
rect 471 104 557 160
rect 613 104 699 160
rect 755 104 841 160
rect 897 104 983 160
rect 1039 104 1125 160
rect 1181 104 1267 160
rect 1323 104 1409 160
rect 1465 104 1551 160
rect 1607 104 1693 160
rect 1749 104 1835 160
rect 1891 104 1977 160
rect 2033 104 2119 160
rect 2175 104 2261 160
rect 2317 104 2403 160
rect 2459 104 2545 160
rect 2601 104 2687 160
rect 2743 104 2829 160
rect 2885 104 2971 160
rect 3027 104 3113 160
rect 3169 104 3255 160
rect 3311 104 3397 160
rect 3453 104 3539 160
rect 3595 104 3681 160
rect 3737 104 3823 160
rect 3879 104 3965 160
rect 4021 104 4107 160
rect 4163 104 4249 160
rect 4305 104 4391 160
rect 4447 104 4533 160
rect 4589 104 4675 160
rect 4731 104 4817 160
rect 4873 104 4959 160
rect 5015 104 5101 160
rect 5157 104 5243 160
rect 5299 104 5385 160
rect 5441 104 5527 160
rect 5583 104 5669 160
rect 5725 104 5811 160
rect 5867 104 5953 160
rect 6009 104 6095 160
rect 6151 104 6237 160
rect 6293 104 6379 160
rect 6435 104 6521 160
rect 6577 104 6663 160
rect 6719 104 6805 160
rect 6861 104 6947 160
rect 7003 104 7089 160
rect 7145 104 7231 160
rect 7287 104 7373 160
rect 7429 104 7515 160
rect 7571 104 7657 160
rect 7713 104 7799 160
rect 7855 104 7941 160
rect 7997 104 8083 160
rect 8139 104 8225 160
rect 8281 104 8367 160
rect 8423 104 8509 160
rect 8565 104 8651 160
rect 8707 104 8793 160
rect 8849 104 8935 160
rect 8991 104 9077 160
rect 9133 104 9219 160
rect 9275 104 9361 160
rect 9417 104 9503 160
rect 9559 104 9645 160
rect 9701 104 9787 160
rect 9843 104 9929 160
rect 9985 104 10071 160
rect 10127 104 10213 160
rect 10269 104 10355 160
rect 10411 104 10497 160
rect 10553 104 10639 160
rect 10695 104 10781 160
rect 10837 104 10923 160
rect 10979 104 11065 160
rect 11121 104 11207 160
rect 11263 104 11349 160
rect 11405 104 11491 160
rect 11547 104 11633 160
rect 11689 104 11775 160
rect 11831 104 11917 160
rect 11973 104 12059 160
rect 12115 104 12201 160
rect 12257 104 12343 160
rect 12399 150 12526 160
rect 12582 150 12650 206
rect 12706 150 12774 206
rect 12830 150 12898 206
rect 12954 150 13022 206
rect 13078 150 13200 206
rect 12399 104 13200 150
rect -400 0 13200 104
<< glass >>
rect 400 400 12400 12400
<< end >>
