magic
tech gf180mcuD
timestamp 1768559988
<< nwell >>
rect -33 -9 32 38
<< nmos >>
rect 0 -31 6 -19
<< pmos >>
rect 0 0 6 24
<< ndiff >>
rect -5 -31 0 -19
rect 6 -31 11 -19
<< pdiff >>
rect -18 15 0 24
rect -18 9 -13 15
rect -7 9 0 15
rect -18 0 0 9
rect 6 0 11 24
<< pdiffc >>
rect -13 9 -7 15
<< polysilicon >>
rect 0 24 6 29
rect 0 -19 6 0
rect 0 -36 6 -31
<< metal1 >>
rect -33 29 32 38
rect -13 15 -7 29
rect -13 7 -7 9
<< end >>
