magic
tech gf180mcuD
magscale 1 5
timestamp 1764281188
use pmos_6p0_esd  pmos_6p0_esd_0
timestamp 1764281188
transform -1 0 1040 0 1 0
box 0 6 598 6126
use pmos_6p0_esd  pmos_6p0_esd_1
timestamp 1764281188
transform 1 0 0 0 1 0
box 0 6 598 6126
<< end >>
