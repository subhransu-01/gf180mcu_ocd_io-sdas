magic
tech gf180mcuD
magscale 1 10
timestamp 1764347740
<< psubdiff >>
rect 13097 70975 69968 71000
rect 13097 70929 13119 70975
rect 13165 70929 13223 70975
rect 13269 70929 13377 70975
rect 13423 70929 13481 70975
rect 13527 70929 13585 70975
rect 13631 70929 13689 70975
rect 13735 70929 13793 70975
rect 13839 70929 13897 70975
rect 13943 70929 14001 70975
rect 14047 70929 14105 70975
rect 14151 70929 14209 70975
rect 14255 70929 14313 70975
rect 14359 70929 14417 70975
rect 14463 70929 14521 70975
rect 14567 70929 14625 70975
rect 14671 70929 14729 70975
rect 14775 70929 14833 70975
rect 14879 70929 14937 70975
rect 14983 70929 15041 70975
rect 15087 70929 15145 70975
rect 15191 70929 15249 70975
rect 15295 70929 15353 70975
rect 15399 70929 15457 70975
rect 15503 70929 15561 70975
rect 15607 70929 15665 70975
rect 15711 70929 15769 70975
rect 15815 70929 15873 70975
rect 15919 70929 15977 70975
rect 16023 70929 16081 70975
rect 16127 70929 16185 70975
rect 16231 70929 16289 70975
rect 16335 70929 16393 70975
rect 16439 70929 16497 70975
rect 16543 70929 16601 70975
rect 16647 70929 16705 70975
rect 16751 70929 16809 70975
rect 16855 70929 16913 70975
rect 16959 70929 17017 70975
rect 17063 70929 17121 70975
rect 17167 70929 17225 70975
rect 17271 70929 17329 70975
rect 17375 70929 17433 70975
rect 17479 70929 17537 70975
rect 17583 70929 17641 70975
rect 17687 70929 17745 70975
rect 17791 70929 17849 70975
rect 17895 70929 17953 70975
rect 17999 70929 18057 70975
rect 18103 70929 18161 70975
rect 18207 70929 18265 70975
rect 18311 70929 18369 70975
rect 18415 70929 18473 70975
rect 18519 70929 18577 70975
rect 18623 70929 18681 70975
rect 18727 70929 18785 70975
rect 18831 70929 18889 70975
rect 18935 70929 18993 70975
rect 19039 70929 19097 70975
rect 19143 70929 19201 70975
rect 19247 70929 19305 70975
rect 19351 70929 19409 70975
rect 19455 70929 19513 70975
rect 19559 70929 19617 70975
rect 19663 70929 19721 70975
rect 19767 70929 19825 70975
rect 19871 70929 19929 70975
rect 19975 70929 20033 70975
rect 20079 70929 20137 70975
rect 20183 70929 20241 70975
rect 20287 70929 20345 70975
rect 20391 70929 20449 70975
rect 20495 70929 20553 70975
rect 20599 70929 20657 70975
rect 20703 70929 20761 70975
rect 20807 70929 20865 70975
rect 20911 70929 20969 70975
rect 21015 70929 21073 70975
rect 21119 70929 21177 70975
rect 21223 70929 21281 70975
rect 21327 70929 21385 70975
rect 21431 70929 21489 70975
rect 21535 70929 21593 70975
rect 21639 70929 21697 70975
rect 21743 70929 21801 70975
rect 21847 70929 21905 70975
rect 21951 70929 22009 70975
rect 22055 70929 22113 70975
rect 22159 70929 22217 70975
rect 22263 70929 22321 70975
rect 22367 70929 22425 70975
rect 22471 70929 22529 70975
rect 22575 70929 22633 70975
rect 22679 70929 22737 70975
rect 22783 70929 22841 70975
rect 22887 70929 22945 70975
rect 22991 70929 23049 70975
rect 23095 70929 23153 70975
rect 23199 70929 23257 70975
rect 23303 70929 23361 70975
rect 23407 70929 23465 70975
rect 23511 70929 23569 70975
rect 23615 70929 23673 70975
rect 23719 70929 23777 70975
rect 23823 70929 23881 70975
rect 23927 70929 23985 70975
rect 24031 70929 24089 70975
rect 24135 70929 24193 70975
rect 24239 70929 24297 70975
rect 24343 70929 24401 70975
rect 24447 70929 24505 70975
rect 24551 70929 24609 70975
rect 24655 70929 24713 70975
rect 24759 70929 24817 70975
rect 24863 70929 24921 70975
rect 24967 70929 25025 70975
rect 25071 70929 25129 70975
rect 25175 70929 25233 70975
rect 25279 70929 25337 70975
rect 25383 70929 25441 70975
rect 25487 70929 25545 70975
rect 25591 70929 25649 70975
rect 25695 70929 25753 70975
rect 25799 70929 25857 70975
rect 25903 70929 25961 70975
rect 26007 70929 26065 70975
rect 26111 70929 26169 70975
rect 26215 70929 26273 70975
rect 26319 70929 26377 70975
rect 26423 70929 26481 70975
rect 26527 70929 26585 70975
rect 26631 70929 26689 70975
rect 26735 70929 26793 70975
rect 26839 70929 26897 70975
rect 26943 70929 27001 70975
rect 27047 70929 27105 70975
rect 27151 70929 27209 70975
rect 27255 70929 27313 70975
rect 27359 70929 27417 70975
rect 27463 70929 27521 70975
rect 27567 70929 27625 70975
rect 27671 70929 27729 70975
rect 27775 70929 27833 70975
rect 27879 70929 27937 70975
rect 27983 70929 28041 70975
rect 28087 70929 28145 70975
rect 28191 70929 28249 70975
rect 28295 70929 28353 70975
rect 28399 70929 28457 70975
rect 28503 70929 28561 70975
rect 28607 70929 28665 70975
rect 28711 70929 28769 70975
rect 28815 70929 28873 70975
rect 28919 70929 28977 70975
rect 29023 70929 29081 70975
rect 29127 70929 29185 70975
rect 29231 70929 29289 70975
rect 29335 70929 29393 70975
rect 29439 70929 29497 70975
rect 29543 70929 29601 70975
rect 29647 70929 29705 70975
rect 29751 70929 29809 70975
rect 29855 70929 29913 70975
rect 29959 70929 30017 70975
rect 30063 70929 30121 70975
rect 30167 70929 30225 70975
rect 30271 70929 30329 70975
rect 30375 70929 30433 70975
rect 30479 70929 30537 70975
rect 30583 70929 30641 70975
rect 30687 70929 30745 70975
rect 30791 70929 30849 70975
rect 30895 70929 30953 70975
rect 30999 70929 31057 70975
rect 31103 70929 31161 70975
rect 31207 70929 31265 70975
rect 31311 70929 31369 70975
rect 31415 70929 31473 70975
rect 31519 70929 31577 70975
rect 31623 70929 31681 70975
rect 31727 70929 31785 70975
rect 31831 70929 31889 70975
rect 31935 70929 31993 70975
rect 32039 70929 32097 70975
rect 32143 70929 32201 70975
rect 32247 70929 32305 70975
rect 32351 70929 32409 70975
rect 32455 70929 32513 70975
rect 32559 70929 32617 70975
rect 32663 70929 32721 70975
rect 32767 70929 32825 70975
rect 32871 70929 32929 70975
rect 32975 70929 33033 70975
rect 33079 70929 33137 70975
rect 33183 70929 33241 70975
rect 33287 70929 33345 70975
rect 33391 70929 33449 70975
rect 33495 70929 33553 70975
rect 33599 70929 33657 70975
rect 33703 70929 33761 70975
rect 33807 70929 33865 70975
rect 33911 70929 33969 70975
rect 34015 70929 34073 70975
rect 34119 70929 34177 70975
rect 34223 70929 34281 70975
rect 34327 70929 34385 70975
rect 34431 70929 34489 70975
rect 34535 70929 34593 70975
rect 34639 70929 34697 70975
rect 34743 70929 34801 70975
rect 34847 70929 34905 70975
rect 34951 70929 35009 70975
rect 35055 70929 35113 70975
rect 35159 70929 35217 70975
rect 35263 70929 35321 70975
rect 35367 70929 35425 70975
rect 35471 70929 35529 70975
rect 35575 70929 35633 70975
rect 35679 70929 35737 70975
rect 35783 70929 35841 70975
rect 35887 70929 35945 70975
rect 35991 70929 36049 70975
rect 36095 70929 36153 70975
rect 36199 70929 36257 70975
rect 36303 70929 36361 70975
rect 36407 70929 36465 70975
rect 36511 70929 36569 70975
rect 36615 70929 36673 70975
rect 36719 70929 36777 70975
rect 36823 70929 36881 70975
rect 36927 70929 36985 70975
rect 37031 70929 37089 70975
rect 37135 70929 37193 70975
rect 37239 70929 37297 70975
rect 37343 70929 37401 70975
rect 37447 70929 37505 70975
rect 37551 70929 37609 70975
rect 37655 70929 37713 70975
rect 37759 70929 37817 70975
rect 37863 70929 37921 70975
rect 37967 70929 38025 70975
rect 38071 70929 38129 70975
rect 38175 70929 38233 70975
rect 38279 70929 38337 70975
rect 38383 70929 38441 70975
rect 38487 70929 38545 70975
rect 38591 70929 38649 70975
rect 38695 70929 38753 70975
rect 38799 70929 38857 70975
rect 38903 70929 38961 70975
rect 39007 70929 39065 70975
rect 39111 70929 39169 70975
rect 39215 70929 39273 70975
rect 39319 70929 39377 70975
rect 39423 70929 39481 70975
rect 39527 70929 39585 70975
rect 39631 70929 39689 70975
rect 39735 70929 39793 70975
rect 39839 70929 39897 70975
rect 39943 70929 40001 70975
rect 40047 70929 40105 70975
rect 40151 70929 40209 70975
rect 40255 70929 40313 70975
rect 40359 70929 40417 70975
rect 40463 70929 40521 70975
rect 40567 70929 40625 70975
rect 40671 70929 40729 70975
rect 40775 70929 40833 70975
rect 40879 70929 40937 70975
rect 40983 70929 41041 70975
rect 41087 70929 41145 70975
rect 41191 70929 41249 70975
rect 41295 70929 41353 70975
rect 41399 70929 41457 70975
rect 41503 70929 41561 70975
rect 41607 70929 41665 70975
rect 41711 70929 41769 70975
rect 41815 70929 41873 70975
rect 41919 70929 41977 70975
rect 42023 70929 42081 70975
rect 42127 70929 42185 70975
rect 42231 70929 42289 70975
rect 42335 70929 42393 70975
rect 42439 70929 42497 70975
rect 42543 70929 42601 70975
rect 42647 70929 42705 70975
rect 42751 70929 42809 70975
rect 42855 70929 42913 70975
rect 42959 70929 43017 70975
rect 43063 70929 43121 70975
rect 43167 70929 43225 70975
rect 43271 70929 43329 70975
rect 43375 70929 43433 70975
rect 43479 70929 43537 70975
rect 43583 70929 43641 70975
rect 43687 70929 43745 70975
rect 43791 70929 43849 70975
rect 43895 70929 43953 70975
rect 43999 70929 44057 70975
rect 44103 70929 44161 70975
rect 44207 70929 44265 70975
rect 44311 70929 44369 70975
rect 44415 70929 44473 70975
rect 44519 70929 44577 70975
rect 44623 70929 44681 70975
rect 44727 70929 44785 70975
rect 44831 70929 44889 70975
rect 44935 70929 44993 70975
rect 45039 70929 45097 70975
rect 45143 70929 45201 70975
rect 45247 70929 45305 70975
rect 45351 70929 45409 70975
rect 45455 70929 45513 70975
rect 45559 70929 45617 70975
rect 45663 70929 45721 70975
rect 45767 70929 45825 70975
rect 45871 70929 45929 70975
rect 45975 70929 46033 70975
rect 46079 70929 46137 70975
rect 46183 70929 46241 70975
rect 46287 70929 46345 70975
rect 46391 70929 46449 70975
rect 46495 70929 46553 70975
rect 46599 70929 46657 70975
rect 46703 70929 46761 70975
rect 46807 70929 46865 70975
rect 46911 70929 46969 70975
rect 47015 70929 47073 70975
rect 47119 70929 47177 70975
rect 47223 70929 47281 70975
rect 47327 70929 47385 70975
rect 47431 70929 47489 70975
rect 47535 70929 47593 70975
rect 47639 70929 47697 70975
rect 47743 70929 47801 70975
rect 47847 70929 47905 70975
rect 47951 70929 48009 70975
rect 48055 70929 48113 70975
rect 48159 70929 48217 70975
rect 48263 70929 48321 70975
rect 48367 70929 48425 70975
rect 48471 70929 48529 70975
rect 48575 70929 48633 70975
rect 48679 70929 48737 70975
rect 48783 70929 48841 70975
rect 48887 70929 48945 70975
rect 48991 70929 49049 70975
rect 49095 70929 49153 70975
rect 49199 70929 49257 70975
rect 49303 70929 49361 70975
rect 49407 70929 49465 70975
rect 49511 70929 49569 70975
rect 49615 70929 49673 70975
rect 49719 70929 49777 70975
rect 49823 70929 49881 70975
rect 49927 70929 49985 70975
rect 50031 70929 50089 70975
rect 50135 70929 50193 70975
rect 50239 70929 50297 70975
rect 50343 70929 50401 70975
rect 50447 70929 50505 70975
rect 50551 70929 50609 70975
rect 50655 70929 50713 70975
rect 50759 70929 50817 70975
rect 50863 70929 50921 70975
rect 50967 70929 51025 70975
rect 51071 70929 51129 70975
rect 51175 70929 51233 70975
rect 51279 70929 51337 70975
rect 51383 70929 51441 70975
rect 51487 70929 51545 70975
rect 51591 70929 51649 70975
rect 51695 70929 51753 70975
rect 51799 70929 51857 70975
rect 51903 70929 51961 70975
rect 52007 70929 52065 70975
rect 52111 70929 52169 70975
rect 52215 70929 52273 70975
rect 52319 70929 52377 70975
rect 52423 70929 52481 70975
rect 52527 70929 52585 70975
rect 52631 70929 52689 70975
rect 52735 70929 52793 70975
rect 52839 70929 52897 70975
rect 52943 70929 53001 70975
rect 53047 70929 53105 70975
rect 53151 70929 53209 70975
rect 53255 70929 53313 70975
rect 53359 70929 53417 70975
rect 53463 70929 53521 70975
rect 53567 70929 53625 70975
rect 53671 70929 53729 70975
rect 53775 70929 53833 70975
rect 53879 70929 53937 70975
rect 53983 70929 54041 70975
rect 54087 70929 54145 70975
rect 54191 70929 54249 70975
rect 54295 70929 54353 70975
rect 54399 70929 54457 70975
rect 54503 70929 54561 70975
rect 54607 70929 54665 70975
rect 54711 70929 54769 70975
rect 54815 70929 54873 70975
rect 54919 70929 54977 70975
rect 55023 70929 55081 70975
rect 55127 70929 55185 70975
rect 55231 70929 55289 70975
rect 55335 70929 55393 70975
rect 55439 70929 55497 70975
rect 55543 70929 55601 70975
rect 55647 70929 55705 70975
rect 55751 70929 55809 70975
rect 55855 70929 55913 70975
rect 55959 70929 56017 70975
rect 56063 70929 56121 70975
rect 56167 70929 56225 70975
rect 56271 70929 56329 70975
rect 56375 70929 56433 70975
rect 56479 70929 56537 70975
rect 56583 70929 56641 70975
rect 56687 70929 56745 70975
rect 56791 70929 56849 70975
rect 56895 70929 56953 70975
rect 56999 70929 57057 70975
rect 57103 70929 57161 70975
rect 57207 70929 57265 70975
rect 57311 70929 57369 70975
rect 57415 70929 57473 70975
rect 57519 70929 57577 70975
rect 57623 70929 57681 70975
rect 57727 70929 57785 70975
rect 57831 70929 57889 70975
rect 57935 70929 57993 70975
rect 58039 70929 58097 70975
rect 58143 70929 58201 70975
rect 58247 70929 58305 70975
rect 58351 70929 58409 70975
rect 58455 70929 58513 70975
rect 58559 70929 58617 70975
rect 58663 70929 58721 70975
rect 58767 70929 58825 70975
rect 58871 70929 58929 70975
rect 58975 70929 59033 70975
rect 59079 70929 59137 70975
rect 59183 70929 59241 70975
rect 59287 70929 59345 70975
rect 59391 70929 59449 70975
rect 59495 70929 59553 70975
rect 59599 70929 59657 70975
rect 59703 70929 59761 70975
rect 59807 70929 59865 70975
rect 59911 70929 59969 70975
rect 60015 70929 60073 70975
rect 60119 70929 60177 70975
rect 60223 70929 60281 70975
rect 60327 70929 60385 70975
rect 60431 70929 60489 70975
rect 60535 70929 60593 70975
rect 60639 70929 60697 70975
rect 60743 70929 60801 70975
rect 60847 70929 60905 70975
rect 60951 70929 61009 70975
rect 61055 70929 61113 70975
rect 61159 70929 61217 70975
rect 61263 70929 61321 70975
rect 61367 70929 61425 70975
rect 61471 70929 61529 70975
rect 61575 70929 61633 70975
rect 61679 70929 61737 70975
rect 61783 70929 61841 70975
rect 61887 70929 61945 70975
rect 61991 70929 62049 70975
rect 62095 70929 62153 70975
rect 62199 70929 62257 70975
rect 62303 70929 62361 70975
rect 62407 70929 62465 70975
rect 62511 70929 62569 70975
rect 62615 70929 62673 70975
rect 62719 70929 62777 70975
rect 62823 70929 62881 70975
rect 62927 70929 62985 70975
rect 63031 70929 63089 70975
rect 63135 70929 63193 70975
rect 63239 70929 63297 70975
rect 63343 70929 63401 70975
rect 63447 70929 63505 70975
rect 63551 70929 63609 70975
rect 63655 70929 63713 70975
rect 63759 70929 63817 70975
rect 63863 70929 63921 70975
rect 63967 70929 64025 70975
rect 64071 70929 64129 70975
rect 64175 70929 64233 70975
rect 64279 70929 64337 70975
rect 64383 70929 64441 70975
rect 64487 70929 64545 70975
rect 64591 70929 64649 70975
rect 64695 70929 64753 70975
rect 64799 70929 64857 70975
rect 64903 70929 64961 70975
rect 65007 70929 65065 70975
rect 65111 70929 65169 70975
rect 65215 70929 65273 70975
rect 65319 70929 65377 70975
rect 65423 70929 65481 70975
rect 65527 70929 65585 70975
rect 65631 70929 65689 70975
rect 65735 70929 65793 70975
rect 65839 70929 65897 70975
rect 65943 70929 66001 70975
rect 66047 70929 66105 70975
rect 66151 70929 66209 70975
rect 66255 70929 66313 70975
rect 66359 70929 66417 70975
rect 66463 70929 66521 70975
rect 66567 70929 66625 70975
rect 66671 70929 66729 70975
rect 66775 70929 66833 70975
rect 66879 70929 66937 70975
rect 66983 70929 67041 70975
rect 67087 70929 67145 70975
rect 67191 70929 67249 70975
rect 67295 70929 67353 70975
rect 67399 70929 67457 70975
rect 67503 70929 67561 70975
rect 67607 70929 67665 70975
rect 67711 70929 67769 70975
rect 67815 70929 67873 70975
rect 67919 70929 67977 70975
rect 68023 70929 68081 70975
rect 68127 70929 68185 70975
rect 68231 70929 68289 70975
rect 68335 70929 68393 70975
rect 68439 70929 68497 70975
rect 68543 70929 68601 70975
rect 68647 70929 68705 70975
rect 68751 70929 68809 70975
rect 68855 70929 68913 70975
rect 68959 70929 69017 70975
rect 69063 70929 69121 70975
rect 69167 70929 69225 70975
rect 69271 70929 69329 70975
rect 69375 70929 69433 70975
rect 69479 70929 69537 70975
rect 69583 70929 69641 70975
rect 69687 70929 69745 70975
rect 69791 70929 69849 70975
rect 69895 70929 69968 70975
rect 13097 70871 69968 70929
rect 13097 70825 13119 70871
rect 13165 70825 13223 70871
rect 13269 70825 13377 70871
rect 13423 70825 13481 70871
rect 13527 70825 13585 70871
rect 13631 70825 13689 70871
rect 13735 70825 13793 70871
rect 13839 70825 13897 70871
rect 13943 70825 14001 70871
rect 14047 70825 14105 70871
rect 14151 70825 14209 70871
rect 14255 70825 14313 70871
rect 14359 70825 14417 70871
rect 14463 70825 14521 70871
rect 14567 70825 14625 70871
rect 14671 70825 14729 70871
rect 14775 70825 14833 70871
rect 14879 70825 14937 70871
rect 14983 70825 15041 70871
rect 15087 70825 15145 70871
rect 15191 70825 15249 70871
rect 15295 70825 15353 70871
rect 15399 70825 15457 70871
rect 15503 70825 15561 70871
rect 15607 70825 15665 70871
rect 15711 70825 15769 70871
rect 15815 70825 15873 70871
rect 15919 70825 15977 70871
rect 16023 70825 16081 70871
rect 16127 70825 16185 70871
rect 16231 70825 16289 70871
rect 16335 70825 16393 70871
rect 16439 70825 16497 70871
rect 16543 70825 16601 70871
rect 16647 70825 16705 70871
rect 16751 70825 16809 70871
rect 16855 70825 16913 70871
rect 16959 70825 17017 70871
rect 17063 70825 17121 70871
rect 17167 70825 17225 70871
rect 17271 70825 17329 70871
rect 17375 70825 17433 70871
rect 17479 70825 17537 70871
rect 17583 70825 17641 70871
rect 17687 70825 17745 70871
rect 17791 70825 17849 70871
rect 17895 70825 17953 70871
rect 17999 70825 18057 70871
rect 18103 70825 18161 70871
rect 18207 70825 18265 70871
rect 18311 70825 18369 70871
rect 18415 70825 18473 70871
rect 18519 70825 18577 70871
rect 18623 70825 18681 70871
rect 18727 70825 18785 70871
rect 18831 70825 18889 70871
rect 18935 70825 18993 70871
rect 19039 70825 19097 70871
rect 19143 70825 19201 70871
rect 19247 70825 19305 70871
rect 19351 70825 19409 70871
rect 19455 70825 19513 70871
rect 19559 70825 19617 70871
rect 19663 70825 19721 70871
rect 19767 70825 19825 70871
rect 19871 70825 19929 70871
rect 19975 70825 20033 70871
rect 20079 70825 20137 70871
rect 20183 70825 20241 70871
rect 20287 70825 20345 70871
rect 20391 70825 20449 70871
rect 20495 70825 20553 70871
rect 20599 70825 20657 70871
rect 20703 70825 20761 70871
rect 20807 70825 20865 70871
rect 20911 70825 20969 70871
rect 21015 70825 21073 70871
rect 21119 70825 21177 70871
rect 21223 70825 21281 70871
rect 21327 70825 21385 70871
rect 21431 70825 21489 70871
rect 21535 70825 21593 70871
rect 21639 70825 21697 70871
rect 21743 70825 21801 70871
rect 21847 70825 21905 70871
rect 21951 70825 22009 70871
rect 22055 70825 22113 70871
rect 22159 70825 22217 70871
rect 22263 70825 22321 70871
rect 22367 70825 22425 70871
rect 22471 70825 22529 70871
rect 22575 70825 22633 70871
rect 22679 70825 22737 70871
rect 22783 70825 22841 70871
rect 22887 70825 22945 70871
rect 22991 70825 23049 70871
rect 23095 70825 23153 70871
rect 23199 70825 23257 70871
rect 23303 70825 23361 70871
rect 23407 70825 23465 70871
rect 23511 70825 23569 70871
rect 23615 70825 23673 70871
rect 23719 70825 23777 70871
rect 23823 70825 23881 70871
rect 23927 70825 23985 70871
rect 24031 70825 24089 70871
rect 24135 70825 24193 70871
rect 24239 70825 24297 70871
rect 24343 70825 24401 70871
rect 24447 70825 24505 70871
rect 24551 70825 24609 70871
rect 24655 70825 24713 70871
rect 24759 70825 24817 70871
rect 24863 70825 24921 70871
rect 24967 70825 25025 70871
rect 25071 70825 25129 70871
rect 25175 70825 25233 70871
rect 25279 70825 25337 70871
rect 25383 70825 25441 70871
rect 25487 70825 25545 70871
rect 25591 70825 25649 70871
rect 25695 70825 25753 70871
rect 25799 70825 25857 70871
rect 25903 70825 25961 70871
rect 26007 70825 26065 70871
rect 26111 70825 26169 70871
rect 26215 70825 26273 70871
rect 26319 70825 26377 70871
rect 26423 70825 26481 70871
rect 26527 70825 26585 70871
rect 26631 70825 26689 70871
rect 26735 70825 26793 70871
rect 26839 70825 26897 70871
rect 26943 70825 27001 70871
rect 27047 70825 27105 70871
rect 27151 70825 27209 70871
rect 27255 70825 27313 70871
rect 27359 70825 27417 70871
rect 27463 70825 27521 70871
rect 27567 70825 27625 70871
rect 27671 70825 27729 70871
rect 27775 70825 27833 70871
rect 27879 70825 27937 70871
rect 27983 70825 28041 70871
rect 28087 70825 28145 70871
rect 28191 70825 28249 70871
rect 28295 70825 28353 70871
rect 28399 70825 28457 70871
rect 28503 70825 28561 70871
rect 28607 70825 28665 70871
rect 28711 70825 28769 70871
rect 28815 70825 28873 70871
rect 28919 70825 28977 70871
rect 29023 70825 29081 70871
rect 29127 70825 29185 70871
rect 29231 70825 29289 70871
rect 29335 70825 29393 70871
rect 29439 70825 29497 70871
rect 29543 70825 29601 70871
rect 29647 70825 29705 70871
rect 29751 70825 29809 70871
rect 29855 70825 29913 70871
rect 29959 70825 30017 70871
rect 30063 70825 30121 70871
rect 30167 70825 30225 70871
rect 30271 70825 30329 70871
rect 30375 70825 30433 70871
rect 30479 70825 30537 70871
rect 30583 70825 30641 70871
rect 30687 70825 30745 70871
rect 30791 70825 30849 70871
rect 30895 70825 30953 70871
rect 30999 70825 31057 70871
rect 31103 70825 31161 70871
rect 31207 70825 31265 70871
rect 31311 70825 31369 70871
rect 31415 70825 31473 70871
rect 31519 70825 31577 70871
rect 31623 70825 31681 70871
rect 31727 70825 31785 70871
rect 31831 70825 31889 70871
rect 31935 70825 31993 70871
rect 32039 70825 32097 70871
rect 32143 70825 32201 70871
rect 32247 70825 32305 70871
rect 32351 70825 32409 70871
rect 32455 70825 32513 70871
rect 32559 70825 32617 70871
rect 32663 70825 32721 70871
rect 32767 70825 32825 70871
rect 32871 70825 32929 70871
rect 32975 70825 33033 70871
rect 33079 70825 33137 70871
rect 33183 70825 33241 70871
rect 33287 70825 33345 70871
rect 33391 70825 33449 70871
rect 33495 70825 33553 70871
rect 33599 70825 33657 70871
rect 33703 70825 33761 70871
rect 33807 70825 33865 70871
rect 33911 70825 33969 70871
rect 34015 70825 34073 70871
rect 34119 70825 34177 70871
rect 34223 70825 34281 70871
rect 34327 70825 34385 70871
rect 34431 70825 34489 70871
rect 34535 70825 34593 70871
rect 34639 70825 34697 70871
rect 34743 70825 34801 70871
rect 34847 70825 34905 70871
rect 34951 70825 35009 70871
rect 35055 70825 35113 70871
rect 35159 70825 35217 70871
rect 35263 70825 35321 70871
rect 35367 70825 35425 70871
rect 35471 70825 35529 70871
rect 35575 70825 35633 70871
rect 35679 70825 35737 70871
rect 35783 70825 35841 70871
rect 35887 70825 35945 70871
rect 35991 70825 36049 70871
rect 36095 70825 36153 70871
rect 36199 70825 36257 70871
rect 36303 70825 36361 70871
rect 36407 70825 36465 70871
rect 36511 70825 36569 70871
rect 36615 70825 36673 70871
rect 36719 70825 36777 70871
rect 36823 70825 36881 70871
rect 36927 70825 36985 70871
rect 37031 70825 37089 70871
rect 37135 70825 37193 70871
rect 37239 70825 37297 70871
rect 37343 70825 37401 70871
rect 37447 70825 37505 70871
rect 37551 70825 37609 70871
rect 37655 70825 37713 70871
rect 37759 70825 37817 70871
rect 37863 70825 37921 70871
rect 37967 70825 38025 70871
rect 38071 70825 38129 70871
rect 38175 70825 38233 70871
rect 38279 70825 38337 70871
rect 38383 70825 38441 70871
rect 38487 70825 38545 70871
rect 38591 70825 38649 70871
rect 38695 70825 38753 70871
rect 38799 70825 38857 70871
rect 38903 70825 38961 70871
rect 39007 70825 39065 70871
rect 39111 70825 39169 70871
rect 39215 70825 39273 70871
rect 39319 70825 39377 70871
rect 39423 70825 39481 70871
rect 39527 70825 39585 70871
rect 39631 70825 39689 70871
rect 39735 70825 39793 70871
rect 39839 70825 39897 70871
rect 39943 70825 40001 70871
rect 40047 70825 40105 70871
rect 40151 70825 40209 70871
rect 40255 70825 40313 70871
rect 40359 70825 40417 70871
rect 40463 70825 40521 70871
rect 40567 70825 40625 70871
rect 40671 70825 40729 70871
rect 40775 70825 40833 70871
rect 40879 70825 40937 70871
rect 40983 70825 41041 70871
rect 41087 70825 41145 70871
rect 41191 70825 41249 70871
rect 41295 70825 41353 70871
rect 41399 70825 41457 70871
rect 41503 70825 41561 70871
rect 41607 70825 41665 70871
rect 41711 70825 41769 70871
rect 41815 70825 41873 70871
rect 41919 70825 41977 70871
rect 42023 70825 42081 70871
rect 42127 70825 42185 70871
rect 42231 70825 42289 70871
rect 42335 70825 42393 70871
rect 42439 70825 42497 70871
rect 42543 70825 42601 70871
rect 42647 70825 42705 70871
rect 42751 70825 42809 70871
rect 42855 70825 42913 70871
rect 42959 70825 43017 70871
rect 43063 70825 43121 70871
rect 43167 70825 43225 70871
rect 43271 70825 43329 70871
rect 43375 70825 43433 70871
rect 43479 70825 43537 70871
rect 43583 70825 43641 70871
rect 43687 70825 43745 70871
rect 43791 70825 43849 70871
rect 43895 70825 43953 70871
rect 43999 70825 44057 70871
rect 44103 70825 44161 70871
rect 44207 70825 44265 70871
rect 44311 70825 44369 70871
rect 44415 70825 44473 70871
rect 44519 70825 44577 70871
rect 44623 70825 44681 70871
rect 44727 70825 44785 70871
rect 44831 70825 44889 70871
rect 44935 70825 44993 70871
rect 45039 70825 45097 70871
rect 45143 70825 45201 70871
rect 45247 70825 45305 70871
rect 45351 70825 45409 70871
rect 45455 70825 45513 70871
rect 45559 70825 45617 70871
rect 45663 70825 45721 70871
rect 45767 70825 45825 70871
rect 45871 70825 45929 70871
rect 45975 70825 46033 70871
rect 46079 70825 46137 70871
rect 46183 70825 46241 70871
rect 46287 70825 46345 70871
rect 46391 70825 46449 70871
rect 46495 70825 46553 70871
rect 46599 70825 46657 70871
rect 46703 70825 46761 70871
rect 46807 70825 46865 70871
rect 46911 70825 46969 70871
rect 47015 70825 47073 70871
rect 47119 70825 47177 70871
rect 47223 70825 47281 70871
rect 47327 70825 47385 70871
rect 47431 70825 47489 70871
rect 47535 70825 47593 70871
rect 47639 70825 47697 70871
rect 47743 70825 47801 70871
rect 47847 70825 47905 70871
rect 47951 70825 48009 70871
rect 48055 70825 48113 70871
rect 48159 70825 48217 70871
rect 48263 70825 48321 70871
rect 48367 70825 48425 70871
rect 48471 70825 48529 70871
rect 48575 70825 48633 70871
rect 48679 70825 48737 70871
rect 48783 70825 48841 70871
rect 48887 70825 48945 70871
rect 48991 70825 49049 70871
rect 49095 70825 49153 70871
rect 49199 70825 49257 70871
rect 49303 70825 49361 70871
rect 49407 70825 49465 70871
rect 49511 70825 49569 70871
rect 49615 70825 49673 70871
rect 49719 70825 49777 70871
rect 49823 70825 49881 70871
rect 49927 70825 49985 70871
rect 50031 70825 50089 70871
rect 50135 70825 50193 70871
rect 50239 70825 50297 70871
rect 50343 70825 50401 70871
rect 50447 70825 50505 70871
rect 50551 70825 50609 70871
rect 50655 70825 50713 70871
rect 50759 70825 50817 70871
rect 50863 70825 50921 70871
rect 50967 70825 51025 70871
rect 51071 70825 51129 70871
rect 51175 70825 51233 70871
rect 51279 70825 51337 70871
rect 51383 70825 51441 70871
rect 51487 70825 51545 70871
rect 51591 70825 51649 70871
rect 51695 70825 51753 70871
rect 51799 70825 51857 70871
rect 51903 70825 51961 70871
rect 52007 70825 52065 70871
rect 52111 70825 52169 70871
rect 52215 70825 52273 70871
rect 52319 70825 52377 70871
rect 52423 70825 52481 70871
rect 52527 70825 52585 70871
rect 52631 70825 52689 70871
rect 52735 70825 52793 70871
rect 52839 70825 52897 70871
rect 52943 70825 53001 70871
rect 53047 70825 53105 70871
rect 53151 70825 53209 70871
rect 53255 70825 53313 70871
rect 53359 70825 53417 70871
rect 53463 70825 53521 70871
rect 53567 70825 53625 70871
rect 53671 70825 53729 70871
rect 53775 70825 53833 70871
rect 53879 70825 53937 70871
rect 53983 70825 54041 70871
rect 54087 70825 54145 70871
rect 54191 70825 54249 70871
rect 54295 70825 54353 70871
rect 54399 70825 54457 70871
rect 54503 70825 54561 70871
rect 54607 70825 54665 70871
rect 54711 70825 54769 70871
rect 54815 70825 54873 70871
rect 54919 70825 54977 70871
rect 55023 70825 55081 70871
rect 55127 70825 55185 70871
rect 55231 70825 55289 70871
rect 55335 70825 55393 70871
rect 55439 70825 55497 70871
rect 55543 70825 55601 70871
rect 55647 70825 55705 70871
rect 55751 70825 55809 70871
rect 55855 70825 55913 70871
rect 55959 70825 56017 70871
rect 56063 70825 56121 70871
rect 56167 70825 56225 70871
rect 56271 70825 56329 70871
rect 56375 70825 56433 70871
rect 56479 70825 56537 70871
rect 56583 70825 56641 70871
rect 56687 70825 56745 70871
rect 56791 70825 56849 70871
rect 56895 70825 56953 70871
rect 56999 70825 57057 70871
rect 57103 70825 57161 70871
rect 57207 70825 57265 70871
rect 57311 70825 57369 70871
rect 57415 70825 57473 70871
rect 57519 70825 57577 70871
rect 57623 70825 57681 70871
rect 57727 70825 57785 70871
rect 57831 70825 57889 70871
rect 57935 70825 57993 70871
rect 58039 70825 58097 70871
rect 58143 70825 58201 70871
rect 58247 70825 58305 70871
rect 58351 70825 58409 70871
rect 58455 70825 58513 70871
rect 58559 70825 58617 70871
rect 58663 70825 58721 70871
rect 58767 70825 58825 70871
rect 58871 70825 58929 70871
rect 58975 70825 59033 70871
rect 59079 70825 59137 70871
rect 59183 70825 59241 70871
rect 59287 70825 59345 70871
rect 59391 70825 59449 70871
rect 59495 70825 59553 70871
rect 59599 70825 59657 70871
rect 59703 70825 59761 70871
rect 59807 70825 59865 70871
rect 59911 70825 59969 70871
rect 60015 70825 60073 70871
rect 60119 70825 60177 70871
rect 60223 70825 60281 70871
rect 60327 70825 60385 70871
rect 60431 70825 60489 70871
rect 60535 70825 60593 70871
rect 60639 70825 60697 70871
rect 60743 70825 60801 70871
rect 60847 70825 60905 70871
rect 60951 70825 61009 70871
rect 61055 70825 61113 70871
rect 61159 70825 61217 70871
rect 61263 70825 61321 70871
rect 61367 70825 61425 70871
rect 61471 70825 61529 70871
rect 61575 70825 61633 70871
rect 61679 70825 61737 70871
rect 61783 70825 61841 70871
rect 61887 70825 61945 70871
rect 61991 70825 62049 70871
rect 62095 70825 62153 70871
rect 62199 70825 62257 70871
rect 62303 70825 62361 70871
rect 62407 70825 62465 70871
rect 62511 70825 62569 70871
rect 62615 70825 62673 70871
rect 62719 70825 62777 70871
rect 62823 70825 62881 70871
rect 62927 70825 62985 70871
rect 63031 70825 63089 70871
rect 63135 70825 63193 70871
rect 63239 70825 63297 70871
rect 63343 70825 63401 70871
rect 63447 70825 63505 70871
rect 63551 70825 63609 70871
rect 63655 70825 63713 70871
rect 63759 70825 63817 70871
rect 63863 70825 63921 70871
rect 63967 70825 64025 70871
rect 64071 70825 64129 70871
rect 64175 70825 64233 70871
rect 64279 70825 64337 70871
rect 64383 70825 64441 70871
rect 64487 70825 64545 70871
rect 64591 70825 64649 70871
rect 64695 70825 64753 70871
rect 64799 70825 64857 70871
rect 64903 70825 64961 70871
rect 65007 70825 65065 70871
rect 65111 70825 65169 70871
rect 65215 70825 65273 70871
rect 65319 70825 65377 70871
rect 65423 70825 65481 70871
rect 65527 70825 65585 70871
rect 65631 70825 65689 70871
rect 65735 70825 65793 70871
rect 65839 70825 65897 70871
rect 65943 70825 66001 70871
rect 66047 70825 66105 70871
rect 66151 70825 66209 70871
rect 66255 70825 66313 70871
rect 66359 70825 66417 70871
rect 66463 70825 66521 70871
rect 66567 70825 66625 70871
rect 66671 70825 66729 70871
rect 66775 70825 66833 70871
rect 66879 70825 66937 70871
rect 66983 70825 67041 70871
rect 67087 70825 67145 70871
rect 67191 70825 67249 70871
rect 67295 70825 67353 70871
rect 67399 70825 67457 70871
rect 67503 70825 67561 70871
rect 67607 70825 67665 70871
rect 67711 70825 67769 70871
rect 67815 70825 67873 70871
rect 67919 70825 67977 70871
rect 68023 70825 68081 70871
rect 68127 70825 68185 70871
rect 68231 70825 68289 70871
rect 68335 70825 68393 70871
rect 68439 70825 68497 70871
rect 68543 70825 68601 70871
rect 68647 70825 68705 70871
rect 68751 70825 68809 70871
rect 68855 70825 68913 70871
rect 68959 70825 69017 70871
rect 69063 70825 69121 70871
rect 69167 70825 69225 70871
rect 69271 70825 69329 70871
rect 69375 70825 69433 70871
rect 69479 70825 69537 70871
rect 69583 70825 69641 70871
rect 69687 70825 69745 70871
rect 69791 70825 69849 70871
rect 69895 70825 69968 70871
rect 13097 70803 69968 70825
rect 13097 70767 13291 70803
rect 13097 70721 13119 70767
rect 13165 70721 13223 70767
rect 13269 70721 13291 70767
rect 13097 70663 13291 70721
rect 13097 70617 13119 70663
rect 13165 70617 13223 70663
rect 13269 70617 13291 70663
rect 13097 70559 13291 70617
rect 13097 70513 13119 70559
rect 13165 70513 13223 70559
rect 13269 70513 13291 70559
rect 13097 70455 13291 70513
rect 13097 70409 13119 70455
rect 13165 70409 13223 70455
rect 13269 70409 13291 70455
rect 13097 70351 13291 70409
rect 13097 70305 13119 70351
rect 13165 70305 13223 70351
rect 13269 70305 13291 70351
rect 13097 70247 13291 70305
rect 13097 70201 13119 70247
rect 13165 70201 13223 70247
rect 13269 70201 13291 70247
rect 13097 70143 13291 70201
rect 13097 70097 13119 70143
rect 13165 70097 13223 70143
rect 13269 70097 13291 70143
rect 13097 70039 13291 70097
rect 13097 69993 13119 70039
rect 13165 69993 13223 70039
rect 13269 69993 13291 70039
rect 13097 69935 13291 69993
rect 13097 69889 13119 69935
rect 13165 69889 13223 69935
rect 13269 69889 13291 69935
rect 13097 69831 13291 69889
rect 13097 69785 13119 69831
rect 13165 69785 13223 69831
rect 13269 69785 13291 69831
rect 13097 69727 13291 69785
rect 69774 70720 69968 70803
rect 69774 70674 69796 70720
rect 69842 70674 69900 70720
rect 69946 70674 69968 70720
rect 69774 70616 69968 70674
rect 69774 70570 69796 70616
rect 69842 70570 69900 70616
rect 69946 70570 69968 70616
rect 69774 70512 69968 70570
rect 69774 70466 69796 70512
rect 69842 70466 69900 70512
rect 69946 70466 69968 70512
rect 69774 70408 69968 70466
rect 69774 70362 69796 70408
rect 69842 70362 69900 70408
rect 69946 70362 69968 70408
rect 69774 70304 69968 70362
rect 69774 70258 69796 70304
rect 69842 70258 69900 70304
rect 69946 70258 69968 70304
rect 69774 70200 69968 70258
rect 69774 70154 69796 70200
rect 69842 70154 69900 70200
rect 69946 70154 69968 70200
rect 69774 70096 69968 70154
rect 69774 70050 69796 70096
rect 69842 70050 69900 70096
rect 69946 70050 69968 70096
rect 69774 69968 69968 70050
rect 69774 69946 71000 69968
rect 69774 69900 69796 69946
rect 69842 69900 69900 69946
rect 69946 69900 70004 69946
rect 70050 69900 70108 69946
rect 70154 69900 70212 69946
rect 70258 69900 70316 69946
rect 70362 69900 70420 69946
rect 70466 69900 70524 69946
rect 70570 69900 70628 69946
rect 70674 69908 71000 69946
rect 70674 69900 70824 69908
rect 69774 69862 70824 69900
rect 70870 69862 70928 69908
rect 70974 69862 71000 69908
rect 69774 69842 71000 69862
rect 69774 69796 69796 69842
rect 69842 69796 69900 69842
rect 69946 69796 70004 69842
rect 70050 69796 70108 69842
rect 70154 69796 70212 69842
rect 70258 69796 70316 69842
rect 70362 69796 70420 69842
rect 70466 69796 70524 69842
rect 70570 69796 70628 69842
rect 70674 69804 71000 69842
rect 70674 69796 70824 69804
rect 69774 69774 70824 69796
rect 13097 69681 13119 69727
rect 13165 69681 13223 69727
rect 13269 69681 13291 69727
rect 13097 69623 13291 69681
rect 13097 69577 13119 69623
rect 13165 69577 13223 69623
rect 13269 69577 13291 69623
rect 13097 69519 13291 69577
rect 13097 69473 13119 69519
rect 13165 69473 13223 69519
rect 13269 69473 13291 69519
rect 13097 69415 13291 69473
rect 13097 69369 13119 69415
rect 13165 69369 13223 69415
rect 13269 69369 13291 69415
rect 13097 69311 13291 69369
rect 13097 69265 13119 69311
rect 13165 69265 13223 69311
rect 13269 69265 13291 69311
rect 13097 69207 13291 69265
rect 13097 69161 13119 69207
rect 13165 69161 13223 69207
rect 13269 69161 13291 69207
rect 13097 69103 13291 69161
rect 13097 69057 13119 69103
rect 13165 69057 13223 69103
rect 13269 69057 13291 69103
rect 13097 68999 13291 69057
rect 13097 68953 13119 68999
rect 13165 68953 13223 68999
rect 13269 68953 13291 68999
rect 13097 68895 13291 68953
rect 13097 68849 13119 68895
rect 13165 68849 13223 68895
rect 13269 68849 13291 68895
rect 13097 68791 13291 68849
rect 13097 68745 13119 68791
rect 13165 68745 13223 68791
rect 13269 68745 13291 68791
rect 13097 68687 13291 68745
rect 13097 68641 13119 68687
rect 13165 68641 13223 68687
rect 13269 68641 13291 68687
rect 13097 68583 13291 68641
rect 13097 68537 13119 68583
rect 13165 68537 13223 68583
rect 13269 68537 13291 68583
rect 13097 68479 13291 68537
rect 13097 68433 13119 68479
rect 13165 68433 13223 68479
rect 13269 68433 13291 68479
rect 13097 68375 13291 68433
rect 13097 68329 13119 68375
rect 13165 68329 13223 68375
rect 13269 68329 13291 68375
rect 13097 68271 13291 68329
rect 13097 68225 13119 68271
rect 13165 68225 13223 68271
rect 13269 68225 13291 68271
rect 13097 68167 13291 68225
rect 13097 68121 13119 68167
rect 13165 68121 13223 68167
rect 13269 68121 13291 68167
rect 13097 68063 13291 68121
rect 13097 68017 13119 68063
rect 13165 68017 13223 68063
rect 13269 68017 13291 68063
rect 13097 67959 13291 68017
rect 13097 67913 13119 67959
rect 13165 67913 13223 67959
rect 13269 67913 13291 67959
rect 13097 67855 13291 67913
rect 13097 67809 13119 67855
rect 13165 67809 13223 67855
rect 13269 67809 13291 67855
rect 13097 67751 13291 67809
rect 13097 67705 13119 67751
rect 13165 67705 13223 67751
rect 13269 67705 13291 67751
rect 13097 67647 13291 67705
rect 13097 67601 13119 67647
rect 13165 67601 13223 67647
rect 13269 67601 13291 67647
rect 13097 67543 13291 67601
rect 13097 67497 13119 67543
rect 13165 67497 13223 67543
rect 13269 67497 13291 67543
rect 13097 67439 13291 67497
rect 13097 67393 13119 67439
rect 13165 67393 13223 67439
rect 13269 67393 13291 67439
rect 13097 67335 13291 67393
rect 13097 67289 13119 67335
rect 13165 67289 13223 67335
rect 13269 67289 13291 67335
rect 13097 67231 13291 67289
rect 13097 67185 13119 67231
rect 13165 67185 13223 67231
rect 13269 67185 13291 67231
rect 13097 67127 13291 67185
rect 13097 67081 13119 67127
rect 13165 67081 13223 67127
rect 13269 67081 13291 67127
rect 13097 67023 13291 67081
rect 13097 66977 13119 67023
rect 13165 66977 13223 67023
rect 13269 66977 13291 67023
rect 13097 66919 13291 66977
rect 13097 66873 13119 66919
rect 13165 66873 13223 66919
rect 13269 66873 13291 66919
rect 13097 66815 13291 66873
rect 13097 66769 13119 66815
rect 13165 66769 13223 66815
rect 13269 66769 13291 66815
rect 13097 66711 13291 66769
rect 13097 66665 13119 66711
rect 13165 66665 13223 66711
rect 13269 66665 13291 66711
rect 13097 66607 13291 66665
rect 13097 66561 13119 66607
rect 13165 66561 13223 66607
rect 13269 66561 13291 66607
rect 13097 66503 13291 66561
rect 13097 66457 13119 66503
rect 13165 66457 13223 66503
rect 13269 66457 13291 66503
rect 13097 66399 13291 66457
rect 13097 66353 13119 66399
rect 13165 66353 13223 66399
rect 13269 66353 13291 66399
rect 13097 66295 13291 66353
rect 13097 66249 13119 66295
rect 13165 66249 13223 66295
rect 13269 66249 13291 66295
rect 13097 66191 13291 66249
rect 13097 66145 13119 66191
rect 13165 66145 13223 66191
rect 13269 66145 13291 66191
rect 13097 66087 13291 66145
rect 13097 66041 13119 66087
rect 13165 66041 13223 66087
rect 13269 66041 13291 66087
rect 13097 65983 13291 66041
rect 13097 65937 13119 65983
rect 13165 65937 13223 65983
rect 13269 65937 13291 65983
rect 13097 65879 13291 65937
rect 13097 65833 13119 65879
rect 13165 65833 13223 65879
rect 13269 65833 13291 65879
rect 13097 65775 13291 65833
rect 13097 65729 13119 65775
rect 13165 65729 13223 65775
rect 13269 65729 13291 65775
rect 13097 65671 13291 65729
rect 13097 65625 13119 65671
rect 13165 65625 13223 65671
rect 13269 65625 13291 65671
rect 13097 65567 13291 65625
rect 13097 65521 13119 65567
rect 13165 65521 13223 65567
rect 13269 65521 13291 65567
rect 13097 65463 13291 65521
rect 13097 65417 13119 65463
rect 13165 65417 13223 65463
rect 13269 65417 13291 65463
rect 13097 65359 13291 65417
rect 13097 65313 13119 65359
rect 13165 65313 13223 65359
rect 13269 65313 13291 65359
rect 13097 65255 13291 65313
rect 13097 65209 13119 65255
rect 13165 65209 13223 65255
rect 13269 65209 13291 65255
rect 13097 65151 13291 65209
rect 13097 65105 13119 65151
rect 13165 65105 13223 65151
rect 13269 65105 13291 65151
rect 13097 65047 13291 65105
rect 13097 65001 13119 65047
rect 13165 65001 13223 65047
rect 13269 65001 13291 65047
rect 13097 64943 13291 65001
rect 13097 64897 13119 64943
rect 13165 64897 13223 64943
rect 13269 64897 13291 64943
rect 13097 64839 13291 64897
rect 13097 64793 13119 64839
rect 13165 64793 13223 64839
rect 13269 64793 13291 64839
rect 13097 64735 13291 64793
rect 13097 64689 13119 64735
rect 13165 64689 13223 64735
rect 13269 64689 13291 64735
rect 13097 64631 13291 64689
rect 13097 64585 13119 64631
rect 13165 64585 13223 64631
rect 13269 64585 13291 64631
rect 13097 64527 13291 64585
rect 13097 64481 13119 64527
rect 13165 64481 13223 64527
rect 13269 64481 13291 64527
rect 13097 64423 13291 64481
rect 13097 64377 13119 64423
rect 13165 64377 13223 64423
rect 13269 64377 13291 64423
rect 13097 64319 13291 64377
rect 13097 64273 13119 64319
rect 13165 64273 13223 64319
rect 13269 64273 13291 64319
rect 13097 64215 13291 64273
rect 13097 64169 13119 64215
rect 13165 64169 13223 64215
rect 13269 64169 13291 64215
rect 13097 64111 13291 64169
rect 13097 64065 13119 64111
rect 13165 64065 13223 64111
rect 13269 64065 13291 64111
rect 13097 64007 13291 64065
rect 13097 63961 13119 64007
rect 13165 63961 13223 64007
rect 13269 63961 13291 64007
rect 13097 63903 13291 63961
rect 13097 63857 13119 63903
rect 13165 63857 13223 63903
rect 13269 63857 13291 63903
rect 13097 63799 13291 63857
rect 13097 63753 13119 63799
rect 13165 63753 13223 63799
rect 13269 63753 13291 63799
rect 13097 63695 13291 63753
rect 13097 63649 13119 63695
rect 13165 63649 13223 63695
rect 13269 63649 13291 63695
rect 13097 63591 13291 63649
rect 13097 63545 13119 63591
rect 13165 63545 13223 63591
rect 13269 63545 13291 63591
rect 13097 63487 13291 63545
rect 13097 63441 13119 63487
rect 13165 63441 13223 63487
rect 13269 63441 13291 63487
rect 13097 63383 13291 63441
rect 13097 63337 13119 63383
rect 13165 63337 13223 63383
rect 13269 63337 13291 63383
rect 13097 63279 13291 63337
rect 13097 63233 13119 63279
rect 13165 63233 13223 63279
rect 13269 63233 13291 63279
rect 13097 63175 13291 63233
rect 13097 63129 13119 63175
rect 13165 63129 13223 63175
rect 13269 63129 13291 63175
rect 13097 63071 13291 63129
rect 13097 63025 13119 63071
rect 13165 63025 13223 63071
rect 13269 63025 13291 63071
rect 13097 62967 13291 63025
rect 13097 62921 13119 62967
rect 13165 62921 13223 62967
rect 13269 62921 13291 62967
rect 13097 62863 13291 62921
rect 13097 62817 13119 62863
rect 13165 62817 13223 62863
rect 13269 62817 13291 62863
rect 13097 62759 13291 62817
rect 13097 62713 13119 62759
rect 13165 62713 13223 62759
rect 13269 62713 13291 62759
rect 13097 62655 13291 62713
rect 13097 62609 13119 62655
rect 13165 62609 13223 62655
rect 13269 62609 13291 62655
rect 13097 62551 13291 62609
rect 13097 62505 13119 62551
rect 13165 62505 13223 62551
rect 13269 62505 13291 62551
rect 13097 62447 13291 62505
rect 13097 62401 13119 62447
rect 13165 62401 13223 62447
rect 13269 62401 13291 62447
rect 13097 62343 13291 62401
rect 13097 62297 13119 62343
rect 13165 62297 13223 62343
rect 13269 62297 13291 62343
rect 13097 62239 13291 62297
rect 13097 62193 13119 62239
rect 13165 62193 13223 62239
rect 13269 62193 13291 62239
rect 13097 62135 13291 62193
rect 13097 62089 13119 62135
rect 13165 62089 13223 62135
rect 13269 62089 13291 62135
rect 13097 62031 13291 62089
rect 13097 61985 13119 62031
rect 13165 61985 13223 62031
rect 13269 61985 13291 62031
rect 13097 61927 13291 61985
rect 13097 61881 13119 61927
rect 13165 61881 13223 61927
rect 13269 61881 13291 61927
rect 13097 61823 13291 61881
rect 13097 61777 13119 61823
rect 13165 61777 13223 61823
rect 13269 61777 13291 61823
rect 13097 61719 13291 61777
rect 13097 61673 13119 61719
rect 13165 61673 13223 61719
rect 13269 61673 13291 61719
rect 13097 61615 13291 61673
rect 13097 61569 13119 61615
rect 13165 61569 13223 61615
rect 13269 61569 13291 61615
rect 13097 61511 13291 61569
rect 13097 61465 13119 61511
rect 13165 61465 13223 61511
rect 13269 61465 13291 61511
rect 13097 61407 13291 61465
rect 13097 61361 13119 61407
rect 13165 61361 13223 61407
rect 13269 61361 13291 61407
rect 13097 61303 13291 61361
rect 13097 61257 13119 61303
rect 13165 61257 13223 61303
rect 13269 61257 13291 61303
rect 13097 61199 13291 61257
rect 13097 61153 13119 61199
rect 13165 61153 13223 61199
rect 13269 61153 13291 61199
rect 13097 61095 13291 61153
rect 13097 61049 13119 61095
rect 13165 61049 13223 61095
rect 13269 61049 13291 61095
rect 13097 60991 13291 61049
rect 13097 60945 13119 60991
rect 13165 60945 13223 60991
rect 13269 60945 13291 60991
rect 13097 60887 13291 60945
rect 13097 60841 13119 60887
rect 13165 60841 13223 60887
rect 13269 60841 13291 60887
rect 13097 60783 13291 60841
rect 13097 60737 13119 60783
rect 13165 60737 13223 60783
rect 13269 60737 13291 60783
rect 13097 60679 13291 60737
rect 13097 60633 13119 60679
rect 13165 60633 13223 60679
rect 13269 60633 13291 60679
rect 13097 60575 13291 60633
rect 13097 60529 13119 60575
rect 13165 60529 13223 60575
rect 13269 60529 13291 60575
rect 13097 60471 13291 60529
rect 13097 60425 13119 60471
rect 13165 60425 13223 60471
rect 13269 60425 13291 60471
rect 13097 60367 13291 60425
rect 13097 60321 13119 60367
rect 13165 60321 13223 60367
rect 13269 60321 13291 60367
rect 13097 60263 13291 60321
rect 13097 60217 13119 60263
rect 13165 60217 13223 60263
rect 13269 60217 13291 60263
rect 13097 60159 13291 60217
rect 13097 60113 13119 60159
rect 13165 60113 13223 60159
rect 13269 60113 13291 60159
rect 13097 60055 13291 60113
rect 13097 60009 13119 60055
rect 13165 60009 13223 60055
rect 13269 60009 13291 60055
rect 13097 59951 13291 60009
rect 13097 59905 13119 59951
rect 13165 59905 13223 59951
rect 13269 59905 13291 59951
rect 13097 59847 13291 59905
rect 13097 59801 13119 59847
rect 13165 59801 13223 59847
rect 13269 59801 13291 59847
rect 13097 59743 13291 59801
rect 13097 59697 13119 59743
rect 13165 59697 13223 59743
rect 13269 59697 13291 59743
rect 13097 59639 13291 59697
rect 13097 59593 13119 59639
rect 13165 59593 13223 59639
rect 13269 59593 13291 59639
rect 13097 59535 13291 59593
rect 13097 59489 13119 59535
rect 13165 59489 13223 59535
rect 13269 59489 13291 59535
rect 13097 59431 13291 59489
rect 13097 59385 13119 59431
rect 13165 59385 13223 59431
rect 13269 59385 13291 59431
rect 13097 59327 13291 59385
rect 13097 59281 13119 59327
rect 13165 59281 13223 59327
rect 13269 59281 13291 59327
rect 13097 59223 13291 59281
rect 13097 59177 13119 59223
rect 13165 59177 13223 59223
rect 13269 59177 13291 59223
rect 13097 59119 13291 59177
rect 13097 59073 13119 59119
rect 13165 59073 13223 59119
rect 13269 59073 13291 59119
rect 13097 59015 13291 59073
rect 13097 58969 13119 59015
rect 13165 58969 13223 59015
rect 13269 58969 13291 59015
rect 13097 58911 13291 58969
rect 13097 58865 13119 58911
rect 13165 58865 13223 58911
rect 13269 58865 13291 58911
rect 13097 58807 13291 58865
rect 13097 58761 13119 58807
rect 13165 58761 13223 58807
rect 13269 58761 13291 58807
rect 13097 58703 13291 58761
rect 13097 58657 13119 58703
rect 13165 58657 13223 58703
rect 13269 58657 13291 58703
rect 13097 58599 13291 58657
rect 13097 58553 13119 58599
rect 13165 58553 13223 58599
rect 13269 58553 13291 58599
rect 13097 58495 13291 58553
rect 13097 58449 13119 58495
rect 13165 58449 13223 58495
rect 13269 58449 13291 58495
rect 13097 58391 13291 58449
rect 13097 58345 13119 58391
rect 13165 58345 13223 58391
rect 13269 58345 13291 58391
rect 13097 58287 13291 58345
rect 13097 58241 13119 58287
rect 13165 58241 13223 58287
rect 13269 58241 13291 58287
rect 13097 58183 13291 58241
rect 13097 58137 13119 58183
rect 13165 58137 13223 58183
rect 13269 58137 13291 58183
rect 13097 58079 13291 58137
rect 13097 58033 13119 58079
rect 13165 58033 13223 58079
rect 13269 58033 13291 58079
rect 13097 57975 13291 58033
rect 13097 57929 13119 57975
rect 13165 57929 13223 57975
rect 13269 57929 13291 57975
rect 13097 57871 13291 57929
rect 13097 57825 13119 57871
rect 13165 57825 13223 57871
rect 13269 57825 13291 57871
rect 13097 57767 13291 57825
rect 13097 57721 13119 57767
rect 13165 57721 13223 57767
rect 13269 57721 13291 57767
rect 13097 57663 13291 57721
rect 13097 57617 13119 57663
rect 13165 57617 13223 57663
rect 13269 57617 13291 57663
rect 13097 57559 13291 57617
rect 13097 57513 13119 57559
rect 13165 57513 13223 57559
rect 13269 57513 13291 57559
rect 13097 57455 13291 57513
rect 13097 57409 13119 57455
rect 13165 57409 13223 57455
rect 13269 57409 13291 57455
rect 13097 57351 13291 57409
rect 13097 57305 13119 57351
rect 13165 57305 13223 57351
rect 13269 57305 13291 57351
rect 13097 57247 13291 57305
rect 13097 57201 13119 57247
rect 13165 57201 13223 57247
rect 13269 57201 13291 57247
rect 13097 57143 13291 57201
rect 13097 57097 13119 57143
rect 13165 57097 13223 57143
rect 13269 57097 13291 57143
rect 13097 57039 13291 57097
rect 13097 56993 13119 57039
rect 13165 56993 13223 57039
rect 13269 56993 13291 57039
rect 13097 56935 13291 56993
rect 13097 56889 13119 56935
rect 13165 56889 13223 56935
rect 13269 56889 13291 56935
rect 13097 56831 13291 56889
rect 13097 56785 13119 56831
rect 13165 56785 13223 56831
rect 13269 56785 13291 56831
rect 13097 56727 13291 56785
rect 13097 56681 13119 56727
rect 13165 56681 13223 56727
rect 13269 56681 13291 56727
rect 13097 56623 13291 56681
rect 13097 56577 13119 56623
rect 13165 56577 13223 56623
rect 13269 56577 13291 56623
rect 13097 56519 13291 56577
rect 13097 56473 13119 56519
rect 13165 56473 13223 56519
rect 13269 56473 13291 56519
rect 13097 56415 13291 56473
rect 13097 56369 13119 56415
rect 13165 56369 13223 56415
rect 13269 56369 13291 56415
rect 13097 56311 13291 56369
rect 13097 56265 13119 56311
rect 13165 56265 13223 56311
rect 13269 56265 13291 56311
rect 13097 56207 13291 56265
rect 13097 56161 13119 56207
rect 13165 56161 13223 56207
rect 13269 56161 13291 56207
rect 13097 56103 13291 56161
rect 13097 56057 13119 56103
rect 13165 56057 13223 56103
rect 13269 56057 13291 56103
rect 13097 55999 13291 56057
rect 13097 55953 13119 55999
rect 13165 55953 13223 55999
rect 13269 55953 13291 55999
rect 13097 55895 13291 55953
rect 13097 55849 13119 55895
rect 13165 55849 13223 55895
rect 13269 55849 13291 55895
rect 13097 55791 13291 55849
rect 13097 55745 13119 55791
rect 13165 55745 13223 55791
rect 13269 55745 13291 55791
rect 13097 55687 13291 55745
rect 13097 55641 13119 55687
rect 13165 55641 13223 55687
rect 13269 55641 13291 55687
rect 13097 55583 13291 55641
rect 13097 55537 13119 55583
rect 13165 55537 13223 55583
rect 13269 55537 13291 55583
rect 13097 55479 13291 55537
rect 13097 55433 13119 55479
rect 13165 55433 13223 55479
rect 13269 55433 13291 55479
rect 13097 55375 13291 55433
rect 13097 55329 13119 55375
rect 13165 55329 13223 55375
rect 13269 55329 13291 55375
rect 13097 55271 13291 55329
rect 13097 55225 13119 55271
rect 13165 55225 13223 55271
rect 13269 55225 13291 55271
rect 13097 55167 13291 55225
rect 13097 55121 13119 55167
rect 13165 55121 13223 55167
rect 13269 55121 13291 55167
rect 13097 55063 13291 55121
rect 13097 55017 13119 55063
rect 13165 55017 13223 55063
rect 13269 55017 13291 55063
rect 13097 54959 13291 55017
rect 13097 54913 13119 54959
rect 13165 54913 13223 54959
rect 13269 54913 13291 54959
rect 13097 54855 13291 54913
rect 13097 54809 13119 54855
rect 13165 54809 13223 54855
rect 13269 54809 13291 54855
rect 13097 54751 13291 54809
rect 13097 54705 13119 54751
rect 13165 54705 13223 54751
rect 13269 54705 13291 54751
rect 13097 54647 13291 54705
rect 13097 54601 13119 54647
rect 13165 54601 13223 54647
rect 13269 54601 13291 54647
rect 13097 54543 13291 54601
rect 13097 54497 13119 54543
rect 13165 54497 13223 54543
rect 13269 54497 13291 54543
rect 13097 54439 13291 54497
rect 13097 54393 13119 54439
rect 13165 54393 13223 54439
rect 13269 54393 13291 54439
rect 13097 54335 13291 54393
rect 13097 54289 13119 54335
rect 13165 54289 13223 54335
rect 13269 54289 13291 54335
rect 13097 54231 13291 54289
rect 13097 54185 13119 54231
rect 13165 54185 13223 54231
rect 13269 54185 13291 54231
rect 13097 54127 13291 54185
rect 13097 54081 13119 54127
rect 13165 54081 13223 54127
rect 13269 54081 13291 54127
rect 13097 54023 13291 54081
rect 13097 53977 13119 54023
rect 13165 53977 13223 54023
rect 13269 53977 13291 54023
rect 13097 53919 13291 53977
rect 13097 53873 13119 53919
rect 13165 53873 13223 53919
rect 13269 53873 13291 53919
rect 13097 53815 13291 53873
rect 13097 53769 13119 53815
rect 13165 53769 13223 53815
rect 13269 53769 13291 53815
rect 13097 53711 13291 53769
rect 13097 53665 13119 53711
rect 13165 53665 13223 53711
rect 13269 53665 13291 53711
rect 13097 53607 13291 53665
rect 13097 53561 13119 53607
rect 13165 53561 13223 53607
rect 13269 53561 13291 53607
rect 13097 53503 13291 53561
rect 13097 53457 13119 53503
rect 13165 53457 13223 53503
rect 13269 53457 13291 53503
rect 13097 53399 13291 53457
rect 13097 53353 13119 53399
rect 13165 53353 13223 53399
rect 13269 53353 13291 53399
rect 13097 53295 13291 53353
rect 13097 53249 13119 53295
rect 13165 53249 13223 53295
rect 13269 53249 13291 53295
rect 13097 53191 13291 53249
rect 13097 53145 13119 53191
rect 13165 53145 13223 53191
rect 13269 53145 13291 53191
rect 13097 53087 13291 53145
rect 13097 53041 13119 53087
rect 13165 53041 13223 53087
rect 13269 53041 13291 53087
rect 13097 52983 13291 53041
rect 13097 52937 13119 52983
rect 13165 52937 13223 52983
rect 13269 52937 13291 52983
rect 13097 52879 13291 52937
rect 13097 52833 13119 52879
rect 13165 52833 13223 52879
rect 13269 52833 13291 52879
rect 13097 52775 13291 52833
rect 13097 52729 13119 52775
rect 13165 52729 13223 52775
rect 13269 52729 13291 52775
rect 13097 52671 13291 52729
rect 13097 52625 13119 52671
rect 13165 52625 13223 52671
rect 13269 52625 13291 52671
rect 13097 52567 13291 52625
rect 13097 52521 13119 52567
rect 13165 52521 13223 52567
rect 13269 52521 13291 52567
rect 13097 52463 13291 52521
rect 13097 52417 13119 52463
rect 13165 52417 13223 52463
rect 13269 52417 13291 52463
rect 13097 52359 13291 52417
rect 13097 52313 13119 52359
rect 13165 52313 13223 52359
rect 13269 52313 13291 52359
rect 13097 52255 13291 52313
rect 13097 52209 13119 52255
rect 13165 52209 13223 52255
rect 13269 52209 13291 52255
rect 13097 52151 13291 52209
rect 13097 52105 13119 52151
rect 13165 52105 13223 52151
rect 13269 52105 13291 52151
rect 13097 52047 13291 52105
rect 13097 52001 13119 52047
rect 13165 52001 13223 52047
rect 13269 52001 13291 52047
rect 13097 51943 13291 52001
rect 13097 51897 13119 51943
rect 13165 51897 13223 51943
rect 13269 51897 13291 51943
rect 13097 51839 13291 51897
rect 13097 51793 13119 51839
rect 13165 51793 13223 51839
rect 13269 51793 13291 51839
rect 13097 51735 13291 51793
rect 13097 51689 13119 51735
rect 13165 51689 13223 51735
rect 13269 51689 13291 51735
rect 13097 51631 13291 51689
rect 13097 51585 13119 51631
rect 13165 51585 13223 51631
rect 13269 51585 13291 51631
rect 13097 51527 13291 51585
rect 13097 51481 13119 51527
rect 13165 51481 13223 51527
rect 13269 51481 13291 51527
rect 13097 51423 13291 51481
rect 13097 51377 13119 51423
rect 13165 51377 13223 51423
rect 13269 51377 13291 51423
rect 13097 51319 13291 51377
rect 13097 51273 13119 51319
rect 13165 51273 13223 51319
rect 13269 51273 13291 51319
rect 13097 51215 13291 51273
rect 13097 51169 13119 51215
rect 13165 51169 13223 51215
rect 13269 51169 13291 51215
rect 13097 51111 13291 51169
rect 13097 51065 13119 51111
rect 13165 51065 13223 51111
rect 13269 51065 13291 51111
rect 13097 51007 13291 51065
rect 13097 50961 13119 51007
rect 13165 50961 13223 51007
rect 13269 50961 13291 51007
rect 13097 50903 13291 50961
rect 13097 50857 13119 50903
rect 13165 50857 13223 50903
rect 13269 50857 13291 50903
rect 13097 50799 13291 50857
rect 13097 50753 13119 50799
rect 13165 50753 13223 50799
rect 13269 50753 13291 50799
rect 13097 50695 13291 50753
rect 13097 50649 13119 50695
rect 13165 50649 13223 50695
rect 13269 50649 13291 50695
rect 13097 50591 13291 50649
rect 13097 50545 13119 50591
rect 13165 50545 13223 50591
rect 13269 50545 13291 50591
rect 13097 50487 13291 50545
rect 13097 50441 13119 50487
rect 13165 50441 13223 50487
rect 13269 50441 13291 50487
rect 13097 50383 13291 50441
rect 13097 50337 13119 50383
rect 13165 50337 13223 50383
rect 13269 50337 13291 50383
rect 13097 50279 13291 50337
rect 13097 50233 13119 50279
rect 13165 50233 13223 50279
rect 13269 50233 13291 50279
rect 13097 50175 13291 50233
rect 13097 50129 13119 50175
rect 13165 50129 13223 50175
rect 13269 50129 13291 50175
rect 13097 50071 13291 50129
rect 13097 50025 13119 50071
rect 13165 50025 13223 50071
rect 13269 50025 13291 50071
rect 13097 49967 13291 50025
rect 13097 49921 13119 49967
rect 13165 49921 13223 49967
rect 13269 49921 13291 49967
rect 13097 49863 13291 49921
rect 13097 49817 13119 49863
rect 13165 49817 13223 49863
rect 13269 49817 13291 49863
rect 13097 49759 13291 49817
rect 13097 49713 13119 49759
rect 13165 49713 13223 49759
rect 13269 49713 13291 49759
rect 13097 49655 13291 49713
rect 13097 49609 13119 49655
rect 13165 49609 13223 49655
rect 13269 49609 13291 49655
rect 13097 49551 13291 49609
rect 13097 49505 13119 49551
rect 13165 49505 13223 49551
rect 13269 49505 13291 49551
rect 13097 49447 13291 49505
rect 13097 49401 13119 49447
rect 13165 49401 13223 49447
rect 13269 49401 13291 49447
rect 13097 49343 13291 49401
rect 13097 49297 13119 49343
rect 13165 49297 13223 49343
rect 13269 49297 13291 49343
rect 13097 49239 13291 49297
rect 13097 49193 13119 49239
rect 13165 49193 13223 49239
rect 13269 49193 13291 49239
rect 13097 49135 13291 49193
rect 13097 49089 13119 49135
rect 13165 49089 13223 49135
rect 13269 49089 13291 49135
rect 13097 49031 13291 49089
rect 13097 48985 13119 49031
rect 13165 48985 13223 49031
rect 13269 48985 13291 49031
rect 13097 48927 13291 48985
rect 13097 48881 13119 48927
rect 13165 48881 13223 48927
rect 13269 48881 13291 48927
rect 13097 48823 13291 48881
rect 13097 48777 13119 48823
rect 13165 48777 13223 48823
rect 13269 48777 13291 48823
rect 13097 48719 13291 48777
rect 13097 48673 13119 48719
rect 13165 48673 13223 48719
rect 13269 48673 13291 48719
rect 13097 48615 13291 48673
rect 13097 48569 13119 48615
rect 13165 48569 13223 48615
rect 13269 48569 13291 48615
rect 13097 48511 13291 48569
rect 13097 48465 13119 48511
rect 13165 48465 13223 48511
rect 13269 48465 13291 48511
rect 13097 48407 13291 48465
rect 13097 48361 13119 48407
rect 13165 48361 13223 48407
rect 13269 48361 13291 48407
rect 13097 48303 13291 48361
rect 13097 48257 13119 48303
rect 13165 48257 13223 48303
rect 13269 48257 13291 48303
rect 13097 48199 13291 48257
rect 13097 48153 13119 48199
rect 13165 48153 13223 48199
rect 13269 48153 13291 48199
rect 13097 48095 13291 48153
rect 13097 48049 13119 48095
rect 13165 48049 13223 48095
rect 13269 48049 13291 48095
rect 13097 47991 13291 48049
rect 13097 47945 13119 47991
rect 13165 47945 13223 47991
rect 13269 47945 13291 47991
rect 13097 47887 13291 47945
rect 13097 47841 13119 47887
rect 13165 47841 13223 47887
rect 13269 47841 13291 47887
rect 13097 47783 13291 47841
rect 13097 47737 13119 47783
rect 13165 47737 13223 47783
rect 13269 47737 13291 47783
rect 13097 47679 13291 47737
rect 13097 47633 13119 47679
rect 13165 47633 13223 47679
rect 13269 47633 13291 47679
rect 13097 47575 13291 47633
rect 13097 47529 13119 47575
rect 13165 47529 13223 47575
rect 13269 47529 13291 47575
rect 13097 47471 13291 47529
rect 13097 47425 13119 47471
rect 13165 47425 13223 47471
rect 13269 47425 13291 47471
rect 13097 47367 13291 47425
rect 13097 47321 13119 47367
rect 13165 47321 13223 47367
rect 13269 47321 13291 47367
rect 13097 47263 13291 47321
rect 13097 47217 13119 47263
rect 13165 47217 13223 47263
rect 13269 47217 13291 47263
rect 13097 47159 13291 47217
rect 13097 47113 13119 47159
rect 13165 47113 13223 47159
rect 13269 47113 13291 47159
rect 13097 47055 13291 47113
rect 13097 47009 13119 47055
rect 13165 47009 13223 47055
rect 13269 47009 13291 47055
rect 13097 46951 13291 47009
rect 13097 46905 13119 46951
rect 13165 46905 13223 46951
rect 13269 46905 13291 46951
rect 13097 46847 13291 46905
rect 13097 46801 13119 46847
rect 13165 46801 13223 46847
rect 13269 46801 13291 46847
rect 13097 46743 13291 46801
rect 13097 46697 13119 46743
rect 13165 46697 13223 46743
rect 13269 46697 13291 46743
rect 13097 46639 13291 46697
rect 13097 46593 13119 46639
rect 13165 46593 13223 46639
rect 13269 46593 13291 46639
rect 13097 46535 13291 46593
rect 13097 46489 13119 46535
rect 13165 46489 13223 46535
rect 13269 46489 13291 46535
rect 13097 46431 13291 46489
rect 13097 46385 13119 46431
rect 13165 46385 13223 46431
rect 13269 46385 13291 46431
rect 13097 46327 13291 46385
rect 13097 46281 13119 46327
rect 13165 46281 13223 46327
rect 13269 46281 13291 46327
rect 13097 46223 13291 46281
rect 13097 46177 13119 46223
rect 13165 46177 13223 46223
rect 13269 46177 13291 46223
rect 13097 46119 13291 46177
rect 13097 46073 13119 46119
rect 13165 46073 13223 46119
rect 13269 46073 13291 46119
rect 13097 46015 13291 46073
rect 13097 45969 13119 46015
rect 13165 45969 13223 46015
rect 13269 45969 13291 46015
rect 13097 45911 13291 45969
rect 13097 45865 13119 45911
rect 13165 45865 13223 45911
rect 13269 45865 13291 45911
rect 13097 45807 13291 45865
rect 13097 45761 13119 45807
rect 13165 45761 13223 45807
rect 13269 45761 13291 45807
rect 13097 45703 13291 45761
rect 13097 45657 13119 45703
rect 13165 45657 13223 45703
rect 13269 45657 13291 45703
rect 13097 45599 13291 45657
rect 13097 45553 13119 45599
rect 13165 45553 13223 45599
rect 13269 45553 13291 45599
rect 13097 45495 13291 45553
rect 13097 45449 13119 45495
rect 13165 45449 13223 45495
rect 13269 45449 13291 45495
rect 13097 45391 13291 45449
rect 13097 45345 13119 45391
rect 13165 45345 13223 45391
rect 13269 45345 13291 45391
rect 13097 45287 13291 45345
rect 13097 45241 13119 45287
rect 13165 45241 13223 45287
rect 13269 45241 13291 45287
rect 13097 45183 13291 45241
rect 13097 45137 13119 45183
rect 13165 45137 13223 45183
rect 13269 45137 13291 45183
rect 13097 45079 13291 45137
rect 13097 45033 13119 45079
rect 13165 45033 13223 45079
rect 13269 45033 13291 45079
rect 13097 44843 13291 45033
rect 70802 69758 70824 69774
rect 70870 69758 70928 69804
rect 70974 69758 71000 69804
rect 70802 69700 71000 69758
rect 70802 69654 70824 69700
rect 70870 69654 70928 69700
rect 70974 69654 71000 69700
rect 70802 69596 71000 69654
rect 70802 69550 70824 69596
rect 70870 69550 70928 69596
rect 70974 69550 71000 69596
rect 70802 69492 71000 69550
rect 70802 69446 70824 69492
rect 70870 69446 70928 69492
rect 70974 69446 71000 69492
rect 70802 69388 71000 69446
rect 70802 69342 70824 69388
rect 70870 69342 70928 69388
rect 70974 69342 71000 69388
rect 70802 69284 71000 69342
rect 70802 69238 70824 69284
rect 70870 69238 70928 69284
rect 70974 69238 71000 69284
rect 70802 69180 71000 69238
rect 70802 69134 70824 69180
rect 70870 69134 70928 69180
rect 70974 69134 71000 69180
rect 70802 69076 71000 69134
rect 70802 69030 70824 69076
rect 70870 69030 70928 69076
rect 70974 69030 71000 69076
rect 70802 68972 71000 69030
rect 70802 68926 70824 68972
rect 70870 68926 70928 68972
rect 70974 68926 71000 68972
rect 70802 68868 71000 68926
rect 70802 68822 70824 68868
rect 70870 68822 70928 68868
rect 70974 68822 71000 68868
rect 70802 68764 71000 68822
rect 70802 68718 70824 68764
rect 70870 68718 70928 68764
rect 70974 68718 71000 68764
rect 70802 68660 71000 68718
rect 70802 68614 70824 68660
rect 70870 68614 70928 68660
rect 70974 68614 71000 68660
rect 70802 68556 71000 68614
rect 70802 68510 70824 68556
rect 70870 68510 70928 68556
rect 70974 68510 71000 68556
rect 70802 68452 71000 68510
rect 70802 68406 70824 68452
rect 70870 68406 70928 68452
rect 70974 68406 71000 68452
rect 70802 68348 71000 68406
rect 70802 68302 70824 68348
rect 70870 68302 70928 68348
rect 70974 68302 71000 68348
rect 70802 68244 71000 68302
rect 70802 68198 70824 68244
rect 70870 68198 70928 68244
rect 70974 68198 71000 68244
rect 70802 68140 71000 68198
rect 70802 68094 70824 68140
rect 70870 68094 70928 68140
rect 70974 68094 71000 68140
rect 70802 68036 71000 68094
rect 70802 67990 70824 68036
rect 70870 67990 70928 68036
rect 70974 67990 71000 68036
rect 70802 67932 71000 67990
rect 70802 67886 70824 67932
rect 70870 67886 70928 67932
rect 70974 67886 71000 67932
rect 70802 67828 71000 67886
rect 70802 67782 70824 67828
rect 70870 67782 70928 67828
rect 70974 67782 71000 67828
rect 70802 67724 71000 67782
rect 70802 67678 70824 67724
rect 70870 67678 70928 67724
rect 70974 67678 71000 67724
rect 70802 67620 71000 67678
rect 70802 67574 70824 67620
rect 70870 67574 70928 67620
rect 70974 67574 71000 67620
rect 70802 67516 71000 67574
rect 70802 67470 70824 67516
rect 70870 67470 70928 67516
rect 70974 67470 71000 67516
rect 70802 67412 71000 67470
rect 70802 67366 70824 67412
rect 70870 67366 70928 67412
rect 70974 67366 71000 67412
rect 70802 67308 71000 67366
rect 70802 67262 70824 67308
rect 70870 67262 70928 67308
rect 70974 67262 71000 67308
rect 70802 67204 71000 67262
rect 70802 67158 70824 67204
rect 70870 67158 70928 67204
rect 70974 67158 71000 67204
rect 70802 67100 71000 67158
rect 70802 67054 70824 67100
rect 70870 67054 70928 67100
rect 70974 67054 71000 67100
rect 70802 66996 71000 67054
rect 70802 66950 70824 66996
rect 70870 66950 70928 66996
rect 70974 66950 71000 66996
rect 70802 66892 71000 66950
rect 70802 66846 70824 66892
rect 70870 66846 70928 66892
rect 70974 66846 71000 66892
rect 70802 66788 71000 66846
rect 70802 66742 70824 66788
rect 70870 66742 70928 66788
rect 70974 66742 71000 66788
rect 70802 66684 71000 66742
rect 70802 66638 70824 66684
rect 70870 66638 70928 66684
rect 70974 66638 71000 66684
rect 70802 66580 71000 66638
rect 70802 66534 70824 66580
rect 70870 66534 70928 66580
rect 70974 66534 71000 66580
rect 70802 66476 71000 66534
rect 70802 66430 70824 66476
rect 70870 66430 70928 66476
rect 70974 66430 71000 66476
rect 70802 66372 71000 66430
rect 70802 66326 70824 66372
rect 70870 66326 70928 66372
rect 70974 66326 71000 66372
rect 70802 66268 71000 66326
rect 70802 66222 70824 66268
rect 70870 66222 70928 66268
rect 70974 66222 71000 66268
rect 70802 66164 71000 66222
rect 70802 66118 70824 66164
rect 70870 66118 70928 66164
rect 70974 66118 71000 66164
rect 70802 66060 71000 66118
rect 70802 66014 70824 66060
rect 70870 66014 70928 66060
rect 70974 66014 71000 66060
rect 70802 65956 71000 66014
rect 70802 65910 70824 65956
rect 70870 65910 70928 65956
rect 70974 65910 71000 65956
rect 70802 65852 71000 65910
rect 70802 65806 70824 65852
rect 70870 65806 70928 65852
rect 70974 65806 71000 65852
rect 70802 65748 71000 65806
rect 70802 65702 70824 65748
rect 70870 65702 70928 65748
rect 70974 65702 71000 65748
rect 70802 65644 71000 65702
rect 70802 65598 70824 65644
rect 70870 65598 70928 65644
rect 70974 65598 71000 65644
rect 70802 65540 71000 65598
rect 70802 65494 70824 65540
rect 70870 65494 70928 65540
rect 70974 65494 71000 65540
rect 70802 65436 71000 65494
rect 70802 65390 70824 65436
rect 70870 65390 70928 65436
rect 70974 65390 71000 65436
rect 70802 65332 71000 65390
rect 70802 65286 70824 65332
rect 70870 65286 70928 65332
rect 70974 65286 71000 65332
rect 70802 65228 71000 65286
rect 70802 65182 70824 65228
rect 70870 65182 70928 65228
rect 70974 65182 71000 65228
rect 70802 65124 71000 65182
rect 70802 65078 70824 65124
rect 70870 65078 70928 65124
rect 70974 65078 71000 65124
rect 70802 65020 71000 65078
rect 70802 64974 70824 65020
rect 70870 64974 70928 65020
rect 70974 64974 71000 65020
rect 70802 64916 71000 64974
rect 70802 64870 70824 64916
rect 70870 64870 70928 64916
rect 70974 64870 71000 64916
rect 70802 64812 71000 64870
rect 70802 64766 70824 64812
rect 70870 64766 70928 64812
rect 70974 64766 71000 64812
rect 70802 64708 71000 64766
rect 70802 64662 70824 64708
rect 70870 64662 70928 64708
rect 70974 64662 71000 64708
rect 70802 64604 71000 64662
rect 70802 64558 70824 64604
rect 70870 64558 70928 64604
rect 70974 64558 71000 64604
rect 70802 64500 71000 64558
rect 70802 64454 70824 64500
rect 70870 64454 70928 64500
rect 70974 64454 71000 64500
rect 70802 64396 71000 64454
rect 70802 64350 70824 64396
rect 70870 64350 70928 64396
rect 70974 64350 71000 64396
rect 70802 64292 71000 64350
rect 70802 64246 70824 64292
rect 70870 64246 70928 64292
rect 70974 64246 71000 64292
rect 70802 64188 71000 64246
rect 70802 64142 70824 64188
rect 70870 64142 70928 64188
rect 70974 64142 71000 64188
rect 70802 64084 71000 64142
rect 70802 64038 70824 64084
rect 70870 64038 70928 64084
rect 70974 64038 71000 64084
rect 70802 63980 71000 64038
rect 70802 63934 70824 63980
rect 70870 63934 70928 63980
rect 70974 63934 71000 63980
rect 70802 63876 71000 63934
rect 70802 63830 70824 63876
rect 70870 63830 70928 63876
rect 70974 63830 71000 63876
rect 70802 63772 71000 63830
rect 70802 63726 70824 63772
rect 70870 63726 70928 63772
rect 70974 63726 71000 63772
rect 70802 63668 71000 63726
rect 70802 63622 70824 63668
rect 70870 63622 70928 63668
rect 70974 63622 71000 63668
rect 70802 63564 71000 63622
rect 70802 63518 70824 63564
rect 70870 63518 70928 63564
rect 70974 63518 71000 63564
rect 70802 63460 71000 63518
rect 70802 63414 70824 63460
rect 70870 63414 70928 63460
rect 70974 63414 71000 63460
rect 70802 63356 71000 63414
rect 70802 63310 70824 63356
rect 70870 63310 70928 63356
rect 70974 63310 71000 63356
rect 70802 63252 71000 63310
rect 70802 63206 70824 63252
rect 70870 63206 70928 63252
rect 70974 63206 71000 63252
rect 70802 63148 71000 63206
rect 70802 63102 70824 63148
rect 70870 63102 70928 63148
rect 70974 63102 71000 63148
rect 70802 63044 71000 63102
rect 70802 62998 70824 63044
rect 70870 62998 70928 63044
rect 70974 62998 71000 63044
rect 70802 62940 71000 62998
rect 70802 62894 70824 62940
rect 70870 62894 70928 62940
rect 70974 62894 71000 62940
rect 70802 62836 71000 62894
rect 70802 62790 70824 62836
rect 70870 62790 70928 62836
rect 70974 62790 71000 62836
rect 70802 62732 71000 62790
rect 70802 62686 70824 62732
rect 70870 62686 70928 62732
rect 70974 62686 71000 62732
rect 70802 62628 71000 62686
rect 70802 62582 70824 62628
rect 70870 62582 70928 62628
rect 70974 62582 71000 62628
rect 70802 62524 71000 62582
rect 70802 62478 70824 62524
rect 70870 62478 70928 62524
rect 70974 62478 71000 62524
rect 70802 62420 71000 62478
rect 70802 62374 70824 62420
rect 70870 62374 70928 62420
rect 70974 62374 71000 62420
rect 70802 62316 71000 62374
rect 70802 62270 70824 62316
rect 70870 62270 70928 62316
rect 70974 62270 71000 62316
rect 70802 62212 71000 62270
rect 70802 62166 70824 62212
rect 70870 62166 70928 62212
rect 70974 62166 71000 62212
rect 70802 62108 71000 62166
rect 70802 62062 70824 62108
rect 70870 62062 70928 62108
rect 70974 62062 71000 62108
rect 70802 62004 71000 62062
rect 70802 61958 70824 62004
rect 70870 61958 70928 62004
rect 70974 61958 71000 62004
rect 70802 61900 71000 61958
rect 70802 61854 70824 61900
rect 70870 61854 70928 61900
rect 70974 61854 71000 61900
rect 70802 61796 71000 61854
rect 70802 61750 70824 61796
rect 70870 61750 70928 61796
rect 70974 61750 71000 61796
rect 70802 61692 71000 61750
rect 70802 61646 70824 61692
rect 70870 61646 70928 61692
rect 70974 61646 71000 61692
rect 70802 61588 71000 61646
rect 70802 61542 70824 61588
rect 70870 61542 70928 61588
rect 70974 61542 71000 61588
rect 70802 61484 71000 61542
rect 70802 61438 70824 61484
rect 70870 61438 70928 61484
rect 70974 61438 71000 61484
rect 70802 61380 71000 61438
rect 70802 61334 70824 61380
rect 70870 61334 70928 61380
rect 70974 61334 71000 61380
rect 70802 61276 71000 61334
rect 70802 61230 70824 61276
rect 70870 61230 70928 61276
rect 70974 61230 71000 61276
rect 70802 61172 71000 61230
rect 70802 61126 70824 61172
rect 70870 61126 70928 61172
rect 70974 61126 71000 61172
rect 70802 61068 71000 61126
rect 70802 61022 70824 61068
rect 70870 61022 70928 61068
rect 70974 61022 71000 61068
rect 70802 60964 71000 61022
rect 70802 60918 70824 60964
rect 70870 60918 70928 60964
rect 70974 60918 71000 60964
rect 70802 60860 71000 60918
rect 70802 60814 70824 60860
rect 70870 60814 70928 60860
rect 70974 60814 71000 60860
rect 70802 60756 71000 60814
rect 70802 60710 70824 60756
rect 70870 60710 70928 60756
rect 70974 60710 71000 60756
rect 70802 60652 71000 60710
rect 70802 60606 70824 60652
rect 70870 60606 70928 60652
rect 70974 60606 71000 60652
rect 70802 60548 71000 60606
rect 70802 60502 70824 60548
rect 70870 60502 70928 60548
rect 70974 60502 71000 60548
rect 70802 60444 71000 60502
rect 70802 60398 70824 60444
rect 70870 60398 70928 60444
rect 70974 60398 71000 60444
rect 70802 60340 71000 60398
rect 70802 60294 70824 60340
rect 70870 60294 70928 60340
rect 70974 60294 71000 60340
rect 70802 60236 71000 60294
rect 70802 60190 70824 60236
rect 70870 60190 70928 60236
rect 70974 60190 71000 60236
rect 70802 60132 71000 60190
rect 70802 60086 70824 60132
rect 70870 60086 70928 60132
rect 70974 60086 71000 60132
rect 70802 60028 71000 60086
rect 70802 59982 70824 60028
rect 70870 59982 70928 60028
rect 70974 59982 71000 60028
rect 70802 59924 71000 59982
rect 70802 59878 70824 59924
rect 70870 59878 70928 59924
rect 70974 59878 71000 59924
rect 70802 59820 71000 59878
rect 70802 59774 70824 59820
rect 70870 59774 70928 59820
rect 70974 59774 71000 59820
rect 70802 59716 71000 59774
rect 70802 59670 70824 59716
rect 70870 59670 70928 59716
rect 70974 59670 71000 59716
rect 70802 59612 71000 59670
rect 70802 59566 70824 59612
rect 70870 59566 70928 59612
rect 70974 59566 71000 59612
rect 70802 59508 71000 59566
rect 70802 59462 70824 59508
rect 70870 59462 70928 59508
rect 70974 59462 71000 59508
rect 70802 59404 71000 59462
rect 70802 59358 70824 59404
rect 70870 59358 70928 59404
rect 70974 59358 71000 59404
rect 70802 59300 71000 59358
rect 70802 59254 70824 59300
rect 70870 59254 70928 59300
rect 70974 59254 71000 59300
rect 70802 59196 71000 59254
rect 70802 59150 70824 59196
rect 70870 59150 70928 59196
rect 70974 59150 71000 59196
rect 70802 59092 71000 59150
rect 70802 59046 70824 59092
rect 70870 59046 70928 59092
rect 70974 59046 71000 59092
rect 70802 58988 71000 59046
rect 70802 58942 70824 58988
rect 70870 58942 70928 58988
rect 70974 58942 71000 58988
rect 70802 58884 71000 58942
rect 70802 58838 70824 58884
rect 70870 58838 70928 58884
rect 70974 58838 71000 58884
rect 70802 58780 71000 58838
rect 70802 58734 70824 58780
rect 70870 58734 70928 58780
rect 70974 58734 71000 58780
rect 70802 58676 71000 58734
rect 70802 58630 70824 58676
rect 70870 58630 70928 58676
rect 70974 58630 71000 58676
rect 70802 58572 71000 58630
rect 70802 58526 70824 58572
rect 70870 58526 70928 58572
rect 70974 58526 71000 58572
rect 70802 58468 71000 58526
rect 70802 58422 70824 58468
rect 70870 58422 70928 58468
rect 70974 58422 71000 58468
rect 70802 58364 71000 58422
rect 70802 58318 70824 58364
rect 70870 58318 70928 58364
rect 70974 58318 71000 58364
rect 70802 58260 71000 58318
rect 70802 58214 70824 58260
rect 70870 58214 70928 58260
rect 70974 58214 71000 58260
rect 70802 58156 71000 58214
rect 70802 58110 70824 58156
rect 70870 58110 70928 58156
rect 70974 58110 71000 58156
rect 70802 58052 71000 58110
rect 70802 58006 70824 58052
rect 70870 58006 70928 58052
rect 70974 58006 71000 58052
rect 70802 57948 71000 58006
rect 70802 57902 70824 57948
rect 70870 57902 70928 57948
rect 70974 57902 71000 57948
rect 70802 57844 71000 57902
rect 70802 57798 70824 57844
rect 70870 57798 70928 57844
rect 70974 57798 71000 57844
rect 70802 57740 71000 57798
rect 70802 57694 70824 57740
rect 70870 57694 70928 57740
rect 70974 57694 71000 57740
rect 70802 57636 71000 57694
rect 70802 57590 70824 57636
rect 70870 57590 70928 57636
rect 70974 57590 71000 57636
rect 70802 57532 71000 57590
rect 70802 57486 70824 57532
rect 70870 57486 70928 57532
rect 70974 57486 71000 57532
rect 70802 57428 71000 57486
rect 70802 57382 70824 57428
rect 70870 57382 70928 57428
rect 70974 57382 71000 57428
rect 70802 57324 71000 57382
rect 70802 57278 70824 57324
rect 70870 57278 70928 57324
rect 70974 57278 71000 57324
rect 70802 57220 71000 57278
rect 70802 57174 70824 57220
rect 70870 57174 70928 57220
rect 70974 57174 71000 57220
rect 70802 57116 71000 57174
rect 70802 57070 70824 57116
rect 70870 57070 70928 57116
rect 70974 57070 71000 57116
rect 70802 57012 71000 57070
rect 70802 56966 70824 57012
rect 70870 56966 70928 57012
rect 70974 56966 71000 57012
rect 70802 56908 71000 56966
rect 70802 56862 70824 56908
rect 70870 56862 70928 56908
rect 70974 56862 71000 56908
rect 70802 56804 71000 56862
rect 70802 56758 70824 56804
rect 70870 56758 70928 56804
rect 70974 56758 71000 56804
rect 70802 56700 71000 56758
rect 70802 56654 70824 56700
rect 70870 56654 70928 56700
rect 70974 56654 71000 56700
rect 70802 56596 71000 56654
rect 70802 56550 70824 56596
rect 70870 56550 70928 56596
rect 70974 56550 71000 56596
rect 70802 56492 71000 56550
rect 70802 56446 70824 56492
rect 70870 56446 70928 56492
rect 70974 56446 71000 56492
rect 70802 56388 71000 56446
rect 70802 56342 70824 56388
rect 70870 56342 70928 56388
rect 70974 56342 71000 56388
rect 70802 56284 71000 56342
rect 70802 56238 70824 56284
rect 70870 56238 70928 56284
rect 70974 56238 71000 56284
rect 70802 56180 71000 56238
rect 70802 56134 70824 56180
rect 70870 56134 70928 56180
rect 70974 56134 71000 56180
rect 70802 56076 71000 56134
rect 70802 56030 70824 56076
rect 70870 56030 70928 56076
rect 70974 56030 71000 56076
rect 70802 55972 71000 56030
rect 70802 55926 70824 55972
rect 70870 55926 70928 55972
rect 70974 55926 71000 55972
rect 70802 55868 71000 55926
rect 70802 55822 70824 55868
rect 70870 55822 70928 55868
rect 70974 55822 71000 55868
rect 70802 55764 71000 55822
rect 70802 55718 70824 55764
rect 70870 55718 70928 55764
rect 70974 55718 71000 55764
rect 70802 55660 71000 55718
rect 70802 55614 70824 55660
rect 70870 55614 70928 55660
rect 70974 55614 71000 55660
rect 70802 55556 71000 55614
rect 70802 55510 70824 55556
rect 70870 55510 70928 55556
rect 70974 55510 71000 55556
rect 70802 55452 71000 55510
rect 70802 55406 70824 55452
rect 70870 55406 70928 55452
rect 70974 55406 71000 55452
rect 70802 55348 71000 55406
rect 70802 55302 70824 55348
rect 70870 55302 70928 55348
rect 70974 55302 71000 55348
rect 70802 55244 71000 55302
rect 70802 55198 70824 55244
rect 70870 55198 70928 55244
rect 70974 55198 71000 55244
rect 70802 55140 71000 55198
rect 70802 55094 70824 55140
rect 70870 55094 70928 55140
rect 70974 55094 71000 55140
rect 70802 55036 71000 55094
rect 70802 54990 70824 55036
rect 70870 54990 70928 55036
rect 70974 54990 71000 55036
rect 70802 54932 71000 54990
rect 70802 54886 70824 54932
rect 70870 54886 70928 54932
rect 70974 54886 71000 54932
rect 70802 54828 71000 54886
rect 70802 54782 70824 54828
rect 70870 54782 70928 54828
rect 70974 54782 71000 54828
rect 70802 54724 71000 54782
rect 70802 54678 70824 54724
rect 70870 54678 70928 54724
rect 70974 54678 71000 54724
rect 70802 54620 71000 54678
rect 70802 54574 70824 54620
rect 70870 54574 70928 54620
rect 70974 54574 71000 54620
rect 70802 54516 71000 54574
rect 70802 54470 70824 54516
rect 70870 54470 70928 54516
rect 70974 54470 71000 54516
rect 70802 54412 71000 54470
rect 70802 54366 70824 54412
rect 70870 54366 70928 54412
rect 70974 54366 71000 54412
rect 70802 54308 71000 54366
rect 70802 54262 70824 54308
rect 70870 54262 70928 54308
rect 70974 54262 71000 54308
rect 70802 54204 71000 54262
rect 70802 54158 70824 54204
rect 70870 54158 70928 54204
rect 70974 54158 71000 54204
rect 70802 54100 71000 54158
rect 70802 54054 70824 54100
rect 70870 54054 70928 54100
rect 70974 54054 71000 54100
rect 70802 53996 71000 54054
rect 70802 53950 70824 53996
rect 70870 53950 70928 53996
rect 70974 53950 71000 53996
rect 70802 53892 71000 53950
rect 70802 53846 70824 53892
rect 70870 53846 70928 53892
rect 70974 53846 71000 53892
rect 70802 53788 71000 53846
rect 70802 53742 70824 53788
rect 70870 53742 70928 53788
rect 70974 53742 71000 53788
rect 70802 53684 71000 53742
rect 70802 53638 70824 53684
rect 70870 53638 70928 53684
rect 70974 53638 71000 53684
rect 70802 53580 71000 53638
rect 70802 53534 70824 53580
rect 70870 53534 70928 53580
rect 70974 53534 71000 53580
rect 70802 53476 71000 53534
rect 70802 53430 70824 53476
rect 70870 53430 70928 53476
rect 70974 53430 71000 53476
rect 70802 53372 71000 53430
rect 70802 53326 70824 53372
rect 70870 53326 70928 53372
rect 70974 53326 71000 53372
rect 70802 53268 71000 53326
rect 70802 53222 70824 53268
rect 70870 53222 70928 53268
rect 70974 53222 71000 53268
rect 70802 53164 71000 53222
rect 70802 53118 70824 53164
rect 70870 53118 70928 53164
rect 70974 53118 71000 53164
rect 70802 53060 71000 53118
rect 70802 53014 70824 53060
rect 70870 53014 70928 53060
rect 70974 53014 71000 53060
rect 70802 52956 71000 53014
rect 70802 52910 70824 52956
rect 70870 52910 70928 52956
rect 70974 52910 71000 52956
rect 70802 52852 71000 52910
rect 70802 52806 70824 52852
rect 70870 52806 70928 52852
rect 70974 52806 71000 52852
rect 70802 52748 71000 52806
rect 70802 52702 70824 52748
rect 70870 52702 70928 52748
rect 70974 52702 71000 52748
rect 70802 52644 71000 52702
rect 70802 52598 70824 52644
rect 70870 52598 70928 52644
rect 70974 52598 71000 52644
rect 70802 52540 71000 52598
rect 70802 52494 70824 52540
rect 70870 52494 70928 52540
rect 70974 52494 71000 52540
rect 70802 52436 71000 52494
rect 70802 52390 70824 52436
rect 70870 52390 70928 52436
rect 70974 52390 71000 52436
rect 70802 52332 71000 52390
rect 70802 52286 70824 52332
rect 70870 52286 70928 52332
rect 70974 52286 71000 52332
rect 70802 52228 71000 52286
rect 70802 52182 70824 52228
rect 70870 52182 70928 52228
rect 70974 52182 71000 52228
rect 70802 52124 71000 52182
rect 70802 52078 70824 52124
rect 70870 52078 70928 52124
rect 70974 52078 71000 52124
rect 70802 52020 71000 52078
rect 70802 51974 70824 52020
rect 70870 51974 70928 52020
rect 70974 51974 71000 52020
rect 70802 51916 71000 51974
rect 70802 51870 70824 51916
rect 70870 51870 70928 51916
rect 70974 51870 71000 51916
rect 70802 51812 71000 51870
rect 70802 51766 70824 51812
rect 70870 51766 70928 51812
rect 70974 51766 71000 51812
rect 70802 51708 71000 51766
rect 70802 51662 70824 51708
rect 70870 51662 70928 51708
rect 70974 51662 71000 51708
rect 70802 51604 71000 51662
rect 70802 51558 70824 51604
rect 70870 51558 70928 51604
rect 70974 51558 71000 51604
rect 70802 51500 71000 51558
rect 70802 51454 70824 51500
rect 70870 51454 70928 51500
rect 70974 51454 71000 51500
rect 70802 51396 71000 51454
rect 70802 51350 70824 51396
rect 70870 51350 70928 51396
rect 70974 51350 71000 51396
rect 70802 51292 71000 51350
rect 70802 51246 70824 51292
rect 70870 51246 70928 51292
rect 70974 51246 71000 51292
rect 70802 51188 71000 51246
rect 70802 51142 70824 51188
rect 70870 51142 70928 51188
rect 70974 51142 71000 51188
rect 70802 51084 71000 51142
rect 70802 51038 70824 51084
rect 70870 51038 70928 51084
rect 70974 51038 71000 51084
rect 70802 50980 71000 51038
rect 70802 50934 70824 50980
rect 70870 50934 70928 50980
rect 70974 50934 71000 50980
rect 70802 50876 71000 50934
rect 70802 50830 70824 50876
rect 70870 50830 70928 50876
rect 70974 50830 71000 50876
rect 70802 50772 71000 50830
rect 70802 50726 70824 50772
rect 70870 50726 70928 50772
rect 70974 50726 71000 50772
rect 70802 50668 71000 50726
rect 70802 50622 70824 50668
rect 70870 50622 70928 50668
rect 70974 50622 71000 50668
rect 70802 50564 71000 50622
rect 70802 50518 70824 50564
rect 70870 50518 70928 50564
rect 70974 50518 71000 50564
rect 70802 50460 71000 50518
rect 70802 50414 70824 50460
rect 70870 50414 70928 50460
rect 70974 50414 71000 50460
rect 70802 50356 71000 50414
rect 70802 50310 70824 50356
rect 70870 50310 70928 50356
rect 70974 50310 71000 50356
rect 70802 50252 71000 50310
rect 70802 50206 70824 50252
rect 70870 50206 70928 50252
rect 70974 50206 71000 50252
rect 70802 50148 71000 50206
rect 70802 50102 70824 50148
rect 70870 50102 70928 50148
rect 70974 50102 71000 50148
rect 70802 50044 71000 50102
rect 70802 49998 70824 50044
rect 70870 49998 70928 50044
rect 70974 49998 71000 50044
rect 70802 49940 71000 49998
rect 70802 49894 70824 49940
rect 70870 49894 70928 49940
rect 70974 49894 71000 49940
rect 70802 49836 71000 49894
rect 70802 49790 70824 49836
rect 70870 49790 70928 49836
rect 70974 49790 71000 49836
rect 70802 49732 71000 49790
rect 70802 49686 70824 49732
rect 70870 49686 70928 49732
rect 70974 49686 71000 49732
rect 70802 49628 71000 49686
rect 70802 49582 70824 49628
rect 70870 49582 70928 49628
rect 70974 49582 71000 49628
rect 70802 49524 71000 49582
rect 70802 49478 70824 49524
rect 70870 49478 70928 49524
rect 70974 49478 71000 49524
rect 70802 49420 71000 49478
rect 70802 49374 70824 49420
rect 70870 49374 70928 49420
rect 70974 49374 71000 49420
rect 70802 49316 71000 49374
rect 70802 49270 70824 49316
rect 70870 49270 70928 49316
rect 70974 49270 71000 49316
rect 70802 49212 71000 49270
rect 70802 49166 70824 49212
rect 70870 49166 70928 49212
rect 70974 49166 71000 49212
rect 70802 49108 71000 49166
rect 70802 49062 70824 49108
rect 70870 49062 70928 49108
rect 70974 49062 71000 49108
rect 70802 49004 71000 49062
rect 70802 48958 70824 49004
rect 70870 48958 70928 49004
rect 70974 48958 71000 49004
rect 70802 48900 71000 48958
rect 70802 48854 70824 48900
rect 70870 48854 70928 48900
rect 70974 48854 71000 48900
rect 70802 48796 71000 48854
rect 70802 48750 70824 48796
rect 70870 48750 70928 48796
rect 70974 48750 71000 48796
rect 70802 48692 71000 48750
rect 70802 48646 70824 48692
rect 70870 48646 70928 48692
rect 70974 48646 71000 48692
rect 70802 48588 71000 48646
rect 70802 48542 70824 48588
rect 70870 48542 70928 48588
rect 70974 48542 71000 48588
rect 70802 48484 71000 48542
rect 70802 48438 70824 48484
rect 70870 48438 70928 48484
rect 70974 48438 71000 48484
rect 70802 48380 71000 48438
rect 70802 48334 70824 48380
rect 70870 48334 70928 48380
rect 70974 48334 71000 48380
rect 70802 48276 71000 48334
rect 70802 48230 70824 48276
rect 70870 48230 70928 48276
rect 70974 48230 71000 48276
rect 70802 48172 71000 48230
rect 70802 48126 70824 48172
rect 70870 48126 70928 48172
rect 70974 48126 71000 48172
rect 70802 48068 71000 48126
rect 70802 48022 70824 48068
rect 70870 48022 70928 48068
rect 70974 48022 71000 48068
rect 70802 47964 71000 48022
rect 70802 47918 70824 47964
rect 70870 47918 70928 47964
rect 70974 47918 71000 47964
rect 70802 47860 71000 47918
rect 70802 47814 70824 47860
rect 70870 47814 70928 47860
rect 70974 47814 71000 47860
rect 70802 47756 71000 47814
rect 70802 47710 70824 47756
rect 70870 47710 70928 47756
rect 70974 47710 71000 47756
rect 70802 47652 71000 47710
rect 70802 47606 70824 47652
rect 70870 47606 70928 47652
rect 70974 47606 71000 47652
rect 70802 47548 71000 47606
rect 70802 47502 70824 47548
rect 70870 47502 70928 47548
rect 70974 47502 71000 47548
rect 70802 47444 71000 47502
rect 70802 47398 70824 47444
rect 70870 47398 70928 47444
rect 70974 47398 71000 47444
rect 70802 47340 71000 47398
rect 70802 47294 70824 47340
rect 70870 47294 70928 47340
rect 70974 47294 71000 47340
rect 70802 47236 71000 47294
rect 70802 47190 70824 47236
rect 70870 47190 70928 47236
rect 70974 47190 71000 47236
rect 70802 47132 71000 47190
rect 70802 47086 70824 47132
rect 70870 47086 70928 47132
rect 70974 47086 71000 47132
rect 70802 47028 71000 47086
rect 70802 46982 70824 47028
rect 70870 46982 70928 47028
rect 70974 46982 71000 47028
rect 70802 46924 71000 46982
rect 70802 46878 70824 46924
rect 70870 46878 70928 46924
rect 70974 46878 71000 46924
rect 70802 46820 71000 46878
rect 70802 46774 70824 46820
rect 70870 46774 70928 46820
rect 70974 46774 71000 46820
rect 70802 46716 71000 46774
rect 70802 46670 70824 46716
rect 70870 46670 70928 46716
rect 70974 46670 71000 46716
rect 70802 46612 71000 46670
rect 70802 46566 70824 46612
rect 70870 46566 70928 46612
rect 70974 46566 71000 46612
rect 70802 46508 71000 46566
rect 70802 46462 70824 46508
rect 70870 46462 70928 46508
rect 70974 46462 71000 46508
rect 70802 46404 71000 46462
rect 70802 46358 70824 46404
rect 70870 46358 70928 46404
rect 70974 46358 71000 46404
rect 70802 46300 71000 46358
rect 70802 46254 70824 46300
rect 70870 46254 70928 46300
rect 70974 46254 71000 46300
rect 70802 46196 71000 46254
rect 70802 46150 70824 46196
rect 70870 46150 70928 46196
rect 70974 46150 71000 46196
rect 70802 46092 71000 46150
rect 70802 46046 70824 46092
rect 70870 46046 70928 46092
rect 70974 46046 71000 46092
rect 70802 45988 71000 46046
rect 70802 45942 70824 45988
rect 70870 45942 70928 45988
rect 70974 45942 71000 45988
rect 70802 45884 71000 45942
rect 70802 45838 70824 45884
rect 70870 45838 70928 45884
rect 70974 45838 71000 45884
rect 70802 45780 71000 45838
rect 70802 45734 70824 45780
rect 70870 45734 70928 45780
rect 70974 45734 71000 45780
rect 70802 45676 71000 45734
rect 70802 45630 70824 45676
rect 70870 45630 70928 45676
rect 70974 45630 71000 45676
rect 70802 45572 71000 45630
rect 70802 45526 70824 45572
rect 70870 45526 70928 45572
rect 70974 45526 71000 45572
rect 70802 45468 71000 45526
rect 70802 45422 70824 45468
rect 70870 45422 70928 45468
rect 70974 45422 71000 45468
rect 70802 45364 71000 45422
rect 70802 45318 70824 45364
rect 70870 45318 70928 45364
rect 70974 45318 71000 45364
rect 70802 45260 71000 45318
rect 70802 45214 70824 45260
rect 70870 45214 70928 45260
rect 70974 45214 71000 45260
rect 70802 45156 71000 45214
rect 70802 45110 70824 45156
rect 70870 45110 70928 45156
rect 70974 45110 71000 45156
rect 70802 45052 71000 45110
rect 70802 45006 70824 45052
rect 70870 45006 70928 45052
rect 70974 45006 71000 45052
rect 70802 44948 71000 45006
tri 13097 44708 13232 44843 ne
rect 13232 44837 13291 44843
tri 13291 44837 13379 44925 sw
rect 70802 44902 70824 44948
rect 70870 44902 70928 44948
rect 70974 44902 71000 44948
rect 70802 44844 71000 44902
rect 13232 44824 13379 44837
rect 13232 44778 13254 44824
rect 13300 44778 13379 44824
rect 13232 44708 13379 44778
tri 13232 44561 13379 44708 ne
tri 13379 44696 13520 44837 sw
rect 70802 44798 70824 44844
rect 70870 44798 70928 44844
rect 70974 44798 71000 44844
rect 70802 44740 71000 44798
rect 13379 44692 13520 44696
rect 13379 44646 13386 44692
rect 13432 44646 13520 44692
rect 13379 44561 13520 44646
tri 13520 44561 13655 44696 sw
rect 70802 44694 70824 44740
rect 70870 44694 70928 44740
rect 70974 44694 71000 44740
rect 70802 44636 71000 44694
rect 70802 44590 70824 44636
rect 70870 44590 70928 44636
rect 70974 44590 71000 44636
tri 13379 44466 13474 44561 ne
rect 13474 44560 13655 44561
rect 13474 44514 13518 44560
rect 13564 44514 13655 44560
rect 13474 44466 13655 44514
tri 13474 44290 13650 44466 ne
rect 13650 44451 13655 44466
tri 13655 44451 13765 44561 sw
rect 70802 44532 71000 44590
rect 70802 44486 70824 44532
rect 70870 44486 70928 44532
rect 70974 44486 71000 44532
rect 13650 44428 13765 44451
rect 13696 44382 13765 44428
rect 13650 44330 13765 44382
tri 13765 44330 13886 44451 sw
rect 70802 44428 71000 44486
rect 70802 44382 70824 44428
rect 70870 44382 70928 44428
rect 70974 44382 71000 44428
rect 13650 44296 13886 44330
rect 13650 44290 13782 44296
tri 13650 44175 13765 44290 ne
rect 13765 44250 13782 44290
rect 13828 44250 13886 44296
rect 13765 44175 13886 44250
tri 13886 44175 14041 44330 sw
rect 70802 44324 71000 44382
rect 70802 44278 70824 44324
rect 70870 44278 70928 44324
rect 70974 44278 71000 44324
rect 70802 44220 71000 44278
tri 13765 44069 13871 44175 ne
rect 13871 44164 14041 44175
rect 13871 44118 13914 44164
rect 13960 44118 14041 44164
rect 13871 44069 14041 44118
tri 13871 43919 14021 44069 ne
rect 14021 44054 14041 44069
tri 14041 44054 14162 44175 sw
rect 70802 44174 70824 44220
rect 70870 44174 70928 44220
rect 70974 44174 71000 44220
rect 70802 44116 71000 44174
rect 70802 44070 70824 44116
rect 70870 44070 70928 44116
rect 70974 44070 71000 44116
rect 14021 44032 14162 44054
rect 14021 43986 14046 44032
rect 14092 43986 14162 44032
rect 14021 43919 14162 43986
tri 14162 43919 14297 44054 sw
rect 70802 44012 71000 44070
rect 70802 43966 70824 44012
rect 70870 43966 70928 44012
rect 70974 43966 71000 44012
tri 14021 43764 14176 43919 ne
rect 14176 43900 14297 43919
rect 14176 43854 14178 43900
rect 14224 43854 14297 43900
rect 14176 43809 14297 43854
tri 14297 43809 14407 43919 sw
rect 70802 43908 71000 43966
rect 70802 43862 70824 43908
rect 70870 43862 70928 43908
rect 70974 43862 71000 43908
rect 14176 43768 14407 43809
rect 14176 43764 14310 43768
tri 14176 43646 14294 43764 ne
rect 14294 43722 14310 43764
rect 14356 43722 14407 43768
rect 14294 43646 14407 43722
tri 14294 43556 14384 43646 ne
rect 14384 43643 14407 43646
tri 14407 43643 14573 43809 sw
rect 70802 43804 71000 43862
rect 70802 43758 70824 43804
rect 70870 43758 70928 43804
rect 70974 43758 71000 43804
rect 70802 43700 71000 43758
rect 70802 43654 70824 43700
rect 70870 43654 70928 43700
rect 70974 43654 71000 43700
rect 14384 43636 14573 43643
rect 14384 43590 14442 43636
rect 14488 43590 14573 43636
rect 14384 43556 14573 43590
tri 14384 43398 14542 43556 ne
rect 14542 43547 14573 43556
tri 14573 43547 14669 43643 sw
rect 70802 43596 71000 43654
rect 70802 43550 70824 43596
rect 70870 43550 70928 43596
rect 70974 43550 71000 43596
rect 14542 43504 14669 43547
rect 14542 43458 14574 43504
rect 14620 43458 14669 43504
rect 14542 43398 14669 43458
tri 14669 43398 14818 43547 sw
rect 70802 43492 71000 43550
rect 70802 43446 70824 43492
rect 70870 43446 70928 43492
rect 70974 43446 71000 43492
tri 14542 43237 14703 43398 ne
rect 14703 43372 14818 43398
rect 14703 43326 14706 43372
rect 14752 43326 14818 43372
rect 14703 43271 14818 43326
tri 14818 43271 14945 43398 sw
rect 70802 43388 71000 43446
rect 70802 43342 70824 43388
rect 70870 43342 70928 43388
rect 70974 43342 71000 43388
rect 70802 43284 71000 43342
rect 14703 43240 14945 43271
rect 14703 43237 14838 43240
tri 14703 43122 14818 43237 ne
rect 14818 43194 14838 43237
rect 14884 43194 14945 43240
rect 14818 43122 14945 43194
tri 14945 43122 15094 43271 sw
rect 70802 43238 70824 43284
rect 70870 43238 70928 43284
rect 70974 43238 71000 43284
rect 70802 43180 71000 43238
rect 70802 43134 70824 43180
rect 70870 43134 70928 43180
rect 70974 43134 71000 43180
tri 14818 42971 14969 43122 ne
rect 14969 43108 15094 43122
rect 14969 43062 14970 43108
rect 15016 43062 15094 43108
rect 14969 42987 15094 43062
tri 15094 42987 15229 43122 sw
rect 70802 43076 71000 43134
rect 70802 43030 70824 43076
rect 70870 43030 70928 43076
rect 70974 43030 71000 43076
rect 14969 42976 15229 42987
rect 14969 42971 15102 42976
tri 14969 42860 15080 42971 ne
rect 15080 42930 15102 42971
rect 15148 42930 15229 42976
rect 15080 42860 15229 42930
tri 15229 42860 15356 42987 sw
rect 70802 42972 71000 43030
rect 70802 42926 70824 42972
rect 70870 42926 70928 42972
rect 70974 42926 71000 42972
rect 70802 42868 71000 42926
tri 15080 42711 15229 42860 ne
rect 15229 42844 15356 42860
rect 15229 42798 15234 42844
rect 15280 42798 15356 42844
rect 15229 42756 15356 42798
tri 15356 42756 15460 42860 sw
rect 70802 42822 70824 42868
rect 70870 42822 70928 42868
rect 70974 42822 71000 42868
rect 70802 42764 71000 42822
rect 15229 42712 15460 42756
rect 15229 42711 15366 42712
tri 15229 42584 15356 42711 ne
rect 15356 42666 15366 42711
rect 15412 42666 15460 42712
rect 15356 42584 15460 42666
tri 15460 42584 15632 42756 sw
rect 70802 42718 70824 42764
rect 70870 42718 70928 42764
rect 70974 42718 71000 42764
rect 70802 42660 71000 42718
rect 70802 42614 70824 42660
rect 70870 42614 70928 42660
rect 70974 42614 71000 42660
tri 15356 42462 15478 42584 ne
rect 15478 42580 15632 42584
rect 15478 42534 15498 42580
rect 15544 42534 15632 42580
rect 15478 42488 15632 42534
tri 15632 42488 15728 42584 sw
rect 70802 42556 71000 42614
rect 70802 42510 70824 42556
rect 70870 42510 70928 42556
rect 70974 42510 71000 42556
rect 15478 42462 15728 42488
tri 15478 42345 15595 42462 ne
rect 15595 42448 15728 42462
rect 15595 42402 15630 42448
rect 15676 42402 15728 42448
rect 15595 42345 15728 42402
tri 15728 42345 15871 42488 sw
rect 70802 42452 71000 42510
rect 70802 42406 70824 42452
rect 70870 42406 70928 42452
rect 70974 42406 71000 42452
rect 70802 42348 71000 42406
tri 15595 42187 15753 42345 ne
rect 15753 42316 15871 42345
rect 15753 42270 15762 42316
rect 15808 42270 15871 42316
rect 15753 42210 15871 42270
tri 15871 42210 16006 42345 sw
rect 70802 42302 70824 42348
rect 70870 42302 70928 42348
rect 70974 42302 71000 42348
rect 70802 42244 71000 42302
rect 15753 42187 16006 42210
tri 15753 42077 15863 42187 ne
rect 15863 42184 16006 42187
rect 15863 42138 15894 42184
rect 15940 42138 16006 42184
rect 15863 42077 16006 42138
tri 16006 42077 16139 42210 sw
rect 70802 42198 70824 42244
rect 70870 42198 70928 42244
rect 70974 42198 71000 42244
rect 70802 42140 71000 42198
rect 70802 42094 70824 42140
rect 70870 42094 70928 42140
rect 70974 42094 71000 42140
tri 15863 41934 16006 42077 ne
rect 16006 42052 16139 42077
rect 16006 42006 16026 42052
rect 16072 42006 16139 42052
rect 16006 41934 16139 42006
tri 16139 41934 16282 42077 sw
rect 70802 42036 71000 42094
rect 70802 41990 70824 42036
rect 70870 41990 70928 42036
rect 70974 41990 71000 42036
tri 16006 41801 16139 41934 ne
rect 16139 41920 16282 41934
rect 16139 41874 16158 41920
rect 16204 41874 16282 41920
rect 16139 41801 16282 41874
tri 16282 41801 16415 41934 sw
rect 70802 41932 71000 41990
rect 70802 41886 70824 41932
rect 70870 41886 70928 41932
rect 70974 41886 71000 41932
rect 70802 41828 71000 41886
tri 16139 41658 16282 41801 ne
rect 16282 41788 16415 41801
rect 16282 41742 16290 41788
rect 16336 41742 16415 41788
rect 16282 41658 16415 41742
tri 16415 41658 16558 41801 sw
rect 70802 41782 70824 41828
rect 70870 41782 70928 41828
rect 70974 41782 71000 41828
rect 70802 41724 71000 41782
rect 70802 41678 70824 41724
rect 70870 41678 70928 41724
rect 70974 41678 71000 41724
tri 16282 41525 16415 41658 ne
rect 16415 41656 16558 41658
rect 16415 41610 16422 41656
rect 16468 41610 16558 41656
rect 16415 41525 16558 41610
tri 16558 41525 16691 41658 sw
rect 70802 41620 71000 41678
rect 70802 41574 70824 41620
rect 70870 41574 70928 41620
rect 70974 41574 71000 41620
tri 16415 41413 16527 41525 ne
rect 16527 41524 16691 41525
rect 16527 41478 16554 41524
rect 16600 41478 16691 41524
rect 16527 41435 16691 41478
tri 16691 41435 16781 41525 sw
rect 70802 41516 71000 41574
rect 70802 41470 70824 41516
rect 70870 41470 70928 41516
rect 70974 41470 71000 41516
rect 16527 41413 16781 41435
tri 16527 41254 16686 41413 ne
rect 16686 41392 16781 41413
rect 16732 41346 16781 41392
rect 16686 41294 16781 41346
tri 16781 41294 16922 41435 sw
rect 70802 41412 71000 41470
rect 70802 41366 70824 41412
rect 70870 41366 70928 41412
rect 70974 41366 71000 41412
rect 70802 41308 71000 41366
rect 16686 41260 16922 41294
rect 16686 41254 16818 41260
tri 16686 41138 16802 41254 ne
rect 16802 41214 16818 41254
rect 16864 41214 16922 41260
rect 16802 41157 16922 41214
tri 16922 41157 17059 41294 sw
rect 70802 41262 70824 41308
rect 70870 41262 70928 41308
rect 70974 41262 71000 41308
rect 70802 41204 71000 41262
rect 70802 41158 70824 41204
rect 70870 41158 70928 41204
rect 70974 41158 71000 41204
rect 16802 41138 17059 41157
tri 16802 40990 16950 41138 ne
rect 16950 41128 17059 41138
rect 16996 41082 17059 41128
rect 16950 41018 17059 41082
tri 17059 41018 17198 41157 sw
rect 70802 41100 71000 41158
rect 70802 41054 70824 41100
rect 70870 41054 70928 41100
rect 70974 41054 71000 41100
rect 16950 40996 17198 41018
rect 16950 40990 17082 40996
tri 16950 40881 17059 40990 ne
rect 17059 40950 17082 40990
rect 17128 40950 17198 40996
rect 17059 40881 17198 40950
tri 17198 40881 17335 41018 sw
rect 70802 40996 71000 41054
rect 70802 40950 70824 40996
rect 70870 40950 70928 40996
rect 70974 40950 71000 40996
rect 70802 40892 71000 40950
tri 17059 40726 17214 40881 ne
rect 17214 40864 17335 40881
rect 17260 40818 17335 40864
rect 17214 40742 17335 40818
tri 17335 40742 17474 40881 sw
rect 70802 40846 70824 40892
rect 70870 40846 70928 40892
rect 70974 40846 71000 40892
rect 70802 40788 71000 40846
rect 70802 40742 70824 40788
rect 70870 40742 70928 40788
rect 70974 40742 71000 40788
rect 17214 40732 17474 40742
rect 17214 40726 17346 40732
tri 17214 40607 17333 40726 ne
rect 17333 40686 17346 40726
rect 17392 40686 17474 40732
rect 17333 40607 17474 40686
tri 17333 40470 17470 40607 ne
rect 17470 40605 17474 40607
tri 17474 40605 17611 40742 sw
rect 70802 40684 71000 40742
rect 70802 40638 70824 40684
rect 70870 40638 70928 40684
rect 70974 40638 71000 40684
rect 17470 40600 17611 40605
rect 17470 40554 17478 40600
rect 17524 40554 17611 40600
rect 17470 40470 17611 40554
tri 17611 40470 17746 40605 sw
rect 70802 40580 71000 40638
rect 70802 40534 70824 40580
rect 70870 40534 70928 40580
rect 70974 40534 71000 40580
rect 70802 40476 71000 40534
tri 17470 40363 17577 40470 ne
rect 17577 40468 17746 40470
rect 17577 40422 17610 40468
rect 17656 40422 17746 40468
rect 17577 40376 17746 40422
tri 17746 40376 17840 40470 sw
rect 70802 40430 70824 40476
rect 70870 40430 70928 40476
rect 70974 40430 71000 40476
rect 17577 40363 17840 40376
tri 17577 40228 17712 40363 ne
rect 17712 40336 17840 40363
rect 17712 40290 17742 40336
rect 17788 40290 17840 40336
rect 17712 40239 17840 40290
tri 17840 40239 17977 40376 sw
rect 70802 40372 71000 40430
rect 70802 40326 70824 40372
rect 70870 40326 70928 40372
rect 70974 40326 71000 40372
rect 70802 40268 71000 40326
rect 17712 40228 17977 40239
tri 17712 40100 17840 40228 ne
rect 17840 40204 17977 40228
rect 17840 40158 17874 40204
rect 17920 40158 17977 40204
rect 17840 40104 17977 40158
tri 17977 40104 18112 40239 sw
rect 70802 40222 70824 40268
rect 70870 40222 70928 40268
rect 70974 40222 71000 40268
rect 70802 40164 71000 40222
rect 70802 40118 70824 40164
rect 70870 40118 70928 40164
rect 70974 40118 71000 40164
rect 17840 40100 18112 40104
tri 17840 39953 17987 40100 ne
rect 17987 40072 18112 40100
rect 17987 40026 18006 40072
rect 18052 40026 18112 40072
rect 17987 39959 18112 40026
tri 18112 39959 18257 40104 sw
rect 70802 40060 71000 40118
rect 70802 40014 70824 40060
rect 70870 40014 70928 40060
rect 70974 40014 71000 40060
rect 17987 39953 18257 39959
tri 17987 39824 18116 39953 ne
rect 18116 39940 18257 39953
rect 18116 39894 18138 39940
rect 18184 39894 18257 39940
rect 18116 39828 18257 39894
tri 18257 39828 18388 39959 sw
rect 70802 39956 71000 40014
rect 70802 39910 70824 39956
rect 70870 39910 70928 39956
rect 70974 39910 71000 39956
rect 70802 39852 71000 39910
rect 18116 39824 18388 39828
tri 18116 39679 18261 39824 ne
rect 18261 39808 18388 39824
rect 18261 39762 18270 39808
rect 18316 39762 18388 39808
rect 18261 39683 18388 39762
tri 18388 39683 18533 39828 sw
rect 70802 39806 70824 39852
rect 70870 39806 70928 39852
rect 70974 39806 71000 39852
rect 70802 39748 71000 39806
rect 70802 39702 70824 39748
rect 70870 39702 70928 39748
rect 70974 39702 71000 39748
rect 18261 39679 18533 39683
tri 18261 39548 18392 39679 ne
rect 18392 39676 18533 39679
rect 18392 39630 18402 39676
rect 18448 39630 18533 39676
rect 18392 39548 18533 39630
tri 18533 39548 18668 39683 sw
rect 70802 39644 71000 39702
rect 70802 39598 70824 39644
rect 70870 39598 70928 39644
rect 70974 39598 71000 39644
tri 18392 39417 18523 39548 ne
rect 18523 39544 18668 39548
rect 18523 39498 18534 39544
rect 18580 39498 18668 39544
rect 18523 39417 18668 39498
tri 18668 39417 18799 39548 sw
rect 70802 39540 71000 39598
rect 70802 39494 70824 39540
rect 70870 39494 70928 39540
rect 70974 39494 71000 39540
rect 70802 39436 71000 39494
tri 18523 39317 18623 39417 ne
rect 18623 39412 18799 39417
rect 18623 39366 18666 39412
rect 18712 39366 18799 39412
rect 18623 39317 18799 39366
tri 18799 39317 18899 39417 sw
rect 70802 39390 70824 39436
rect 70870 39390 70928 39436
rect 70974 39390 71000 39436
rect 70802 39332 71000 39390
tri 18623 39179 18761 39317 ne
rect 18761 39280 18899 39317
rect 18761 39234 18798 39280
rect 18844 39234 18899 39280
rect 18761 39186 18899 39234
tri 18899 39186 19030 39317 sw
rect 70802 39286 70824 39332
rect 70870 39286 70928 39332
rect 70974 39286 71000 39332
rect 70802 39228 71000 39286
rect 18761 39179 19030 39186
tri 18761 39041 18899 39179 ne
rect 18899 39148 19030 39179
rect 18899 39102 18930 39148
rect 18976 39102 19030 39148
rect 18899 39041 19030 39102
tri 19030 39041 19175 39186 sw
rect 70802 39182 70824 39228
rect 70870 39182 70928 39228
rect 70974 39182 71000 39228
rect 70802 39124 71000 39182
rect 70802 39078 70824 39124
rect 70870 39078 70928 39124
rect 70974 39078 71000 39124
tri 18899 38904 19036 39041 ne
rect 19036 39016 19175 39041
rect 19036 38970 19062 39016
rect 19108 38970 19175 39016
rect 19036 38904 19175 38970
tri 19036 38765 19175 38904 ne
tri 19175 38900 19316 39041 sw
rect 70802 39020 71000 39078
rect 70802 38974 70824 39020
rect 70870 38974 70928 39020
rect 70974 38974 71000 39020
rect 70802 38916 71000 38974
rect 19175 38884 19316 38900
rect 19175 38838 19194 38884
rect 19240 38838 19316 38884
rect 19175 38765 19316 38838
tri 19316 38765 19451 38900 sw
rect 70802 38870 70824 38916
rect 70870 38870 70928 38916
rect 70974 38870 71000 38916
rect 70802 38812 71000 38870
rect 70802 38766 70824 38812
rect 70870 38766 70928 38812
rect 70974 38766 71000 38812
tri 19175 38640 19300 38765 ne
rect 19300 38752 19451 38765
rect 19300 38706 19326 38752
rect 19372 38706 19451 38752
rect 19300 38640 19451 38706
tri 19451 38640 19576 38765 sw
rect 70802 38708 71000 38766
rect 70802 38662 70824 38708
rect 70870 38662 70928 38708
rect 70974 38662 71000 38708
tri 19300 38489 19451 38640 ne
rect 19451 38620 19576 38640
rect 19451 38574 19458 38620
rect 19504 38574 19576 38620
rect 19451 38489 19576 38574
tri 19576 38489 19727 38640 sw
rect 70802 38604 71000 38662
rect 70802 38558 70824 38604
rect 70870 38558 70928 38604
rect 70974 38558 71000 38604
rect 70802 38500 71000 38558
tri 19451 38354 19586 38489 ne
rect 19586 38488 19727 38489
rect 19586 38442 19590 38488
rect 19636 38442 19727 38488
rect 19586 38364 19727 38442
tri 19727 38364 19852 38489 sw
rect 70802 38454 70824 38500
rect 70870 38454 70928 38500
rect 70974 38454 71000 38500
rect 70802 38396 71000 38454
rect 19586 38356 19852 38364
rect 19586 38354 19722 38356
tri 19586 38218 19722 38354 ne
rect 19768 38310 19852 38356
rect 19722 38258 19852 38310
tri 19852 38258 19958 38364 sw
rect 70802 38350 70824 38396
rect 70870 38350 70928 38396
rect 70974 38350 71000 38396
rect 70802 38292 71000 38350
rect 19722 38224 19958 38258
rect 19722 38218 19854 38224
tri 19722 38129 19811 38218 ne
rect 19811 38178 19854 38218
rect 19900 38178 19958 38224
rect 19811 38129 19958 38178
tri 19811 37982 19958 38129 ne
tri 19958 38123 20093 38258 sw
rect 70802 38246 70824 38292
rect 70870 38246 70928 38292
rect 70974 38246 71000 38292
rect 70802 38188 71000 38246
rect 70802 38142 70824 38188
rect 70870 38142 70928 38188
rect 70974 38142 71000 38188
rect 19958 38092 20093 38123
rect 19958 38046 19986 38092
rect 20032 38046 20093 38092
rect 19958 37998 20093 38046
tri 20093 37998 20218 38123 sw
rect 70802 38084 71000 38142
rect 70802 38038 70824 38084
rect 70870 38038 70928 38084
rect 70974 38038 71000 38084
rect 19958 37982 20218 37998
tri 19958 37855 20085 37982 ne
rect 20085 37960 20218 37982
rect 20085 37914 20118 37960
rect 20164 37914 20218 37960
rect 20085 37863 20218 37914
tri 20218 37863 20353 37998 sw
rect 70802 37980 71000 38038
rect 70802 37934 70824 37980
rect 70870 37934 70928 37980
rect 70974 37934 71000 37980
rect 70802 37876 71000 37934
rect 20085 37855 20353 37863
tri 20085 37690 20250 37855 ne
rect 20250 37828 20353 37855
rect 20296 37782 20353 37828
rect 20250 37706 20353 37782
tri 20353 37706 20510 37863 sw
rect 70802 37830 70824 37876
rect 70870 37830 70928 37876
rect 70974 37830 71000 37876
rect 70802 37772 71000 37830
rect 70802 37726 70824 37772
rect 70870 37726 70928 37772
rect 70974 37726 71000 37772
rect 20250 37696 20510 37706
rect 20250 37690 20382 37696
tri 20250 37587 20353 37690 ne
rect 20353 37650 20382 37690
rect 20428 37650 20510 37696
rect 20353 37587 20510 37650
tri 20510 37587 20629 37706 sw
rect 70802 37668 71000 37726
rect 70802 37622 70824 37668
rect 70870 37622 70928 37668
rect 70974 37622 71000 37668
tri 20353 37426 20514 37587 ne
rect 20514 37564 20629 37587
rect 20560 37518 20629 37564
rect 20514 37475 20629 37518
tri 20629 37475 20741 37587 sw
rect 70802 37564 71000 37622
rect 70802 37518 70824 37564
rect 70870 37518 70928 37564
rect 70974 37518 71000 37564
rect 20514 37432 20741 37475
rect 20514 37426 20646 37432
tri 20514 37295 20645 37426 ne
rect 20645 37386 20646 37426
rect 20692 37386 20741 37432
rect 20645 37311 20741 37386
tri 20741 37311 20905 37475 sw
rect 70802 37460 71000 37518
rect 70802 37414 70824 37460
rect 70870 37414 70928 37460
rect 70974 37414 71000 37460
rect 70802 37356 71000 37414
rect 20645 37300 20905 37311
rect 20645 37295 20778 37300
tri 20645 37162 20778 37295 ne
rect 20824 37254 20905 37300
rect 20778 37176 20905 37254
tri 20905 37176 21040 37311 sw
rect 70802 37310 70824 37356
rect 70870 37310 70928 37356
rect 70974 37310 71000 37356
rect 70802 37252 71000 37310
rect 70802 37206 70824 37252
rect 70870 37206 70928 37252
rect 70974 37206 71000 37252
rect 20778 37168 21040 37176
rect 20778 37162 20910 37168
tri 20778 37035 20905 37162 ne
rect 20905 37122 20910 37162
rect 20956 37122 21040 37168
rect 20905 37064 21040 37122
tri 21040 37064 21152 37176 sw
rect 70802 37148 71000 37206
rect 70802 37102 70824 37148
rect 70870 37102 70928 37148
rect 70974 37102 71000 37148
rect 20905 37036 21152 37064
rect 20905 37035 21042 37036
tri 20905 36900 21040 37035 ne
rect 21040 36990 21042 37035
rect 21088 36990 21152 37036
rect 21040 36945 21152 36990
tri 21152 36945 21271 37064 sw
rect 70802 37044 71000 37102
rect 70802 36998 70824 37044
rect 70870 36998 70928 37044
rect 70974 36998 71000 37044
rect 21040 36904 21271 36945
rect 21040 36900 21174 36904
tri 21040 36788 21152 36900 ne
rect 21152 36858 21174 36900
rect 21220 36858 21271 36904
rect 21152 36810 21271 36858
tri 21271 36810 21406 36945 sw
rect 70802 36940 71000 36998
rect 70802 36894 70824 36940
rect 70870 36894 70928 36940
rect 70974 36894 71000 36940
rect 70802 36836 71000 36894
rect 21152 36788 21406 36810
tri 21152 36670 21270 36788 ne
rect 21270 36772 21406 36788
rect 21270 36726 21306 36772
rect 21352 36726 21406 36772
rect 21270 36670 21406 36726
tri 21270 36534 21406 36670 ne
tri 21406 36647 21569 36810 sw
rect 70802 36790 70824 36836
rect 70870 36790 70928 36836
rect 70974 36790 71000 36836
rect 70802 36732 71000 36790
rect 70802 36686 70824 36732
rect 70870 36686 70928 36732
rect 70974 36686 71000 36732
rect 21406 36640 21569 36647
rect 21406 36594 21438 36640
rect 21484 36594 21569 36640
rect 21406 36534 21569 36594
tri 21569 36534 21682 36647 sw
rect 70802 36628 71000 36686
rect 70802 36582 70824 36628
rect 70870 36582 70928 36628
rect 70974 36582 71000 36628
tri 21406 36395 21545 36534 ne
rect 21545 36508 21682 36534
rect 21545 36462 21570 36508
rect 21616 36462 21682 36508
rect 21545 36399 21682 36462
tri 21682 36399 21817 36534 sw
rect 70802 36524 71000 36582
rect 70802 36478 70824 36524
rect 70870 36478 70928 36524
rect 70974 36478 71000 36524
rect 70802 36420 71000 36478
rect 21545 36395 21817 36399
tri 21545 36281 21659 36395 ne
rect 21659 36376 21817 36395
rect 21659 36330 21702 36376
rect 21748 36330 21817 36376
rect 21659 36281 21817 36330
tri 21817 36281 21935 36399 sw
rect 70802 36374 70824 36420
rect 70870 36374 70928 36420
rect 70974 36374 71000 36420
rect 70802 36316 71000 36374
tri 21659 36123 21817 36281 ne
rect 21817 36244 21935 36281
rect 21817 36198 21834 36244
rect 21880 36198 21935 36244
rect 21817 36123 21935 36198
tri 21935 36123 22093 36281 sw
rect 70802 36270 70824 36316
rect 70870 36270 70928 36316
rect 70974 36270 71000 36316
rect 70802 36212 71000 36270
rect 70802 36166 70824 36212
rect 70870 36166 70928 36212
rect 70974 36166 71000 36212
tri 21817 35986 21954 36123 ne
rect 21954 36112 22093 36123
rect 21954 36066 21966 36112
rect 22012 36066 22093 36112
rect 21954 36005 22093 36066
tri 22093 36005 22211 36123 sw
rect 70802 36108 71000 36166
rect 70802 36062 70824 36108
rect 70870 36062 70928 36108
rect 70974 36062 71000 36108
rect 21954 35986 22211 36005
tri 21954 35851 22089 35986 ne
rect 22089 35980 22211 35986
rect 22089 35934 22098 35980
rect 22144 35934 22211 35980
rect 22089 35892 22211 35934
tri 22211 35892 22324 36005 sw
rect 70802 36004 71000 36062
rect 70802 35958 70824 36004
rect 70870 35958 70928 36004
rect 70974 35958 71000 36004
rect 70802 35900 71000 35958
rect 22089 35851 22324 35892
tri 22089 35729 22211 35851 ne
rect 22211 35848 22324 35851
rect 22211 35802 22230 35848
rect 22276 35802 22324 35848
rect 22211 35729 22324 35802
tri 22324 35729 22487 35892 sw
rect 70802 35854 70824 35900
rect 70870 35854 70928 35900
rect 70974 35854 71000 35900
rect 70802 35796 71000 35854
rect 70802 35750 70824 35796
rect 70870 35750 70928 35796
rect 70974 35750 71000 35796
tri 22211 35621 22319 35729 ne
rect 22319 35716 22487 35729
rect 22319 35670 22362 35716
rect 22408 35670 22487 35716
rect 22319 35621 22487 35670
tri 22319 35453 22487 35621 ne
tri 22487 35588 22628 35729 sw
rect 70802 35692 71000 35750
rect 70802 35646 70824 35692
rect 70870 35646 70928 35692
rect 70974 35646 71000 35692
rect 70802 35588 71000 35646
rect 22487 35584 22628 35588
rect 22487 35538 22494 35584
rect 22540 35538 22628 35584
rect 22487 35453 22628 35538
tri 22628 35453 22763 35588 sw
rect 70802 35542 70824 35588
rect 70870 35542 70928 35588
rect 70974 35542 71000 35588
rect 70802 35484 71000 35542
tri 22487 35346 22594 35453 ne
rect 22594 35452 22763 35453
rect 22594 35406 22626 35452
rect 22672 35406 22763 35452
rect 22594 35346 22763 35406
tri 22763 35346 22870 35453 sw
rect 70802 35438 70824 35484
rect 70870 35438 70928 35484
rect 70974 35438 71000 35484
rect 70802 35380 71000 35438
tri 22594 35182 22758 35346 ne
rect 22758 35320 22870 35346
rect 22804 35274 22870 35320
rect 22758 35222 22870 35274
tri 22870 35222 22994 35346 sw
rect 70802 35334 70824 35380
rect 70870 35334 70928 35380
rect 70974 35334 71000 35380
rect 70802 35276 71000 35334
rect 70802 35230 70824 35276
rect 70870 35230 70928 35276
rect 70974 35230 71000 35276
rect 22758 35188 22994 35222
rect 22758 35182 22890 35188
tri 22758 35070 22870 35182 ne
rect 22870 35142 22890 35182
rect 22936 35142 22994 35188
rect 22870 35070 22994 35142
tri 22994 35070 23146 35222 sw
rect 70802 35172 71000 35230
rect 70802 35126 70824 35172
rect 70870 35126 70928 35172
rect 70974 35126 71000 35172
tri 22870 34918 23022 35070 ne
rect 23022 35056 23146 35070
rect 23068 35010 23146 35056
rect 23022 34946 23146 35010
tri 23146 34946 23270 35070 sw
rect 70802 35068 71000 35126
rect 70802 35022 70824 35068
rect 70870 35022 70928 35068
rect 70974 35022 71000 35068
rect 70802 34964 71000 35022
rect 23022 34924 23270 34946
rect 23022 34918 23154 34924
tri 23022 34801 23139 34918 ne
rect 23139 34878 23154 34918
rect 23200 34878 23270 34924
rect 23139 34801 23270 34878
tri 23139 34670 23270 34801 ne
tri 23270 34794 23422 34946 sw
rect 70802 34918 70824 34964
rect 70870 34918 70928 34964
rect 70974 34918 71000 34964
rect 70802 34860 71000 34918
rect 70802 34814 70824 34860
rect 70870 34814 70928 34860
rect 70974 34814 71000 34860
rect 23270 34792 23422 34794
rect 23270 34746 23286 34792
rect 23332 34746 23422 34792
rect 23270 34704 23422 34746
tri 23422 34704 23512 34794 sw
rect 70802 34756 71000 34814
rect 70802 34710 70824 34756
rect 70870 34710 70928 34756
rect 70974 34710 71000 34756
rect 23270 34670 23512 34704
tri 23270 34526 23414 34670 ne
rect 23414 34660 23512 34670
rect 23414 34614 23418 34660
rect 23464 34614 23512 34660
rect 23414 34569 23512 34614
tri 23512 34569 23647 34704 sw
rect 70802 34652 71000 34710
rect 70802 34606 70824 34652
rect 70870 34606 70928 34652
rect 70974 34606 71000 34652
rect 23414 34528 23647 34569
rect 23414 34526 23550 34528
tri 23414 34390 23550 34526 ne
rect 23596 34482 23647 34528
rect 23550 34439 23647 34482
tri 23647 34439 23777 34569 sw
rect 70802 34548 71000 34606
rect 70802 34502 70824 34548
rect 70870 34502 70928 34548
rect 70974 34502 71000 34548
rect 70802 34444 71000 34502
rect 23550 34396 23777 34439
rect 23550 34390 23682 34396
tri 23550 34293 23647 34390 ne
rect 23647 34350 23682 34390
rect 23728 34350 23777 34396
rect 23647 34293 23777 34350
tri 23777 34293 23923 34439 sw
rect 70802 34398 70824 34444
rect 70870 34398 70928 34444
rect 70974 34398 71000 34444
rect 70802 34340 71000 34398
rect 70802 34294 70824 34340
rect 70870 34294 70928 34340
rect 70974 34294 71000 34340
tri 23647 34126 23814 34293 ne
rect 23814 34264 23923 34293
rect 23860 34218 23923 34264
rect 23814 34163 23923 34218
tri 23923 34163 24053 34293 sw
rect 70802 34236 71000 34294
rect 70802 34190 70824 34236
rect 70870 34190 70928 34236
rect 70974 34190 71000 34236
rect 23814 34132 24053 34163
rect 23814 34126 23946 34132
tri 23814 34028 23912 34126 ne
rect 23912 34086 23946 34126
rect 23992 34086 24053 34132
rect 23912 34028 24053 34086
tri 23912 33927 24013 34028 ne
rect 24013 34017 24053 34028
tri 24053 34017 24199 34163 sw
rect 70802 34132 71000 34190
rect 70802 34086 70824 34132
rect 70870 34086 70928 34132
rect 70974 34086 71000 34132
rect 70802 34028 71000 34086
rect 24013 34000 24199 34017
rect 24013 33954 24078 34000
rect 24124 33954 24199 34000
rect 24013 33927 24199 33954
tri 24013 33752 24188 33927 ne
rect 24188 33882 24199 33927
tri 24199 33882 24334 34017 sw
rect 70802 33982 70824 34028
rect 70870 33982 70928 34028
rect 70974 33982 71000 34028
rect 70802 33924 71000 33982
rect 24188 33868 24334 33882
rect 24188 33822 24210 33868
rect 24256 33822 24334 33868
rect 24188 33752 24334 33822
tri 24334 33752 24464 33882 sw
rect 70802 33878 70824 33924
rect 70870 33878 70928 33924
rect 70974 33878 71000 33924
rect 70802 33820 71000 33878
rect 70802 33774 70824 33820
rect 70870 33774 70928 33820
rect 70974 33774 71000 33820
tri 24188 33606 24334 33752 ne
rect 24334 33736 24464 33752
rect 24334 33690 24342 33736
rect 24388 33690 24464 33736
rect 24334 33606 24464 33690
tri 24464 33606 24610 33752 sw
rect 70802 33716 71000 33774
rect 70802 33670 70824 33716
rect 70870 33670 70928 33716
rect 70974 33670 71000 33716
rect 70802 33612 71000 33670
tri 24334 33476 24464 33606 ne
rect 24464 33604 24610 33606
rect 24464 33558 24474 33604
rect 24520 33558 24610 33604
rect 24464 33516 24610 33558
tri 24610 33516 24700 33606 sw
rect 70802 33566 70824 33612
rect 70870 33566 70928 33612
rect 70974 33566 71000 33612
rect 24464 33476 24700 33516
tri 24464 33342 24598 33476 ne
rect 24598 33472 24700 33476
rect 24598 33426 24606 33472
rect 24652 33426 24700 33472
rect 24598 33380 24700 33426
tri 24700 33380 24836 33516 sw
rect 70802 33508 71000 33566
rect 70802 33462 70824 33508
rect 70870 33462 70928 33508
rect 70974 33462 71000 33508
rect 70802 33404 71000 33462
rect 24598 33342 24836 33380
tri 24598 33240 24700 33342 ne
rect 24700 33340 24836 33342
rect 24700 33294 24738 33340
rect 24784 33294 24836 33340
rect 24700 33240 24836 33294
tri 24836 33240 24976 33380 sw
rect 70802 33358 70824 33404
rect 70870 33358 70928 33404
rect 70974 33358 71000 33404
rect 70802 33300 71000 33358
rect 70802 33254 70824 33300
rect 70870 33254 70928 33300
rect 70974 33254 71000 33300
tri 24700 33112 24828 33240 ne
rect 24828 33208 24976 33240
rect 24828 33162 24870 33208
rect 24916 33162 24976 33208
rect 24828 33112 24976 33162
tri 24828 32969 24971 33112 ne
rect 24971 33105 24976 33112
tri 24976 33105 25111 33240 sw
rect 70802 33196 71000 33254
rect 70802 33150 70824 33196
rect 70870 33150 70928 33196
rect 70974 33150 71000 33196
rect 24971 33076 25111 33105
rect 24971 33030 25002 33076
rect 25048 33030 25111 33076
rect 24971 32969 25111 33030
tri 25111 32969 25247 33105 sw
rect 70802 33092 71000 33150
rect 70802 33046 70824 33092
rect 70870 33046 70928 33092
rect 70974 33046 71000 33092
rect 70802 32988 71000 33046
tri 24971 32829 25111 32969 ne
rect 25111 32944 25247 32969
rect 25111 32898 25134 32944
rect 25180 32898 25247 32944
rect 25111 32829 25247 32898
tri 25247 32829 25387 32969 sw
rect 70802 32942 70824 32988
rect 70870 32942 70928 32988
rect 70974 32942 71000 32988
rect 70802 32884 71000 32942
rect 70802 32838 70824 32884
rect 70870 32838 70928 32884
rect 70974 32838 71000 32884
tri 25111 32693 25247 32829 ne
rect 25247 32812 25387 32829
rect 25247 32766 25266 32812
rect 25312 32766 25387 32812
rect 25247 32693 25387 32766
tri 25387 32693 25523 32829 sw
rect 70802 32780 71000 32838
rect 70802 32734 70824 32780
rect 70870 32734 70928 32780
rect 70974 32734 71000 32780
tri 25247 32558 25382 32693 ne
rect 25382 32680 25523 32693
rect 25382 32634 25398 32680
rect 25444 32634 25523 32680
rect 25382 32558 25523 32634
tri 25382 32417 25523 32558 ne
tri 25523 32553 25663 32693 sw
rect 70802 32676 71000 32734
rect 70802 32630 70824 32676
rect 70870 32630 70928 32676
rect 70974 32630 71000 32676
rect 70802 32572 71000 32630
rect 25523 32548 25663 32553
rect 25523 32502 25530 32548
rect 25576 32502 25663 32548
rect 25523 32417 25663 32502
tri 25663 32417 25799 32553 sw
rect 70802 32526 70824 32572
rect 70870 32526 70928 32572
rect 70974 32526 71000 32572
rect 70802 32468 71000 32526
rect 70802 32422 70824 32468
rect 70870 32422 70928 32468
rect 70974 32422 71000 32468
tri 25523 32293 25647 32417 ne
rect 25647 32416 25799 32417
rect 25647 32370 25662 32416
rect 25708 32370 25799 32416
rect 25647 32327 25799 32370
tri 25799 32327 25889 32417 sw
rect 70802 32364 71000 32422
rect 25647 32293 25889 32327
tri 25647 32146 25794 32293 ne
rect 25794 32284 25889 32293
rect 25840 32238 25889 32284
rect 25794 32186 25889 32238
tri 25889 32186 26030 32327 sw
rect 70802 32318 70824 32364
rect 70870 32318 70928 32364
rect 70974 32318 71000 32364
rect 70802 32260 71000 32318
rect 70802 32214 70824 32260
rect 70870 32214 70928 32260
rect 70974 32214 71000 32260
rect 25794 32152 26030 32186
rect 25794 32146 25926 32152
tri 25794 32018 25922 32146 ne
rect 25922 32106 25926 32146
rect 25972 32106 26030 32152
rect 25922 32052 26030 32106
tri 26030 32052 26164 32186 sw
rect 70802 32156 71000 32214
rect 70802 32110 70824 32156
rect 70870 32110 70928 32156
rect 70974 32110 71000 32156
rect 70802 32052 71000 32110
rect 25922 32020 26164 32052
rect 25922 32018 26058 32020
tri 25922 31882 26058 32018 ne
rect 26104 31974 26164 32020
rect 26058 31910 26164 31974
tri 26164 31910 26306 32052 sw
rect 70802 32006 70824 32052
rect 70870 32006 70928 32052
rect 70974 32006 71000 32052
rect 70802 31948 71000 32006
rect 26058 31888 26306 31910
rect 26058 31882 26190 31888
tri 26058 31775 26165 31882 ne
rect 26165 31842 26190 31882
rect 26236 31842 26306 31888
rect 26165 31776 26306 31842
tri 26306 31776 26440 31910 sw
rect 70802 31902 70824 31948
rect 70870 31902 70928 31948
rect 70974 31902 71000 31948
rect 70802 31844 71000 31902
rect 70802 31798 70824 31844
rect 70870 31798 70928 31844
rect 70974 31798 71000 31844
rect 26165 31775 26440 31776
tri 26165 31618 26322 31775 ne
rect 26322 31756 26440 31775
rect 26368 31710 26440 31756
rect 26322 31634 26440 31710
tri 26440 31634 26582 31776 sw
rect 70802 31740 71000 31798
rect 70802 31694 70824 31740
rect 70870 31694 70928 31740
rect 70974 31694 71000 31740
rect 70802 31636 71000 31694
rect 26322 31624 26582 31634
rect 26322 31618 26454 31624
tri 26322 31499 26441 31618 ne
rect 26441 31578 26454 31618
rect 26500 31578 26582 31624
rect 26441 31499 26582 31578
tri 26582 31499 26717 31634 sw
rect 70802 31590 70824 31636
rect 70870 31590 70928 31636
rect 70974 31590 71000 31636
rect 70802 31532 71000 31590
tri 26441 31354 26586 31499 ne
rect 26586 31492 26717 31499
rect 26632 31446 26717 31492
rect 26586 31365 26717 31446
tri 26717 31365 26851 31499 sw
rect 70802 31486 70824 31532
rect 70870 31486 70928 31532
rect 70974 31486 71000 31532
rect 70802 31428 71000 31486
rect 70802 31382 70824 31428
rect 70870 31382 70928 31428
rect 70974 31382 71000 31428
rect 26586 31360 26851 31365
rect 26586 31354 26718 31360
tri 26586 31243 26697 31354 ne
rect 26697 31314 26718 31354
rect 26764 31314 26851 31360
rect 26697 31268 26851 31314
tri 26851 31268 26948 31365 sw
rect 70802 31324 71000 31382
rect 70802 31278 70824 31324
rect 70870 31278 70928 31324
rect 70974 31278 71000 31324
rect 26697 31243 26948 31268
tri 26697 31090 26850 31243 ne
rect 26850 31228 26948 31243
rect 26896 31182 26948 31228
rect 26850 31127 26948 31182
tri 26948 31127 27089 31268 sw
rect 70802 31220 71000 31278
rect 70802 31174 70824 31220
rect 70870 31174 70928 31220
rect 70974 31174 71000 31220
rect 26850 31096 27089 31127
rect 26850 31090 26982 31096
tri 26850 30999 26941 31090 ne
rect 26941 31050 26982 31090
rect 27028 31050 27089 31096
rect 26941 30999 27089 31050
tri 27089 30999 27217 31127 sw
rect 70802 31116 71000 31174
rect 70802 31070 70824 31116
rect 70870 31070 70928 31116
rect 70974 31070 71000 31116
rect 70802 31012 71000 31070
tri 26941 30826 27114 30999 ne
rect 27114 30964 27217 30999
rect 27160 30918 27217 30964
rect 27114 30851 27217 30918
tri 27217 30851 27365 30999 sw
rect 70802 30966 70824 31012
rect 70870 30966 70928 31012
rect 70974 30966 71000 31012
rect 70802 30908 71000 30966
rect 70802 30862 70824 30908
rect 70870 30862 70928 30908
rect 70974 30862 71000 30908
rect 27114 30832 27365 30851
rect 27114 30826 27246 30832
tri 27114 30716 27224 30826 ne
rect 27224 30786 27246 30826
rect 27292 30786 27365 30832
rect 27224 30716 27365 30786
tri 27365 30716 27500 30851 sw
rect 70802 30804 71000 30862
rect 70802 30758 70824 30804
rect 70870 30758 70928 30804
rect 70974 30758 71000 30804
tri 27224 30562 27378 30716 ne
rect 27378 30700 27500 30716
rect 27424 30654 27500 30700
rect 27378 30588 27500 30654
tri 27500 30588 27628 30716 sw
rect 70802 30700 71000 30758
rect 70802 30654 70824 30700
rect 70870 30654 70928 30700
rect 70974 30654 71000 30700
rect 70802 30596 71000 30654
rect 27378 30568 27628 30588
rect 27378 30562 27510 30568
tri 27378 30440 27500 30562 ne
rect 27500 30522 27510 30562
rect 27556 30522 27628 30568
rect 27500 30440 27628 30522
tri 27628 30440 27776 30588 sw
rect 70802 30550 70824 30596
rect 70870 30550 70928 30596
rect 70974 30550 71000 30596
rect 70802 30492 71000 30550
rect 70802 30446 70824 30492
rect 70870 30446 70928 30492
rect 70974 30446 71000 30492
tri 27500 30298 27642 30440 ne
rect 27642 30436 27776 30440
rect 27688 30390 27776 30436
rect 27642 30312 27776 30390
tri 27776 30312 27904 30440 sw
rect 70802 30388 71000 30446
rect 70802 30342 70824 30388
rect 70870 30342 70928 30388
rect 70974 30342 71000 30388
rect 27642 30304 27904 30312
rect 27642 30298 27774 30304
tri 27642 30209 27731 30298 ne
rect 27731 30258 27774 30298
rect 27820 30258 27904 30304
rect 27731 30209 27904 30258
tri 27904 30209 28007 30312 sw
rect 70802 30284 71000 30342
rect 70802 30238 70824 30284
rect 70870 30238 70928 30284
rect 70974 30238 71000 30284
tri 27731 30059 27881 30209 ne
rect 27881 30172 28007 30209
rect 27881 30126 27906 30172
rect 27952 30126 28007 30172
rect 27881 30068 28007 30126
tri 28007 30068 28148 30209 sw
rect 70802 30180 71000 30238
rect 70802 30134 70824 30180
rect 70870 30134 70928 30180
rect 70974 30134 71000 30180
rect 70802 30076 71000 30134
rect 27881 30059 28148 30068
tri 27881 29933 28007 30059 ne
rect 28007 30040 28148 30059
rect 28007 29994 28038 30040
rect 28084 29994 28148 30040
rect 28007 29933 28148 29994
tri 28148 29933 28283 30068 sw
rect 70802 30030 70824 30076
rect 70870 30030 70928 30076
rect 70974 30030 71000 30076
rect 70802 29972 71000 30030
tri 28007 29784 28156 29933 ne
rect 28156 29908 28283 29933
rect 28156 29862 28170 29908
rect 28216 29862 28283 29908
rect 28156 29811 28283 29862
tri 28283 29811 28405 29933 sw
rect 70802 29926 70824 29972
rect 70870 29926 70928 29972
rect 70974 29926 71000 29972
rect 70802 29868 71000 29926
rect 70802 29822 70824 29868
rect 70870 29822 70928 29868
rect 70974 29822 71000 29868
rect 28156 29784 28405 29811
tri 28156 29657 28283 29784 ne
rect 28283 29776 28405 29784
rect 28283 29730 28302 29776
rect 28348 29730 28405 29776
rect 28283 29657 28405 29730
tri 28405 29657 28559 29811 sw
rect 70802 29764 71000 29822
rect 70802 29718 70824 29764
rect 70870 29718 70928 29764
rect 70974 29718 71000 29764
rect 70802 29660 71000 29718
tri 28283 29535 28405 29657 ne
rect 28405 29644 28559 29657
rect 28405 29598 28434 29644
rect 28480 29598 28559 29644
rect 28405 29535 28559 29598
tri 28559 29535 28681 29657 sw
rect 70802 29614 70824 29660
rect 70870 29614 70928 29660
rect 70974 29614 71000 29660
rect 70802 29556 71000 29614
tri 28405 29381 28559 29535 ne
rect 28559 29512 28681 29535
rect 28559 29466 28566 29512
rect 28612 29466 28681 29512
rect 28559 29381 28681 29466
tri 28681 29381 28835 29535 sw
rect 70802 29510 70824 29556
rect 70870 29510 70928 29556
rect 70974 29510 71000 29556
rect 70802 29452 71000 29510
rect 70802 29406 70824 29452
rect 70870 29406 70928 29452
rect 70974 29406 71000 29452
tri 28559 29246 28694 29381 ne
rect 28694 29380 28835 29381
rect 28694 29334 28698 29380
rect 28744 29334 28835 29380
rect 28694 29259 28835 29334
tri 28835 29259 28957 29381 sw
rect 70802 29348 71000 29406
rect 70802 29302 70824 29348
rect 70870 29302 70928 29348
rect 70974 29302 71000 29348
rect 28694 29248 28957 29259
rect 28694 29246 28830 29248
tri 28694 29110 28830 29246 ne
rect 28876 29202 28957 29248
rect 28830 29124 28957 29202
tri 28957 29124 29092 29259 sw
rect 70802 29244 71000 29302
rect 70802 29198 70824 29244
rect 70870 29198 70928 29244
rect 70974 29198 71000 29244
rect 70802 29140 71000 29198
rect 28830 29116 29092 29124
rect 28830 29110 28962 29116
tri 28830 29009 28931 29110 ne
rect 28931 29070 28962 29110
rect 29008 29070 29092 29116
rect 28931 29015 29092 29070
tri 29092 29015 29201 29124 sw
rect 70802 29094 70824 29140
rect 70870 29094 70928 29140
rect 70974 29094 71000 29140
rect 70802 29036 71000 29094
rect 28931 29009 29201 29015
tri 28931 28846 29094 29009 ne
rect 29094 28984 29201 29009
rect 29140 28938 29201 28984
rect 29094 28874 29201 28938
tri 29201 28874 29342 29015 sw
rect 70802 28990 70824 29036
rect 70870 28990 70928 29036
rect 70974 28990 71000 29036
rect 70802 28932 71000 28990
rect 70802 28886 70824 28932
rect 70870 28886 70928 28932
rect 70974 28886 71000 28932
rect 29094 28852 29342 28874
rect 29094 28846 29226 28852
tri 29094 28735 29205 28846 ne
rect 29205 28806 29226 28846
rect 29272 28806 29342 28852
rect 29205 28758 29342 28806
tri 29342 28758 29458 28874 sw
rect 70802 28828 71000 28886
rect 70802 28782 70824 28828
rect 70870 28782 70928 28828
rect 70974 28782 71000 28828
rect 29205 28735 29458 28758
tri 29205 28582 29358 28735 ne
rect 29358 28720 29458 28735
rect 29404 28674 29458 28720
rect 29358 28598 29458 28674
tri 29458 28598 29618 28758 sw
rect 70802 28724 71000 28782
rect 70802 28678 70824 28724
rect 70870 28678 70928 28724
rect 70974 28678 71000 28724
rect 70802 28620 71000 28678
rect 29358 28588 29618 28598
rect 29358 28582 29490 28588
tri 29358 28463 29477 28582 ne
rect 29477 28542 29490 28582
rect 29536 28542 29618 28588
rect 29477 28482 29618 28542
tri 29618 28482 29734 28598 sw
rect 70802 28574 70824 28620
rect 70870 28574 70928 28620
rect 70974 28574 71000 28620
rect 70802 28516 71000 28574
rect 29477 28463 29734 28482
tri 29477 28318 29622 28463 ne
rect 29622 28456 29734 28463
rect 29668 28410 29734 28456
rect 29622 28347 29734 28410
tri 29734 28347 29869 28482 sw
rect 70802 28470 70824 28516
rect 70870 28470 70928 28516
rect 70974 28470 71000 28516
rect 70802 28412 71000 28470
rect 70802 28366 70824 28412
rect 70870 28366 70928 28412
rect 70974 28366 71000 28412
rect 29622 28324 29869 28347
rect 29622 28318 29754 28324
tri 29622 28187 29753 28318 ne
rect 29753 28278 29754 28318
rect 29800 28278 29869 28324
rect 29753 28232 29869 28278
tri 29869 28232 29984 28347 sw
rect 70802 28308 71000 28366
rect 70802 28262 70824 28308
rect 70870 28262 70928 28308
rect 70974 28262 71000 28308
rect 29753 28192 29984 28232
rect 29753 28187 29886 28192
tri 29753 28054 29886 28187 ne
rect 29932 28146 29984 28192
rect 29886 28071 29984 28146
tri 29984 28071 30145 28232 sw
rect 70802 28204 71000 28262
rect 70802 28158 70824 28204
rect 70870 28158 70928 28204
rect 70974 28158 71000 28204
rect 70802 28100 71000 28158
rect 29886 28060 30145 28071
rect 29886 28054 30018 28060
tri 29886 27960 29980 28054 ne
rect 29980 28014 30018 28054
rect 30064 28014 30145 28060
rect 29980 27960 30145 28014
tri 29980 27795 30145 27960 ne
tri 30145 27956 30260 28071 sw
rect 70802 28054 70824 28100
rect 70870 28054 70928 28100
rect 70974 28054 71000 28100
rect 70802 27996 71000 28054
rect 30145 27928 30260 27956
rect 30145 27882 30150 27928
rect 30196 27882 30260 27928
rect 30145 27815 30260 27882
tri 30260 27815 30401 27956 sw
rect 70802 27950 70824 27996
rect 70870 27950 70928 27996
rect 70974 27950 71000 27996
rect 70802 27892 71000 27950
rect 70802 27846 70824 27892
rect 70870 27846 70928 27892
rect 70974 27846 71000 27892
rect 30145 27796 30401 27815
rect 30145 27795 30282 27796
tri 30145 27660 30280 27795 ne
rect 30280 27750 30282 27795
rect 30328 27750 30401 27796
rect 30280 27705 30401 27750
tri 30401 27705 30511 27815 sw
rect 70802 27788 71000 27846
rect 70802 27742 70824 27788
rect 70870 27742 70928 27788
rect 70974 27742 71000 27788
rect 30280 27664 30511 27705
rect 30280 27660 30414 27664
tri 30280 27526 30414 27660 ne
rect 30460 27618 30511 27664
rect 30414 27539 30511 27618
tri 30511 27539 30677 27705 sw
rect 70802 27684 71000 27742
rect 70802 27638 70824 27684
rect 70870 27638 70928 27684
rect 70974 27638 71000 27684
rect 70802 27580 71000 27638
rect 30414 27532 30677 27539
rect 30414 27526 30546 27532
tri 30414 27404 30536 27526 ne
rect 30536 27486 30546 27526
rect 30592 27486 30677 27532
rect 30536 27404 30677 27486
tri 30677 27404 30812 27539 sw
rect 70802 27534 70824 27580
rect 70870 27534 70928 27580
rect 70974 27534 71000 27580
rect 70802 27476 71000 27534
rect 70802 27430 70824 27476
rect 70870 27430 70928 27476
rect 70974 27430 71000 27476
tri 30536 27262 30678 27404 ne
rect 30678 27400 30812 27404
rect 30724 27354 30812 27400
rect 30678 27294 30812 27354
tri 30812 27294 30922 27404 sw
rect 70802 27372 71000 27430
rect 70802 27326 70824 27372
rect 70870 27326 70928 27372
rect 70974 27326 71000 27372
rect 30678 27268 30922 27294
rect 30678 27262 30810 27268
tri 30678 27173 30767 27262 ne
rect 30767 27222 30810 27262
rect 30856 27222 30922 27268
rect 30767 27173 30922 27222
tri 30922 27173 31043 27294 sw
rect 70802 27268 71000 27326
rect 70802 27222 70824 27268
rect 70870 27222 70928 27268
rect 70974 27222 71000 27268
tri 30767 26998 30942 27173 ne
rect 30942 27136 31043 27173
rect 30988 27090 31043 27136
rect 30942 27018 31043 27090
tri 31043 27018 31198 27173 sw
rect 70802 27164 71000 27222
rect 70802 27118 70824 27164
rect 70870 27118 70928 27164
rect 70974 27118 71000 27164
rect 70802 27060 71000 27118
rect 30942 27004 31198 27018
rect 30942 26998 31074 27004
tri 30942 26866 31074 26998 ne
rect 31120 26958 31198 27004
rect 31074 26897 31198 26958
tri 31198 26897 31319 27018 sw
rect 70802 27014 70824 27060
rect 70870 27014 70928 27060
rect 70974 27014 71000 27060
rect 70802 26956 71000 27014
rect 70802 26910 70824 26956
rect 70870 26910 70928 26956
rect 70974 26910 71000 26956
rect 31074 26872 31319 26897
rect 31074 26866 31206 26872
tri 31074 26734 31206 26866 ne
rect 31252 26826 31319 26872
rect 31206 26756 31319 26826
tri 31319 26756 31460 26897 sw
rect 70802 26852 71000 26910
rect 70802 26806 70824 26852
rect 70870 26806 70928 26852
rect 70974 26806 71000 26852
rect 31206 26740 31460 26756
rect 31206 26734 31338 26740
tri 31206 26607 31333 26734 ne
rect 31333 26694 31338 26734
rect 31384 26694 31460 26740
rect 31333 26621 31460 26694
tri 31460 26621 31595 26756 sw
rect 70802 26748 71000 26806
rect 70802 26702 70824 26748
rect 70870 26702 70928 26748
rect 70974 26702 71000 26748
rect 70802 26644 71000 26702
rect 31333 26608 31595 26621
rect 31333 26607 31470 26608
tri 31333 26501 31439 26607 ne
rect 31439 26562 31470 26607
rect 31516 26562 31595 26608
rect 31439 26517 31595 26562
tri 31595 26517 31699 26621 sw
rect 70802 26598 70824 26644
rect 70870 26598 70928 26644
rect 70974 26598 71000 26644
rect 70802 26540 71000 26598
rect 31439 26501 31699 26517
tri 31439 26345 31595 26501 ne
rect 31595 26476 31699 26501
rect 31595 26430 31602 26476
rect 31648 26430 31699 26476
rect 31595 26345 31699 26430
tri 31699 26345 31871 26517 sw
rect 70802 26494 70824 26540
rect 70870 26494 70928 26540
rect 70974 26494 71000 26540
rect 70802 26436 71000 26494
rect 70802 26390 70824 26436
rect 70870 26390 70928 26436
rect 70974 26390 71000 26436
tri 31595 26241 31699 26345 ne
rect 31699 26344 31871 26345
rect 31699 26298 31734 26344
rect 31780 26298 31871 26344
rect 31699 26241 31871 26298
tri 31871 26241 31975 26345 sw
rect 70802 26332 71000 26390
rect 70802 26286 70824 26332
rect 70870 26286 70928 26332
rect 70974 26286 71000 26332
tri 31699 26074 31866 26241 ne
rect 31866 26212 31975 26241
rect 31912 26166 31975 26212
rect 31866 26114 31975 26166
tri 31975 26114 32102 26241 sw
rect 70802 26228 71000 26286
rect 70802 26182 70824 26228
rect 70870 26182 70928 26228
rect 70974 26182 71000 26228
rect 70802 26124 71000 26182
rect 31866 26080 32102 26114
rect 31866 26074 31998 26080
tri 31866 25979 31961 26074 ne
rect 31961 26034 31998 26074
rect 32044 26034 32102 26080
rect 31961 25979 32102 26034
tri 31961 25838 32102 25979 ne
tri 32102 25965 32251 26114 sw
rect 70802 26078 70824 26124
rect 70870 26078 70928 26124
rect 70974 26078 71000 26124
rect 70802 26020 71000 26078
rect 70802 25974 70824 26020
rect 70870 25974 70928 26020
rect 70974 25974 71000 26020
rect 32102 25948 32251 25965
rect 32102 25902 32130 25948
rect 32176 25902 32251 25948
rect 32102 25838 32251 25902
tri 32102 25726 32214 25838 ne
rect 32214 25830 32251 25838
tri 32251 25830 32386 25965 sw
rect 70802 25916 71000 25974
rect 70802 25870 70824 25916
rect 70870 25870 70928 25916
rect 70974 25870 71000 25916
rect 32214 25816 32386 25830
rect 32214 25770 32262 25816
rect 32308 25770 32386 25816
rect 32214 25726 32386 25770
tri 32214 25554 32386 25726 ne
tri 32386 25703 32513 25830 sw
rect 70802 25812 71000 25870
rect 70802 25766 70824 25812
rect 70870 25766 70928 25812
rect 70974 25766 71000 25812
rect 70802 25708 71000 25766
rect 32386 25684 32513 25703
rect 32386 25638 32394 25684
rect 32440 25638 32513 25684
rect 32386 25562 32513 25638
tri 32513 25562 32654 25703 sw
rect 70802 25662 70824 25708
rect 70870 25662 70928 25708
rect 70974 25662 71000 25708
rect 70802 25604 71000 25662
rect 32386 25554 32654 25562
tri 32386 25451 32489 25554 ne
rect 32489 25552 32654 25554
rect 32489 25506 32526 25552
rect 32572 25506 32654 25552
rect 32489 25464 32654 25506
tri 32654 25464 32752 25562 sw
rect 70802 25558 70824 25604
rect 70870 25558 70928 25604
rect 70974 25558 71000 25604
rect 70802 25500 71000 25558
rect 32489 25451 32752 25464
tri 32489 25282 32658 25451 ne
rect 32658 25420 32752 25451
rect 32704 25374 32752 25420
rect 32658 25331 32752 25374
tri 32752 25331 32885 25464 sw
rect 70802 25454 70824 25500
rect 70870 25454 70928 25500
rect 70974 25454 71000 25500
rect 70802 25396 71000 25454
rect 70802 25350 70824 25396
rect 70870 25350 70928 25396
rect 70974 25350 71000 25396
rect 32658 25288 32885 25331
rect 32658 25282 32790 25288
tri 32658 25151 32789 25282 ne
rect 32789 25242 32790 25282
rect 32836 25242 32885 25288
rect 32789 25188 32885 25242
tri 32885 25188 33028 25331 sw
rect 70802 25292 71000 25350
rect 70802 25246 70824 25292
rect 70870 25246 70928 25292
rect 70974 25246 71000 25292
rect 70802 25188 71000 25246
rect 32789 25156 33028 25188
rect 32789 25151 32922 25156
tri 32789 25018 32922 25151 ne
rect 32968 25110 33028 25156
rect 32922 25053 33028 25110
tri 33028 25053 33163 25188 sw
rect 70802 25142 70824 25188
rect 70870 25142 70928 25188
rect 70974 25142 71000 25188
rect 70802 25084 71000 25142
rect 32922 25024 33163 25053
rect 32922 25018 33054 25024
tri 32922 24920 33020 25018 ne
rect 33020 24978 33054 25018
rect 33100 24978 33163 25024
rect 33020 24920 33163 24978
tri 33163 24920 33296 25053 sw
rect 70802 25038 70824 25084
rect 70870 25038 70928 25084
rect 70974 25038 71000 25084
rect 70802 24980 71000 25038
rect 70802 24934 70824 24980
rect 70870 24934 70928 24980
rect 70974 24934 71000 24980
tri 33020 24754 33186 24920 ne
rect 33186 24892 33296 24920
rect 33232 24846 33296 24892
rect 33186 24777 33296 24846
tri 33296 24777 33439 24920 sw
rect 70802 24876 71000 24934
rect 70802 24830 70824 24876
rect 70870 24830 70928 24876
rect 70974 24830 71000 24876
rect 33186 24760 33439 24777
rect 33186 24754 33318 24760
tri 33186 24632 33308 24754 ne
rect 33308 24714 33318 24754
rect 33364 24714 33439 24760
rect 33308 24644 33439 24714
tri 33439 24644 33572 24777 sw
rect 70802 24772 71000 24830
rect 70802 24726 70824 24772
rect 70870 24726 70928 24772
rect 70974 24726 71000 24772
rect 70802 24668 71000 24726
rect 33308 24632 33572 24644
tri 33308 24490 33450 24632 ne
rect 33450 24628 33572 24632
rect 33496 24582 33572 24628
rect 33450 24503 33572 24582
tri 33572 24503 33713 24644 sw
rect 70802 24622 70824 24668
rect 70870 24622 70928 24668
rect 70974 24622 71000 24668
rect 70802 24564 71000 24622
rect 70802 24518 70824 24564
rect 70870 24518 70928 24564
rect 70974 24518 71000 24564
rect 33450 24496 33713 24503
rect 33450 24490 33582 24496
tri 33450 24366 33574 24490 ne
rect 33574 24450 33582 24490
rect 33628 24450 33713 24496
rect 33574 24366 33713 24450
tri 33713 24366 33850 24503 sw
rect 70802 24460 71000 24518
rect 70802 24414 70824 24460
rect 70870 24414 70928 24460
rect 70974 24414 71000 24460
tri 33574 24226 33714 24366 ne
rect 33714 24364 33850 24366
rect 33760 24318 33850 24364
rect 33714 24272 33850 24318
tri 33850 24272 33944 24366 sw
rect 70802 24356 71000 24414
rect 70802 24310 70824 24356
rect 70870 24310 70928 24356
rect 70974 24310 71000 24356
rect 33714 24232 33944 24272
rect 33714 24226 33846 24232
tri 33714 24137 33803 24226 ne
rect 33803 24186 33846 24226
rect 33892 24186 33944 24232
rect 33803 24137 33944 24186
tri 33944 24137 34079 24272 sw
rect 70802 24252 71000 24310
rect 70802 24206 70824 24252
rect 70870 24206 70928 24252
rect 70974 24206 71000 24252
rect 70802 24148 71000 24206
tri 33803 23962 33978 24137 ne
rect 33978 24100 34079 24137
rect 34024 24054 34079 24100
rect 33978 24000 34079 24054
tri 34079 24000 34216 24137 sw
rect 70802 24102 70824 24148
rect 70870 24102 70928 24148
rect 70974 24102 71000 24148
rect 70802 24044 71000 24102
rect 33978 23968 34216 24000
rect 33978 23962 34110 23968
tri 33978 23861 34079 23962 ne
rect 34079 23922 34110 23962
rect 34156 23922 34216 23968
rect 34079 23861 34216 23922
tri 34216 23861 34355 24000 sw
rect 70802 23998 70824 24044
rect 70870 23998 70928 24044
rect 70974 23998 71000 24044
rect 70802 23940 71000 23998
rect 70802 23894 70824 23940
rect 70870 23894 70928 23940
rect 70974 23894 71000 23940
tri 34079 23698 34242 23861 ne
rect 34242 23836 34355 23861
rect 34288 23790 34355 23836
rect 34242 23724 34355 23790
tri 34355 23724 34492 23861 sw
rect 70802 23836 71000 23894
rect 70802 23790 70824 23836
rect 70870 23790 70928 23836
rect 70974 23790 71000 23836
rect 70802 23732 71000 23790
rect 34242 23704 34492 23724
rect 34242 23698 34374 23704
tri 34242 23582 34358 23698 ne
rect 34358 23658 34374 23698
rect 34420 23658 34492 23704
rect 34358 23585 34492 23658
tri 34492 23585 34631 23724 sw
rect 70802 23686 70824 23732
rect 70870 23686 70928 23732
rect 70974 23686 71000 23732
rect 70802 23628 71000 23686
rect 34358 23582 34631 23585
tri 34358 23434 34506 23582 ne
rect 34506 23572 34631 23582
rect 34552 23526 34631 23572
rect 34506 23448 34631 23526
tri 34631 23448 34768 23585 sw
rect 70802 23582 70824 23628
rect 70870 23582 70928 23628
rect 70974 23582 71000 23628
rect 70802 23524 71000 23582
rect 70802 23478 70824 23524
rect 70870 23478 70928 23524
rect 70974 23478 71000 23524
rect 34506 23440 34768 23448
rect 34506 23434 34638 23440
tri 34506 23309 34631 23434 ne
rect 34631 23394 34638 23434
rect 34684 23394 34768 23440
rect 34631 23309 34768 23394
tri 34768 23309 34907 23448 sw
rect 70802 23420 71000 23478
rect 70802 23374 70824 23420
rect 70870 23374 70928 23420
rect 70974 23374 71000 23420
rect 70802 23316 71000 23374
tri 34631 23173 34767 23309 ne
rect 34767 23308 34907 23309
rect 34767 23262 34770 23308
rect 34816 23262 34907 23308
rect 34767 23178 34907 23262
tri 34907 23178 35038 23309 sw
rect 70802 23270 70824 23316
rect 70870 23270 70928 23316
rect 70974 23270 71000 23316
rect 70802 23212 71000 23270
rect 34767 23176 35038 23178
rect 34767 23173 34902 23176
tri 34767 23038 34902 23173 ne
rect 34948 23130 35038 23176
rect 34902 23078 35038 23130
tri 35038 23078 35138 23178 sw
rect 70802 23166 70824 23212
rect 70870 23166 70928 23212
rect 70974 23166 71000 23212
rect 70802 23108 71000 23166
rect 34902 23044 35138 23078
rect 34902 23038 35034 23044
tri 34902 22947 34993 23038 ne
rect 34993 22998 35034 23038
rect 35080 22998 35138 23044
rect 34993 22947 35138 22998
tri 35138 22947 35269 23078 sw
rect 70802 23062 70824 23108
rect 70870 23062 70928 23108
rect 70974 23062 71000 23108
rect 70802 23004 71000 23062
rect 70802 22958 70824 23004
rect 70870 22958 70928 23004
rect 70974 22958 71000 23004
tri 34993 22774 35166 22947 ne
rect 35166 22912 35269 22947
rect 35212 22866 35269 22912
rect 35166 22802 35269 22866
tri 35269 22802 35414 22947 sw
rect 70802 22900 71000 22958
rect 70802 22854 70824 22900
rect 70870 22854 70928 22900
rect 70974 22854 71000 22900
rect 35166 22780 35414 22802
rect 35166 22774 35298 22780
tri 35166 22667 35273 22774 ne
rect 35273 22734 35298 22774
rect 35344 22734 35414 22780
rect 35273 22671 35414 22734
tri 35414 22671 35545 22802 sw
rect 70802 22796 71000 22854
rect 70802 22750 70824 22796
rect 70870 22750 70928 22796
rect 70974 22750 71000 22796
rect 70802 22692 71000 22750
rect 35273 22667 35545 22671
tri 35273 22510 35430 22667 ne
rect 35430 22648 35545 22667
rect 35476 22602 35545 22648
rect 35430 22526 35545 22602
tri 35545 22526 35690 22671 sw
rect 70802 22646 70824 22692
rect 70870 22646 70928 22692
rect 70974 22646 71000 22692
rect 70802 22588 71000 22646
rect 70802 22542 70824 22588
rect 70870 22542 70928 22588
rect 70974 22542 71000 22588
rect 35430 22516 35690 22526
rect 35430 22510 35562 22516
tri 35430 22391 35549 22510 ne
rect 35549 22470 35562 22510
rect 35608 22470 35690 22516
rect 35549 22391 35690 22470
tri 35690 22391 35825 22526 sw
rect 70802 22484 71000 22542
rect 70802 22438 70824 22484
rect 70870 22438 70928 22484
rect 70974 22438 71000 22484
tri 35549 22246 35694 22391 ne
rect 35694 22384 35825 22391
rect 35740 22338 35825 22384
rect 35694 22260 35825 22338
tri 35825 22260 35956 22391 sw
rect 70802 22380 71000 22438
rect 70802 22334 70824 22380
rect 70870 22334 70928 22380
rect 70974 22334 71000 22380
rect 70802 22276 71000 22334
rect 35694 22252 35956 22260
rect 35694 22246 35826 22252
tri 35694 22123 35817 22246 ne
rect 35817 22206 35826 22246
rect 35872 22206 35956 22252
rect 35817 22125 35956 22206
tri 35956 22125 36091 22260 sw
rect 70802 22230 70824 22276
rect 70870 22230 70928 22276
rect 70974 22230 71000 22276
rect 70802 22172 71000 22230
rect 70802 22126 70824 22172
rect 70870 22126 70928 22172
rect 70974 22126 71000 22172
rect 35817 22123 36091 22125
tri 35817 21982 35958 22123 ne
rect 35958 22120 36091 22123
rect 36004 22074 36091 22120
rect 35958 22019 36091 22074
tri 36091 22019 36197 22125 sw
rect 70802 22068 71000 22126
rect 70802 22022 70824 22068
rect 70870 22022 70928 22068
rect 70974 22022 71000 22068
rect 35958 21988 36197 22019
rect 35958 21982 36090 21988
tri 35958 21884 36056 21982 ne
rect 36056 21942 36090 21982
rect 36136 21942 36197 21988
rect 36056 21894 36197 21942
tri 36197 21894 36322 22019 sw
rect 70802 21964 71000 22022
rect 70802 21918 70824 21964
rect 70870 21918 70928 21964
rect 70974 21918 71000 21964
rect 36056 21884 36322 21894
tri 36056 21718 36222 21884 ne
rect 36222 21856 36322 21884
rect 36268 21810 36322 21856
rect 36222 21743 36322 21810
tri 36322 21743 36473 21894 sw
rect 70802 21860 71000 21918
rect 70802 21814 70824 21860
rect 70870 21814 70928 21860
rect 70974 21814 71000 21860
rect 70802 21756 71000 21814
rect 36222 21724 36473 21743
rect 36222 21718 36354 21724
tri 36222 21608 36332 21718 ne
rect 36332 21678 36354 21718
rect 36400 21678 36473 21724
rect 36332 21608 36473 21678
tri 36473 21608 36608 21743 sw
rect 70802 21710 70824 21756
rect 70870 21710 70928 21756
rect 70974 21710 71000 21756
rect 70802 21652 71000 21710
tri 36332 21454 36486 21608 ne
rect 36486 21592 36608 21608
rect 36532 21546 36608 21592
rect 36486 21483 36608 21546
tri 36608 21483 36733 21608 sw
rect 70802 21606 70824 21652
rect 70870 21606 70928 21652
rect 70974 21606 71000 21652
rect 70802 21548 71000 21606
rect 70802 21502 70824 21548
rect 70870 21502 70928 21548
rect 70974 21502 71000 21548
rect 36486 21460 36733 21483
rect 36486 21454 36618 21460
tri 36486 21332 36608 21454 ne
rect 36608 21414 36618 21454
rect 36664 21414 36733 21460
rect 36608 21332 36733 21414
tri 36733 21332 36884 21483 sw
rect 70802 21444 71000 21502
rect 70802 21398 70824 21444
rect 70870 21398 70928 21444
rect 70974 21398 71000 21444
rect 70802 21340 71000 21398
tri 36608 21190 36750 21332 ne
rect 36750 21328 36884 21332
rect 36796 21282 36884 21328
rect 36750 21207 36884 21282
tri 36884 21207 37009 21332 sw
rect 70802 21294 70824 21340
rect 70870 21294 70928 21340
rect 70974 21294 71000 21340
rect 70802 21236 71000 21294
rect 36750 21196 37009 21207
rect 36750 21190 36882 21196
tri 36750 21101 36839 21190 ne
rect 36839 21150 36882 21190
rect 36928 21150 37009 21196
rect 36839 21101 37009 21150
tri 36839 20931 37009 21101 ne
tri 37009 21072 37144 21207 sw
rect 70802 21190 70824 21236
rect 70870 21190 70928 21236
rect 70974 21190 71000 21236
rect 70802 21132 71000 21190
rect 70802 21086 70824 21132
rect 70870 21086 70928 21132
rect 70974 21086 71000 21132
rect 37009 21064 37144 21072
rect 37009 21018 37014 21064
rect 37060 21018 37144 21064
rect 37009 20960 37144 21018
tri 37144 20960 37256 21072 sw
rect 70802 21028 71000 21086
rect 70802 20982 70824 21028
rect 70870 20982 70928 21028
rect 70974 20982 71000 21028
rect 37009 20932 37256 20960
rect 37009 20931 37146 20932
tri 37009 20796 37144 20931 ne
rect 37144 20886 37146 20931
rect 37192 20886 37256 20932
rect 37144 20825 37256 20886
tri 37256 20825 37391 20960 sw
rect 70802 20924 71000 20982
rect 70802 20878 70824 20924
rect 70870 20878 70928 20924
rect 70974 20878 71000 20924
rect 37144 20800 37391 20825
rect 37144 20796 37278 20800
tri 37144 20662 37278 20796 ne
rect 37324 20754 37391 20800
rect 37278 20706 37391 20754
tri 37391 20706 37510 20825 sw
rect 70802 20820 71000 20878
rect 70802 20774 70824 20820
rect 70870 20774 70928 20820
rect 70974 20774 71000 20820
rect 70802 20716 71000 20774
rect 37278 20668 37510 20706
rect 37278 20662 37410 20668
tri 37278 20549 37391 20662 ne
rect 37391 20622 37410 20662
rect 37456 20622 37510 20668
rect 37391 20549 37510 20622
tri 37510 20549 37667 20706 sw
rect 70802 20670 70824 20716
rect 70870 20670 70928 20716
rect 70974 20670 71000 20716
rect 70802 20612 71000 20670
rect 70802 20566 70824 20612
rect 70870 20566 70928 20612
rect 70974 20566 71000 20612
tri 37391 20398 37542 20549 ne
rect 37542 20536 37667 20549
rect 37588 20490 37667 20536
rect 37542 20430 37667 20490
tri 37667 20430 37786 20549 sw
rect 70802 20508 71000 20566
rect 70802 20462 70824 20508
rect 70870 20462 70928 20508
rect 70974 20462 71000 20508
rect 37542 20404 37786 20430
rect 37542 20398 37674 20404
tri 37542 20273 37667 20398 ne
rect 37667 20358 37674 20398
rect 37720 20358 37786 20404
rect 37667 20273 37786 20358
tri 37786 20273 37943 20430 sw
rect 70802 20404 71000 20462
rect 70802 20358 70824 20404
rect 70870 20358 70928 20404
rect 70974 20358 71000 20404
rect 70802 20300 71000 20358
tri 37667 20134 37806 20273 ne
rect 37806 20272 37943 20273
rect 37852 20226 37943 20272
rect 37806 20154 37943 20226
tri 37943 20154 38062 20273 sw
rect 70802 20254 70824 20300
rect 70870 20254 70928 20300
rect 70974 20254 71000 20300
rect 70802 20196 71000 20254
rect 37806 20140 38062 20154
rect 37806 20134 37938 20140
tri 37806 20002 37938 20134 ne
rect 37984 20094 38062 20140
rect 37938 20019 38062 20094
tri 38062 20019 38197 20154 sw
rect 70802 20150 70824 20196
rect 70870 20150 70928 20196
rect 70974 20150 71000 20196
rect 70802 20092 71000 20150
rect 70802 20046 70824 20092
rect 70870 20046 70928 20092
rect 70974 20046 71000 20092
rect 37938 20008 38197 20019
rect 37938 20002 38070 20008
tri 37938 19870 38070 20002 ne
rect 38116 19962 38197 20008
rect 38070 19884 38197 19962
tri 38197 19884 38332 20019 sw
rect 70802 19988 71000 20046
rect 70802 19942 70824 19988
rect 70870 19942 70928 19988
rect 70974 19942 71000 19988
rect 70802 19884 71000 19942
rect 38070 19876 38332 19884
rect 38070 19870 38202 19876
tri 38070 19738 38202 19870 ne
rect 38248 19830 38332 19876
rect 38202 19766 38332 19830
tri 38332 19766 38450 19884 sw
rect 70802 19838 70824 19884
rect 70870 19838 70928 19884
rect 70974 19838 71000 19884
rect 70802 19780 71000 19838
rect 38202 19744 38450 19766
rect 38202 19738 38334 19744
tri 38202 19608 38332 19738 ne
rect 38332 19698 38334 19738
rect 38380 19698 38450 19744
rect 38332 19653 38450 19698
tri 38450 19653 38563 19766 sw
rect 70802 19734 70824 19780
rect 70870 19734 70928 19780
rect 70974 19734 71000 19780
rect 70802 19676 71000 19734
rect 38332 19612 38563 19653
rect 38332 19608 38466 19612
tri 38332 19474 38466 19608 ne
rect 38512 19566 38563 19612
rect 38466 19490 38563 19566
tri 38563 19490 38726 19653 sw
rect 70802 19630 70824 19676
rect 70870 19630 70928 19676
rect 70974 19630 71000 19676
rect 70802 19572 71000 19630
rect 70802 19526 70824 19572
rect 70870 19526 70928 19572
rect 70974 19526 71000 19572
rect 38466 19480 38726 19490
rect 38466 19474 38598 19480
tri 38466 19355 38585 19474 ne
rect 38585 19434 38598 19474
rect 38644 19434 38726 19480
rect 38585 19377 38726 19434
tri 38726 19377 38839 19490 sw
rect 70802 19468 71000 19526
rect 70802 19422 70824 19468
rect 70870 19422 70928 19468
rect 70974 19422 71000 19468
rect 38585 19355 38839 19377
tri 38585 19210 38730 19355 ne
rect 38730 19348 38839 19355
rect 38776 19302 38839 19348
rect 38730 19242 38839 19302
tri 38839 19242 38974 19377 sw
rect 70802 19364 71000 19422
rect 70802 19318 70824 19364
rect 70870 19318 70928 19364
rect 70974 19318 71000 19364
rect 70802 19260 71000 19318
rect 38730 19216 38974 19242
rect 38730 19210 38862 19216
tri 38730 19079 38861 19210 ne
rect 38861 19170 38862 19210
rect 38908 19170 38974 19216
rect 38861 19124 38974 19170
tri 38974 19124 39092 19242 sw
rect 70802 19214 70824 19260
rect 70870 19214 70928 19260
rect 70974 19214 71000 19260
rect 70802 19156 71000 19214
rect 38861 19084 39092 19124
rect 38861 19079 38994 19084
tri 38861 18946 38994 19079 ne
rect 39040 19038 39092 19084
rect 38994 18966 39092 19038
tri 39092 18966 39250 19124 sw
rect 70802 19110 70824 19156
rect 70870 19110 70928 19156
rect 70974 19110 71000 19156
rect 70802 19052 71000 19110
rect 70802 19006 70824 19052
rect 70870 19006 70928 19052
rect 70974 19006 71000 19052
rect 38994 18952 39250 18966
rect 38994 18946 39126 18952
tri 38994 18840 39100 18946 ne
rect 39100 18906 39126 18946
rect 39172 18906 39250 18952
rect 39100 18840 39250 18906
tri 39100 18690 39250 18840 ne
tri 39250 18831 39385 18966 sw
rect 70802 18948 71000 19006
rect 70802 18902 70824 18948
rect 70870 18902 70928 18948
rect 70974 18902 71000 18948
rect 70802 18844 71000 18902
rect 39250 18820 39385 18831
rect 39250 18774 39258 18820
rect 39304 18774 39385 18820
rect 39250 18707 39385 18774
tri 39385 18707 39509 18831 sw
rect 70802 18798 70824 18844
rect 70870 18798 70928 18844
rect 70974 18798 71000 18844
rect 70802 18740 71000 18798
rect 39250 18690 39509 18707
tri 39250 18555 39385 18690 ne
rect 39385 18688 39509 18690
rect 39385 18642 39390 18688
rect 39436 18642 39509 18688
rect 39385 18600 39509 18642
tri 39509 18600 39616 18707 sw
rect 70802 18694 70824 18740
rect 70870 18694 70928 18740
rect 70974 18694 71000 18740
rect 70802 18636 71000 18694
rect 39385 18556 39616 18600
rect 39385 18555 39522 18556
tri 39385 18418 39522 18555 ne
rect 39568 18510 39616 18556
rect 39522 18431 39616 18510
tri 39616 18431 39785 18600 sw
rect 70802 18590 70824 18636
rect 70870 18590 70928 18636
rect 70974 18590 71000 18636
rect 70802 18532 71000 18590
rect 70802 18486 70824 18532
rect 70870 18486 70928 18532
rect 70974 18486 71000 18532
rect 39522 18424 39785 18431
rect 39522 18418 39654 18424
tri 39522 18296 39644 18418 ne
rect 39644 18378 39654 18418
rect 39700 18378 39785 18424
rect 39644 18296 39785 18378
tri 39785 18296 39920 18431 sw
rect 70802 18428 71000 18486
rect 70802 18382 70824 18428
rect 70870 18382 70928 18428
rect 70974 18382 71000 18428
rect 70802 18324 71000 18382
tri 39644 18154 39786 18296 ne
rect 39786 18292 39920 18296
rect 39832 18246 39920 18292
rect 39786 18189 39920 18246
tri 39920 18189 40027 18296 sw
rect 70802 18278 70824 18324
rect 70870 18278 70928 18324
rect 70974 18278 71000 18324
rect 70802 18220 71000 18278
rect 39786 18160 40027 18189
rect 39786 18154 39918 18160
tri 39786 18065 39875 18154 ne
rect 39875 18114 39918 18154
rect 39964 18114 40027 18160
rect 39875 18065 40027 18114
tri 40027 18065 40151 18189 sw
rect 70802 18174 70824 18220
rect 70870 18174 70928 18220
rect 70974 18174 71000 18220
rect 70802 18116 71000 18174
rect 70802 18070 70824 18116
rect 70870 18070 70928 18116
rect 70974 18070 71000 18116
tri 39875 17890 40050 18065 ne
rect 40050 18028 40151 18065
rect 40096 17982 40151 18028
rect 40050 17913 40151 17982
tri 40151 17913 40303 18065 sw
rect 70802 18012 71000 18070
rect 70802 17966 70824 18012
rect 70870 17966 70928 18012
rect 70974 17966 71000 18012
rect 40050 17896 40303 17913
rect 40050 17890 40182 17896
tri 40050 17789 40151 17890 ne
rect 40151 17850 40182 17890
rect 40228 17850 40303 17896
rect 40151 17789 40303 17850
tri 40151 17637 40303 17789 ne
tri 40303 17778 40438 17913 sw
rect 70802 17908 71000 17966
rect 70802 17862 70824 17908
rect 70870 17862 70928 17908
rect 70974 17862 71000 17908
rect 70802 17804 71000 17862
rect 40303 17764 40438 17778
rect 40303 17718 40314 17764
rect 40360 17718 40438 17764
rect 40303 17648 40438 17718
tri 40438 17648 40568 17778 sw
rect 70802 17758 70824 17804
rect 70870 17758 70928 17804
rect 70974 17758 71000 17804
rect 70802 17700 71000 17758
rect 70802 17654 70824 17700
rect 70870 17654 70928 17700
rect 70974 17654 71000 17700
rect 40303 17637 40568 17648
tri 40303 17502 40438 17637 ne
rect 40438 17632 40568 17637
rect 40438 17586 40446 17632
rect 40492 17586 40568 17632
rect 40438 17502 40568 17586
tri 40568 17502 40714 17648 sw
rect 70802 17596 71000 17654
rect 70802 17550 70824 17596
rect 70870 17550 70928 17596
rect 70974 17550 71000 17596
tri 40438 17362 40578 17502 ne
rect 40578 17500 40714 17502
rect 40624 17454 40714 17500
rect 40578 17412 40714 17454
tri 40714 17412 40804 17502 sw
rect 70802 17492 71000 17550
rect 70802 17446 70824 17492
rect 70870 17446 70928 17492
rect 70974 17446 71000 17492
rect 40578 17368 40804 17412
rect 40578 17362 40710 17368
tri 40578 17237 40703 17362 ne
rect 40703 17322 40710 17362
rect 40756 17322 40804 17368
rect 40703 17237 40804 17322
tri 40804 17237 40979 17412 sw
rect 70802 17388 71000 17446
rect 70802 17342 70824 17388
rect 70870 17342 70928 17388
rect 70974 17342 71000 17388
rect 70802 17284 71000 17342
rect 70802 17238 70824 17284
rect 70870 17238 70928 17284
rect 70974 17238 71000 17284
tri 40703 17098 40842 17237 ne
rect 40842 17236 40979 17237
rect 40888 17190 40979 17236
rect 40842 17136 40979 17190
tri 40979 17136 41080 17237 sw
rect 70802 17180 71000 17238
rect 40842 17104 41080 17136
rect 40842 17098 40974 17104
tri 40842 16966 40974 17098 ne
rect 41020 17058 41080 17104
rect 40974 17006 41080 17058
tri 41080 17006 41210 17136 sw
rect 70802 17134 70824 17180
rect 70870 17134 70928 17180
rect 70974 17134 71000 17180
rect 70802 17076 71000 17134
rect 70802 17030 70824 17076
rect 70870 17030 70928 17076
rect 70974 17030 71000 17076
rect 40974 16972 41210 17006
rect 40974 16966 41106 16972
tri 40974 16834 41106 16966 ne
rect 41152 16926 41210 16972
rect 41106 16860 41210 16926
tri 41210 16860 41356 17006 sw
rect 70802 16972 71000 17030
rect 70802 16926 70824 16972
rect 70870 16926 70928 16972
rect 70974 16926 71000 16972
rect 70802 16868 71000 16926
rect 41106 16840 41356 16860
rect 41106 16834 41238 16840
tri 41106 16702 41238 16834 ne
rect 41284 16794 41356 16840
rect 41238 16725 41356 16794
tri 41356 16725 41491 16860 sw
rect 70802 16822 70824 16868
rect 70870 16822 70928 16868
rect 70974 16822 71000 16868
rect 70802 16764 71000 16822
rect 41238 16708 41491 16725
rect 41238 16702 41370 16708
tri 41238 16570 41370 16702 ne
rect 41416 16662 41491 16708
rect 41370 16590 41491 16662
tri 41491 16590 41626 16725 sw
rect 70802 16718 70824 16764
rect 70870 16718 70928 16764
rect 70974 16718 71000 16764
rect 70802 16660 71000 16718
rect 70802 16614 70824 16660
rect 70870 16614 70928 16660
rect 70974 16614 71000 16660
rect 41370 16576 41626 16590
rect 41370 16570 41502 16576
tri 41370 16438 41502 16570 ne
rect 41548 16530 41626 16576
rect 41502 16454 41626 16530
tri 41626 16454 41762 16590 sw
rect 70802 16556 71000 16614
rect 70802 16510 70824 16556
rect 70870 16510 70928 16556
rect 70974 16510 71000 16556
rect 41502 16444 41762 16454
rect 41502 16438 41634 16444
tri 41502 16306 41634 16438 ne
rect 41680 16398 41762 16444
rect 41634 16314 41762 16398
tri 41762 16314 41902 16454 sw
rect 70802 16452 71000 16510
rect 70802 16406 70824 16452
rect 70870 16406 70928 16452
rect 70974 16406 71000 16452
rect 70802 16348 71000 16406
rect 41634 16312 41902 16314
rect 41634 16306 41766 16312
tri 41634 16174 41766 16306 ne
rect 41812 16266 41902 16312
rect 41766 16223 41902 16266
tri 41902 16223 41993 16314 sw
rect 70802 16302 70824 16348
rect 70870 16302 70928 16348
rect 70974 16302 71000 16348
rect 70802 16244 71000 16302
rect 41766 16180 41993 16223
rect 41766 16174 41898 16180
tri 41766 16043 41897 16174 ne
rect 41897 16134 41898 16174
rect 41944 16134 41993 16180
rect 41897 16083 41993 16134
tri 41993 16083 42133 16223 sw
rect 70802 16198 70824 16244
rect 70870 16198 70928 16244
rect 70974 16198 71000 16244
rect 70802 16140 71000 16198
rect 70802 16094 70824 16140
rect 70870 16094 70928 16140
rect 70974 16094 71000 16140
rect 41897 16048 42133 16083
rect 41897 16043 42030 16048
tri 41897 15910 42030 16043 ne
rect 42076 16002 42133 16048
rect 42030 15948 42133 16002
tri 42133 15948 42268 16083 sw
rect 70802 16036 71000 16094
rect 70802 15990 70824 16036
rect 70870 15990 70928 16036
rect 70974 15990 71000 16036
rect 42030 15916 42268 15948
rect 42030 15910 42162 15916
tri 42030 15812 42128 15910 ne
rect 42128 15870 42162 15910
rect 42208 15870 42268 15916
rect 42128 15812 42268 15870
tri 42268 15812 42404 15948 sw
rect 70802 15932 71000 15990
rect 70802 15886 70824 15932
rect 70870 15886 70928 15932
rect 70974 15886 71000 15932
rect 70802 15828 71000 15886
tri 42128 15646 42294 15812 ne
rect 42294 15784 42404 15812
rect 42340 15738 42404 15784
rect 42294 15672 42404 15738
tri 42404 15672 42544 15812 sw
rect 70802 15782 70824 15828
rect 70870 15782 70928 15828
rect 70974 15782 71000 15828
rect 70802 15724 71000 15782
rect 70802 15678 70824 15724
rect 70870 15678 70928 15724
rect 70974 15678 71000 15724
rect 42294 15652 42544 15672
rect 42294 15646 42426 15652
tri 42294 15557 42383 15646 ne
rect 42383 15606 42426 15646
rect 42472 15606 42544 15652
rect 42383 15557 42544 15606
tri 42383 15396 42544 15557 ne
tri 42544 15536 42680 15672 sw
rect 70802 15620 71000 15678
rect 70802 15574 70824 15620
rect 70870 15574 70928 15620
rect 70974 15574 71000 15620
rect 42544 15520 42680 15536
rect 42544 15474 42558 15520
rect 42604 15474 42680 15520
rect 42544 15396 42680 15474
tri 42544 15261 42679 15396 ne
rect 42679 15395 42680 15396
tri 42680 15395 42821 15536 sw
rect 70802 15516 71000 15574
rect 70802 15470 70824 15516
rect 70870 15470 70928 15516
rect 70974 15470 71000 15516
rect 70802 15412 71000 15470
rect 42679 15388 42821 15395
rect 42679 15342 42690 15388
rect 42736 15342 42821 15388
rect 42679 15261 42821 15342
tri 42821 15261 42955 15395 sw
rect 70802 15366 70824 15412
rect 70870 15366 70928 15412
rect 70974 15366 71000 15412
rect 70802 15308 71000 15366
rect 70802 15262 70824 15308
rect 70870 15262 70928 15308
rect 70974 15262 71000 15308
tri 42679 15118 42822 15261 ne
rect 42822 15256 42955 15261
rect 42868 15210 42955 15256
rect 42822 15126 42955 15210
tri 42955 15126 43090 15261 sw
rect 70802 15204 71000 15262
rect 70802 15158 70824 15204
rect 70870 15158 70928 15204
rect 70974 15158 71000 15204
rect 42822 15124 43090 15126
rect 42822 15118 42954 15124
tri 42822 15029 42911 15118 ne
rect 42911 15078 42954 15118
rect 43000 15078 43090 15124
rect 42911 15029 43090 15078
tri 43090 15029 43187 15126 sw
rect 70802 15100 71000 15158
rect 70802 15054 70824 15100
rect 70870 15054 70928 15100
rect 70974 15054 71000 15100
tri 42911 14854 43086 15029 ne
rect 43086 14992 43187 15029
rect 43132 14946 43187 14992
rect 43086 14895 43187 14946
tri 43187 14895 43321 15029 sw
rect 70802 14996 71000 15054
rect 70802 14950 70824 14996
rect 70870 14950 70928 14996
rect 70974 14950 71000 14996
rect 43086 14860 43321 14895
rect 43086 14854 43218 14860
tri 43086 14753 43187 14854 ne
rect 43187 14814 43218 14854
rect 43264 14814 43321 14860
rect 43187 14753 43321 14814
tri 43321 14753 43463 14895 sw
rect 70802 14892 71000 14950
rect 70802 14846 70824 14892
rect 70870 14846 70928 14892
rect 70974 14846 71000 14892
rect 70802 14788 71000 14846
tri 43187 14590 43350 14753 ne
rect 43350 14728 43463 14753
rect 43396 14682 43463 14728
rect 43350 14619 43463 14682
tri 43463 14619 43597 14753 sw
rect 70802 14742 70824 14788
rect 70870 14742 70928 14788
rect 70974 14742 71000 14788
rect 70802 14684 71000 14742
rect 70802 14638 70824 14684
rect 70870 14638 70928 14684
rect 70974 14638 71000 14684
rect 43350 14596 43597 14619
rect 43350 14590 43482 14596
tri 43350 14462 43478 14590 ne
rect 43478 14550 43482 14590
rect 43528 14550 43597 14596
rect 43478 14477 43597 14550
tri 43597 14477 43739 14619 sw
rect 70802 14580 71000 14638
rect 70802 14534 70824 14580
rect 70870 14534 70928 14580
rect 70974 14534 71000 14580
rect 43478 14464 43739 14477
rect 43478 14462 43614 14464
tri 43478 14326 43614 14462 ne
rect 43660 14418 43739 14464
rect 43614 14336 43739 14418
tri 43739 14336 43880 14477 sw
rect 70802 14476 71000 14534
rect 70802 14430 70824 14476
rect 70870 14430 70928 14476
rect 70974 14430 71000 14476
rect 70802 14372 71000 14430
rect 43614 14332 43880 14336
rect 43614 14326 43746 14332
tri 43614 14201 43739 14326 ne
rect 43739 14286 43746 14326
rect 43792 14286 43880 14332
rect 43739 14201 43880 14286
tri 43880 14201 44015 14336 sw
rect 70802 14326 70824 14372
rect 70870 14326 70928 14372
rect 70974 14326 71000 14372
rect 70802 14268 71000 14326
rect 70802 14222 70824 14268
rect 70870 14222 70928 14268
rect 70974 14222 71000 14268
tri 43739 14062 43878 14201 ne
rect 43878 14200 44015 14201
rect 43924 14154 44015 14200
rect 43878 14073 44015 14154
tri 44015 14073 44143 14201 sw
rect 70802 14164 71000 14222
rect 70802 14118 70824 14164
rect 70870 14118 70928 14164
rect 70974 14118 71000 14164
rect 43878 14068 44143 14073
rect 43878 14062 44010 14068
tri 43878 13930 44010 14062 ne
rect 44056 14022 44143 14068
rect 44010 13970 44143 14022
tri 44143 13970 44246 14073 sw
rect 70802 14060 71000 14118
rect 70802 14014 70824 14060
rect 70870 14014 70928 14060
rect 70974 14014 71000 14060
rect 44010 13936 44246 13970
rect 44010 13930 44142 13936
tri 44010 13798 44142 13930 ne
rect 44188 13890 44246 13936
rect 44142 13842 44246 13890
tri 44246 13842 44374 13970 sw
rect 70802 13956 71000 14014
rect 70802 13910 70824 13956
rect 70870 13910 70928 13956
rect 70974 13910 71000 13956
rect 70802 13852 71000 13910
rect 44142 13804 44374 13842
rect 44142 13798 44274 13804
tri 44142 13666 44274 13798 ne
rect 44320 13758 44374 13804
rect 44274 13694 44374 13758
tri 44374 13694 44522 13842 sw
rect 70802 13806 70824 13852
rect 70870 13806 70928 13852
rect 70974 13806 71000 13852
rect 70802 13748 71000 13806
rect 70802 13702 70824 13748
rect 70870 13702 70928 13748
rect 70974 13702 71000 13748
rect 44274 13672 44522 13694
rect 44274 13666 44406 13672
tri 44274 13534 44406 13666 ne
rect 44452 13626 44522 13672
rect 44406 13559 44522 13626
tri 44522 13559 44657 13694 sw
rect 70802 13644 71000 13702
rect 70802 13598 70824 13644
rect 70870 13598 70928 13644
rect 70974 13598 71000 13644
rect 44406 13540 44657 13559
rect 44406 13534 44538 13540
tri 44406 13402 44538 13534 ne
rect 44584 13494 44657 13540
rect 44538 13431 44657 13494
tri 44657 13431 44785 13559 sw
rect 70802 13540 71000 13598
rect 70802 13494 70824 13540
rect 70870 13494 70928 13540
rect 70974 13494 71000 13540
rect 70802 13436 71000 13494
rect 44538 13408 44785 13431
rect 44538 13402 44670 13408
tri 44538 13291 44649 13402 ne
rect 44649 13362 44670 13402
rect 44716 13362 44785 13408
rect 44649 13291 44785 13362
tri 44785 13291 44925 13431 sw
rect 70802 13390 70824 13436
rect 70870 13390 70928 13436
rect 70974 13390 71000 13436
rect 70802 13291 71000 13390
tri 44649 13097 44843 13291 ne
rect 44843 13269 71000 13291
rect 44843 13256 45088 13269
rect 44843 13210 44850 13256
rect 44896 13223 45088 13256
rect 45134 13223 45192 13269
rect 45238 13223 45296 13269
rect 45342 13223 45400 13269
rect 45446 13223 45504 13269
rect 45550 13223 45608 13269
rect 45654 13223 45712 13269
rect 45758 13223 45816 13269
rect 45862 13223 45920 13269
rect 45966 13223 46024 13269
rect 46070 13223 46128 13269
rect 46174 13223 46232 13269
rect 46278 13223 46336 13269
rect 46382 13223 46440 13269
rect 46486 13223 46544 13269
rect 46590 13223 46648 13269
rect 46694 13223 46752 13269
rect 46798 13223 46856 13269
rect 46902 13223 46960 13269
rect 47006 13223 47064 13269
rect 47110 13223 47168 13269
rect 47214 13223 47272 13269
rect 47318 13223 47376 13269
rect 47422 13223 47480 13269
rect 47526 13223 47584 13269
rect 47630 13223 47688 13269
rect 47734 13223 47792 13269
rect 47838 13223 47896 13269
rect 47942 13223 48000 13269
rect 48046 13223 48104 13269
rect 48150 13223 48208 13269
rect 48254 13223 48312 13269
rect 48358 13223 48416 13269
rect 48462 13223 48520 13269
rect 48566 13223 48624 13269
rect 48670 13223 48728 13269
rect 48774 13223 48832 13269
rect 48878 13223 48936 13269
rect 48982 13223 49040 13269
rect 49086 13223 49144 13269
rect 49190 13223 49248 13269
rect 49294 13223 49352 13269
rect 49398 13223 49456 13269
rect 49502 13223 49560 13269
rect 49606 13223 49664 13269
rect 49710 13223 49768 13269
rect 49814 13223 49872 13269
rect 49918 13223 49976 13269
rect 50022 13223 50080 13269
rect 50126 13223 50184 13269
rect 50230 13223 50288 13269
rect 50334 13223 50392 13269
rect 50438 13223 50496 13269
rect 50542 13223 50600 13269
rect 50646 13223 50704 13269
rect 50750 13223 50808 13269
rect 50854 13223 50912 13269
rect 50958 13223 51016 13269
rect 51062 13223 51120 13269
rect 51166 13223 51224 13269
rect 51270 13223 51328 13269
rect 51374 13223 51432 13269
rect 51478 13223 51536 13269
rect 51582 13223 51640 13269
rect 51686 13223 51744 13269
rect 51790 13223 51848 13269
rect 51894 13223 51952 13269
rect 51998 13223 52056 13269
rect 52102 13223 52160 13269
rect 52206 13223 52264 13269
rect 52310 13223 52368 13269
rect 52414 13223 52472 13269
rect 52518 13223 52576 13269
rect 52622 13223 52680 13269
rect 52726 13223 52784 13269
rect 52830 13223 52888 13269
rect 52934 13223 52992 13269
rect 53038 13223 53096 13269
rect 53142 13223 53200 13269
rect 53246 13223 53304 13269
rect 53350 13223 53408 13269
rect 53454 13223 53512 13269
rect 53558 13223 53616 13269
rect 53662 13223 53720 13269
rect 53766 13223 53824 13269
rect 53870 13223 53928 13269
rect 53974 13223 54032 13269
rect 54078 13223 54136 13269
rect 54182 13223 54240 13269
rect 54286 13223 54344 13269
rect 54390 13223 54448 13269
rect 54494 13223 54552 13269
rect 54598 13223 54656 13269
rect 54702 13223 54760 13269
rect 54806 13223 54864 13269
rect 54910 13223 54968 13269
rect 55014 13223 55072 13269
rect 55118 13223 55176 13269
rect 55222 13223 55280 13269
rect 55326 13223 55384 13269
rect 55430 13223 55488 13269
rect 55534 13223 55592 13269
rect 55638 13223 55696 13269
rect 55742 13223 55800 13269
rect 55846 13223 55904 13269
rect 55950 13223 56008 13269
rect 56054 13223 56112 13269
rect 56158 13223 56216 13269
rect 56262 13223 56320 13269
rect 56366 13223 56424 13269
rect 56470 13223 56528 13269
rect 56574 13223 56632 13269
rect 56678 13223 56736 13269
rect 56782 13223 56840 13269
rect 56886 13223 56944 13269
rect 56990 13223 57048 13269
rect 57094 13223 57152 13269
rect 57198 13223 57256 13269
rect 57302 13223 57360 13269
rect 57406 13223 57464 13269
rect 57510 13223 57568 13269
rect 57614 13223 57672 13269
rect 57718 13223 57776 13269
rect 57822 13223 57880 13269
rect 57926 13223 57984 13269
rect 58030 13223 58088 13269
rect 58134 13223 58192 13269
rect 58238 13223 58296 13269
rect 58342 13223 58400 13269
rect 58446 13223 58504 13269
rect 58550 13223 58608 13269
rect 58654 13223 58712 13269
rect 58758 13223 58816 13269
rect 58862 13223 58920 13269
rect 58966 13223 59024 13269
rect 59070 13223 59128 13269
rect 59174 13223 59232 13269
rect 59278 13223 59336 13269
rect 59382 13223 59440 13269
rect 59486 13223 59544 13269
rect 59590 13223 59648 13269
rect 59694 13223 59752 13269
rect 59798 13223 59856 13269
rect 59902 13223 59960 13269
rect 60006 13223 60064 13269
rect 60110 13223 60168 13269
rect 60214 13223 60272 13269
rect 60318 13223 60376 13269
rect 60422 13223 60480 13269
rect 60526 13223 60584 13269
rect 60630 13223 60688 13269
rect 60734 13223 60792 13269
rect 60838 13223 60896 13269
rect 60942 13223 61000 13269
rect 61046 13223 61104 13269
rect 61150 13223 61208 13269
rect 61254 13223 61312 13269
rect 61358 13223 61416 13269
rect 61462 13223 61520 13269
rect 61566 13223 61624 13269
rect 61670 13223 61728 13269
rect 61774 13223 61832 13269
rect 61878 13223 61936 13269
rect 61982 13223 62040 13269
rect 62086 13223 62144 13269
rect 62190 13223 62248 13269
rect 62294 13223 62352 13269
rect 62398 13223 62456 13269
rect 62502 13223 62560 13269
rect 62606 13223 62664 13269
rect 62710 13223 62768 13269
rect 62814 13223 62872 13269
rect 62918 13223 62976 13269
rect 63022 13223 63080 13269
rect 63126 13223 63184 13269
rect 63230 13223 63288 13269
rect 63334 13223 63392 13269
rect 63438 13223 63496 13269
rect 63542 13223 63600 13269
rect 63646 13223 63704 13269
rect 63750 13223 63808 13269
rect 63854 13223 63912 13269
rect 63958 13223 64016 13269
rect 64062 13223 64120 13269
rect 64166 13223 64224 13269
rect 64270 13223 64328 13269
rect 64374 13223 64432 13269
rect 64478 13223 64536 13269
rect 64582 13223 64640 13269
rect 64686 13223 64744 13269
rect 64790 13223 64848 13269
rect 64894 13223 64952 13269
rect 64998 13223 65056 13269
rect 65102 13223 65160 13269
rect 65206 13223 65264 13269
rect 65310 13223 65368 13269
rect 65414 13223 65472 13269
rect 65518 13223 65576 13269
rect 65622 13223 65680 13269
rect 65726 13223 65784 13269
rect 65830 13223 65888 13269
rect 65934 13223 65992 13269
rect 66038 13223 66096 13269
rect 66142 13223 66200 13269
rect 66246 13223 66304 13269
rect 66350 13223 66408 13269
rect 66454 13223 66512 13269
rect 66558 13223 66616 13269
rect 66662 13223 66720 13269
rect 66766 13223 66824 13269
rect 66870 13223 66928 13269
rect 66974 13223 67032 13269
rect 67078 13223 67136 13269
rect 67182 13223 67240 13269
rect 67286 13223 67344 13269
rect 67390 13223 67448 13269
rect 67494 13223 67552 13269
rect 67598 13223 67656 13269
rect 67702 13223 67760 13269
rect 67806 13223 67864 13269
rect 67910 13223 67968 13269
rect 68014 13223 68072 13269
rect 68118 13223 68176 13269
rect 68222 13223 68280 13269
rect 68326 13223 68384 13269
rect 68430 13223 68488 13269
rect 68534 13223 68592 13269
rect 68638 13223 68696 13269
rect 68742 13223 68800 13269
rect 68846 13223 68904 13269
rect 68950 13223 69008 13269
rect 69054 13223 69112 13269
rect 69158 13223 69216 13269
rect 69262 13223 69320 13269
rect 69366 13223 69424 13269
rect 69470 13223 69528 13269
rect 69574 13223 69632 13269
rect 69678 13223 69736 13269
rect 69782 13223 69840 13269
rect 69886 13223 69944 13269
rect 69990 13223 70048 13269
rect 70094 13223 70152 13269
rect 70198 13223 70256 13269
rect 70302 13223 70360 13269
rect 70406 13223 70464 13269
rect 70510 13223 70568 13269
rect 70614 13223 70672 13269
rect 70718 13223 70776 13269
rect 70822 13223 70880 13269
rect 70926 13223 71000 13269
rect 44896 13210 71000 13223
rect 44843 13165 71000 13210
rect 44843 13119 45088 13165
rect 45134 13119 45192 13165
rect 45238 13119 45296 13165
rect 45342 13119 45400 13165
rect 45446 13119 45504 13165
rect 45550 13119 45608 13165
rect 45654 13119 45712 13165
rect 45758 13119 45816 13165
rect 45862 13119 45920 13165
rect 45966 13119 46024 13165
rect 46070 13119 46128 13165
rect 46174 13119 46232 13165
rect 46278 13119 46336 13165
rect 46382 13119 46440 13165
rect 46486 13119 46544 13165
rect 46590 13119 46648 13165
rect 46694 13119 46752 13165
rect 46798 13119 46856 13165
rect 46902 13119 46960 13165
rect 47006 13119 47064 13165
rect 47110 13119 47168 13165
rect 47214 13119 47272 13165
rect 47318 13119 47376 13165
rect 47422 13119 47480 13165
rect 47526 13119 47584 13165
rect 47630 13119 47688 13165
rect 47734 13119 47792 13165
rect 47838 13119 47896 13165
rect 47942 13119 48000 13165
rect 48046 13119 48104 13165
rect 48150 13119 48208 13165
rect 48254 13119 48312 13165
rect 48358 13119 48416 13165
rect 48462 13119 48520 13165
rect 48566 13119 48624 13165
rect 48670 13119 48728 13165
rect 48774 13119 48832 13165
rect 48878 13119 48936 13165
rect 48982 13119 49040 13165
rect 49086 13119 49144 13165
rect 49190 13119 49248 13165
rect 49294 13119 49352 13165
rect 49398 13119 49456 13165
rect 49502 13119 49560 13165
rect 49606 13119 49664 13165
rect 49710 13119 49768 13165
rect 49814 13119 49872 13165
rect 49918 13119 49976 13165
rect 50022 13119 50080 13165
rect 50126 13119 50184 13165
rect 50230 13119 50288 13165
rect 50334 13119 50392 13165
rect 50438 13119 50496 13165
rect 50542 13119 50600 13165
rect 50646 13119 50704 13165
rect 50750 13119 50808 13165
rect 50854 13119 50912 13165
rect 50958 13119 51016 13165
rect 51062 13119 51120 13165
rect 51166 13119 51224 13165
rect 51270 13119 51328 13165
rect 51374 13119 51432 13165
rect 51478 13119 51536 13165
rect 51582 13119 51640 13165
rect 51686 13119 51744 13165
rect 51790 13119 51848 13165
rect 51894 13119 51952 13165
rect 51998 13119 52056 13165
rect 52102 13119 52160 13165
rect 52206 13119 52264 13165
rect 52310 13119 52368 13165
rect 52414 13119 52472 13165
rect 52518 13119 52576 13165
rect 52622 13119 52680 13165
rect 52726 13119 52784 13165
rect 52830 13119 52888 13165
rect 52934 13119 52992 13165
rect 53038 13119 53096 13165
rect 53142 13119 53200 13165
rect 53246 13119 53304 13165
rect 53350 13119 53408 13165
rect 53454 13119 53512 13165
rect 53558 13119 53616 13165
rect 53662 13119 53720 13165
rect 53766 13119 53824 13165
rect 53870 13119 53928 13165
rect 53974 13119 54032 13165
rect 54078 13119 54136 13165
rect 54182 13119 54240 13165
rect 54286 13119 54344 13165
rect 54390 13119 54448 13165
rect 54494 13119 54552 13165
rect 54598 13119 54656 13165
rect 54702 13119 54760 13165
rect 54806 13119 54864 13165
rect 54910 13119 54968 13165
rect 55014 13119 55072 13165
rect 55118 13119 55176 13165
rect 55222 13119 55280 13165
rect 55326 13119 55384 13165
rect 55430 13119 55488 13165
rect 55534 13119 55592 13165
rect 55638 13119 55696 13165
rect 55742 13119 55800 13165
rect 55846 13119 55904 13165
rect 55950 13119 56008 13165
rect 56054 13119 56112 13165
rect 56158 13119 56216 13165
rect 56262 13119 56320 13165
rect 56366 13119 56424 13165
rect 56470 13119 56528 13165
rect 56574 13119 56632 13165
rect 56678 13119 56736 13165
rect 56782 13119 56840 13165
rect 56886 13119 56944 13165
rect 56990 13119 57048 13165
rect 57094 13119 57152 13165
rect 57198 13119 57256 13165
rect 57302 13119 57360 13165
rect 57406 13119 57464 13165
rect 57510 13119 57568 13165
rect 57614 13119 57672 13165
rect 57718 13119 57776 13165
rect 57822 13119 57880 13165
rect 57926 13119 57984 13165
rect 58030 13119 58088 13165
rect 58134 13119 58192 13165
rect 58238 13119 58296 13165
rect 58342 13119 58400 13165
rect 58446 13119 58504 13165
rect 58550 13119 58608 13165
rect 58654 13119 58712 13165
rect 58758 13119 58816 13165
rect 58862 13119 58920 13165
rect 58966 13119 59024 13165
rect 59070 13119 59128 13165
rect 59174 13119 59232 13165
rect 59278 13119 59336 13165
rect 59382 13119 59440 13165
rect 59486 13119 59544 13165
rect 59590 13119 59648 13165
rect 59694 13119 59752 13165
rect 59798 13119 59856 13165
rect 59902 13119 59960 13165
rect 60006 13119 60064 13165
rect 60110 13119 60168 13165
rect 60214 13119 60272 13165
rect 60318 13119 60376 13165
rect 60422 13119 60480 13165
rect 60526 13119 60584 13165
rect 60630 13119 60688 13165
rect 60734 13119 60792 13165
rect 60838 13119 60896 13165
rect 60942 13119 61000 13165
rect 61046 13119 61104 13165
rect 61150 13119 61208 13165
rect 61254 13119 61312 13165
rect 61358 13119 61416 13165
rect 61462 13119 61520 13165
rect 61566 13119 61624 13165
rect 61670 13119 61728 13165
rect 61774 13119 61832 13165
rect 61878 13119 61936 13165
rect 61982 13119 62040 13165
rect 62086 13119 62144 13165
rect 62190 13119 62248 13165
rect 62294 13119 62352 13165
rect 62398 13119 62456 13165
rect 62502 13119 62560 13165
rect 62606 13119 62664 13165
rect 62710 13119 62768 13165
rect 62814 13119 62872 13165
rect 62918 13119 62976 13165
rect 63022 13119 63080 13165
rect 63126 13119 63184 13165
rect 63230 13119 63288 13165
rect 63334 13119 63392 13165
rect 63438 13119 63496 13165
rect 63542 13119 63600 13165
rect 63646 13119 63704 13165
rect 63750 13119 63808 13165
rect 63854 13119 63912 13165
rect 63958 13119 64016 13165
rect 64062 13119 64120 13165
rect 64166 13119 64224 13165
rect 64270 13119 64328 13165
rect 64374 13119 64432 13165
rect 64478 13119 64536 13165
rect 64582 13119 64640 13165
rect 64686 13119 64744 13165
rect 64790 13119 64848 13165
rect 64894 13119 64952 13165
rect 64998 13119 65056 13165
rect 65102 13119 65160 13165
rect 65206 13119 65264 13165
rect 65310 13119 65368 13165
rect 65414 13119 65472 13165
rect 65518 13119 65576 13165
rect 65622 13119 65680 13165
rect 65726 13119 65784 13165
rect 65830 13119 65888 13165
rect 65934 13119 65992 13165
rect 66038 13119 66096 13165
rect 66142 13119 66200 13165
rect 66246 13119 66304 13165
rect 66350 13119 66408 13165
rect 66454 13119 66512 13165
rect 66558 13119 66616 13165
rect 66662 13119 66720 13165
rect 66766 13119 66824 13165
rect 66870 13119 66928 13165
rect 66974 13119 67032 13165
rect 67078 13119 67136 13165
rect 67182 13119 67240 13165
rect 67286 13119 67344 13165
rect 67390 13119 67448 13165
rect 67494 13119 67552 13165
rect 67598 13119 67656 13165
rect 67702 13119 67760 13165
rect 67806 13119 67864 13165
rect 67910 13119 67968 13165
rect 68014 13119 68072 13165
rect 68118 13119 68176 13165
rect 68222 13119 68280 13165
rect 68326 13119 68384 13165
rect 68430 13119 68488 13165
rect 68534 13119 68592 13165
rect 68638 13119 68696 13165
rect 68742 13119 68800 13165
rect 68846 13119 68904 13165
rect 68950 13119 69008 13165
rect 69054 13119 69112 13165
rect 69158 13119 69216 13165
rect 69262 13119 69320 13165
rect 69366 13119 69424 13165
rect 69470 13119 69528 13165
rect 69574 13119 69632 13165
rect 69678 13119 69736 13165
rect 69782 13119 69840 13165
rect 69886 13119 69944 13165
rect 69990 13119 70048 13165
rect 70094 13119 70152 13165
rect 70198 13119 70256 13165
rect 70302 13119 70360 13165
rect 70406 13119 70464 13165
rect 70510 13119 70568 13165
rect 70614 13119 70672 13165
rect 70718 13119 70776 13165
rect 70822 13119 70880 13165
rect 70926 13119 71000 13165
rect 44843 13097 71000 13119
<< psubdiffcont >>
rect 13119 70929 13165 70975
rect 13223 70929 13269 70975
rect 13377 70929 13423 70975
rect 13481 70929 13527 70975
rect 13585 70929 13631 70975
rect 13689 70929 13735 70975
rect 13793 70929 13839 70975
rect 13897 70929 13943 70975
rect 14001 70929 14047 70975
rect 14105 70929 14151 70975
rect 14209 70929 14255 70975
rect 14313 70929 14359 70975
rect 14417 70929 14463 70975
rect 14521 70929 14567 70975
rect 14625 70929 14671 70975
rect 14729 70929 14775 70975
rect 14833 70929 14879 70975
rect 14937 70929 14983 70975
rect 15041 70929 15087 70975
rect 15145 70929 15191 70975
rect 15249 70929 15295 70975
rect 15353 70929 15399 70975
rect 15457 70929 15503 70975
rect 15561 70929 15607 70975
rect 15665 70929 15711 70975
rect 15769 70929 15815 70975
rect 15873 70929 15919 70975
rect 15977 70929 16023 70975
rect 16081 70929 16127 70975
rect 16185 70929 16231 70975
rect 16289 70929 16335 70975
rect 16393 70929 16439 70975
rect 16497 70929 16543 70975
rect 16601 70929 16647 70975
rect 16705 70929 16751 70975
rect 16809 70929 16855 70975
rect 16913 70929 16959 70975
rect 17017 70929 17063 70975
rect 17121 70929 17167 70975
rect 17225 70929 17271 70975
rect 17329 70929 17375 70975
rect 17433 70929 17479 70975
rect 17537 70929 17583 70975
rect 17641 70929 17687 70975
rect 17745 70929 17791 70975
rect 17849 70929 17895 70975
rect 17953 70929 17999 70975
rect 18057 70929 18103 70975
rect 18161 70929 18207 70975
rect 18265 70929 18311 70975
rect 18369 70929 18415 70975
rect 18473 70929 18519 70975
rect 18577 70929 18623 70975
rect 18681 70929 18727 70975
rect 18785 70929 18831 70975
rect 18889 70929 18935 70975
rect 18993 70929 19039 70975
rect 19097 70929 19143 70975
rect 19201 70929 19247 70975
rect 19305 70929 19351 70975
rect 19409 70929 19455 70975
rect 19513 70929 19559 70975
rect 19617 70929 19663 70975
rect 19721 70929 19767 70975
rect 19825 70929 19871 70975
rect 19929 70929 19975 70975
rect 20033 70929 20079 70975
rect 20137 70929 20183 70975
rect 20241 70929 20287 70975
rect 20345 70929 20391 70975
rect 20449 70929 20495 70975
rect 20553 70929 20599 70975
rect 20657 70929 20703 70975
rect 20761 70929 20807 70975
rect 20865 70929 20911 70975
rect 20969 70929 21015 70975
rect 21073 70929 21119 70975
rect 21177 70929 21223 70975
rect 21281 70929 21327 70975
rect 21385 70929 21431 70975
rect 21489 70929 21535 70975
rect 21593 70929 21639 70975
rect 21697 70929 21743 70975
rect 21801 70929 21847 70975
rect 21905 70929 21951 70975
rect 22009 70929 22055 70975
rect 22113 70929 22159 70975
rect 22217 70929 22263 70975
rect 22321 70929 22367 70975
rect 22425 70929 22471 70975
rect 22529 70929 22575 70975
rect 22633 70929 22679 70975
rect 22737 70929 22783 70975
rect 22841 70929 22887 70975
rect 22945 70929 22991 70975
rect 23049 70929 23095 70975
rect 23153 70929 23199 70975
rect 23257 70929 23303 70975
rect 23361 70929 23407 70975
rect 23465 70929 23511 70975
rect 23569 70929 23615 70975
rect 23673 70929 23719 70975
rect 23777 70929 23823 70975
rect 23881 70929 23927 70975
rect 23985 70929 24031 70975
rect 24089 70929 24135 70975
rect 24193 70929 24239 70975
rect 24297 70929 24343 70975
rect 24401 70929 24447 70975
rect 24505 70929 24551 70975
rect 24609 70929 24655 70975
rect 24713 70929 24759 70975
rect 24817 70929 24863 70975
rect 24921 70929 24967 70975
rect 25025 70929 25071 70975
rect 25129 70929 25175 70975
rect 25233 70929 25279 70975
rect 25337 70929 25383 70975
rect 25441 70929 25487 70975
rect 25545 70929 25591 70975
rect 25649 70929 25695 70975
rect 25753 70929 25799 70975
rect 25857 70929 25903 70975
rect 25961 70929 26007 70975
rect 26065 70929 26111 70975
rect 26169 70929 26215 70975
rect 26273 70929 26319 70975
rect 26377 70929 26423 70975
rect 26481 70929 26527 70975
rect 26585 70929 26631 70975
rect 26689 70929 26735 70975
rect 26793 70929 26839 70975
rect 26897 70929 26943 70975
rect 27001 70929 27047 70975
rect 27105 70929 27151 70975
rect 27209 70929 27255 70975
rect 27313 70929 27359 70975
rect 27417 70929 27463 70975
rect 27521 70929 27567 70975
rect 27625 70929 27671 70975
rect 27729 70929 27775 70975
rect 27833 70929 27879 70975
rect 27937 70929 27983 70975
rect 28041 70929 28087 70975
rect 28145 70929 28191 70975
rect 28249 70929 28295 70975
rect 28353 70929 28399 70975
rect 28457 70929 28503 70975
rect 28561 70929 28607 70975
rect 28665 70929 28711 70975
rect 28769 70929 28815 70975
rect 28873 70929 28919 70975
rect 28977 70929 29023 70975
rect 29081 70929 29127 70975
rect 29185 70929 29231 70975
rect 29289 70929 29335 70975
rect 29393 70929 29439 70975
rect 29497 70929 29543 70975
rect 29601 70929 29647 70975
rect 29705 70929 29751 70975
rect 29809 70929 29855 70975
rect 29913 70929 29959 70975
rect 30017 70929 30063 70975
rect 30121 70929 30167 70975
rect 30225 70929 30271 70975
rect 30329 70929 30375 70975
rect 30433 70929 30479 70975
rect 30537 70929 30583 70975
rect 30641 70929 30687 70975
rect 30745 70929 30791 70975
rect 30849 70929 30895 70975
rect 30953 70929 30999 70975
rect 31057 70929 31103 70975
rect 31161 70929 31207 70975
rect 31265 70929 31311 70975
rect 31369 70929 31415 70975
rect 31473 70929 31519 70975
rect 31577 70929 31623 70975
rect 31681 70929 31727 70975
rect 31785 70929 31831 70975
rect 31889 70929 31935 70975
rect 31993 70929 32039 70975
rect 32097 70929 32143 70975
rect 32201 70929 32247 70975
rect 32305 70929 32351 70975
rect 32409 70929 32455 70975
rect 32513 70929 32559 70975
rect 32617 70929 32663 70975
rect 32721 70929 32767 70975
rect 32825 70929 32871 70975
rect 32929 70929 32975 70975
rect 33033 70929 33079 70975
rect 33137 70929 33183 70975
rect 33241 70929 33287 70975
rect 33345 70929 33391 70975
rect 33449 70929 33495 70975
rect 33553 70929 33599 70975
rect 33657 70929 33703 70975
rect 33761 70929 33807 70975
rect 33865 70929 33911 70975
rect 33969 70929 34015 70975
rect 34073 70929 34119 70975
rect 34177 70929 34223 70975
rect 34281 70929 34327 70975
rect 34385 70929 34431 70975
rect 34489 70929 34535 70975
rect 34593 70929 34639 70975
rect 34697 70929 34743 70975
rect 34801 70929 34847 70975
rect 34905 70929 34951 70975
rect 35009 70929 35055 70975
rect 35113 70929 35159 70975
rect 35217 70929 35263 70975
rect 35321 70929 35367 70975
rect 35425 70929 35471 70975
rect 35529 70929 35575 70975
rect 35633 70929 35679 70975
rect 35737 70929 35783 70975
rect 35841 70929 35887 70975
rect 35945 70929 35991 70975
rect 36049 70929 36095 70975
rect 36153 70929 36199 70975
rect 36257 70929 36303 70975
rect 36361 70929 36407 70975
rect 36465 70929 36511 70975
rect 36569 70929 36615 70975
rect 36673 70929 36719 70975
rect 36777 70929 36823 70975
rect 36881 70929 36927 70975
rect 36985 70929 37031 70975
rect 37089 70929 37135 70975
rect 37193 70929 37239 70975
rect 37297 70929 37343 70975
rect 37401 70929 37447 70975
rect 37505 70929 37551 70975
rect 37609 70929 37655 70975
rect 37713 70929 37759 70975
rect 37817 70929 37863 70975
rect 37921 70929 37967 70975
rect 38025 70929 38071 70975
rect 38129 70929 38175 70975
rect 38233 70929 38279 70975
rect 38337 70929 38383 70975
rect 38441 70929 38487 70975
rect 38545 70929 38591 70975
rect 38649 70929 38695 70975
rect 38753 70929 38799 70975
rect 38857 70929 38903 70975
rect 38961 70929 39007 70975
rect 39065 70929 39111 70975
rect 39169 70929 39215 70975
rect 39273 70929 39319 70975
rect 39377 70929 39423 70975
rect 39481 70929 39527 70975
rect 39585 70929 39631 70975
rect 39689 70929 39735 70975
rect 39793 70929 39839 70975
rect 39897 70929 39943 70975
rect 40001 70929 40047 70975
rect 40105 70929 40151 70975
rect 40209 70929 40255 70975
rect 40313 70929 40359 70975
rect 40417 70929 40463 70975
rect 40521 70929 40567 70975
rect 40625 70929 40671 70975
rect 40729 70929 40775 70975
rect 40833 70929 40879 70975
rect 40937 70929 40983 70975
rect 41041 70929 41087 70975
rect 41145 70929 41191 70975
rect 41249 70929 41295 70975
rect 41353 70929 41399 70975
rect 41457 70929 41503 70975
rect 41561 70929 41607 70975
rect 41665 70929 41711 70975
rect 41769 70929 41815 70975
rect 41873 70929 41919 70975
rect 41977 70929 42023 70975
rect 42081 70929 42127 70975
rect 42185 70929 42231 70975
rect 42289 70929 42335 70975
rect 42393 70929 42439 70975
rect 42497 70929 42543 70975
rect 42601 70929 42647 70975
rect 42705 70929 42751 70975
rect 42809 70929 42855 70975
rect 42913 70929 42959 70975
rect 43017 70929 43063 70975
rect 43121 70929 43167 70975
rect 43225 70929 43271 70975
rect 43329 70929 43375 70975
rect 43433 70929 43479 70975
rect 43537 70929 43583 70975
rect 43641 70929 43687 70975
rect 43745 70929 43791 70975
rect 43849 70929 43895 70975
rect 43953 70929 43999 70975
rect 44057 70929 44103 70975
rect 44161 70929 44207 70975
rect 44265 70929 44311 70975
rect 44369 70929 44415 70975
rect 44473 70929 44519 70975
rect 44577 70929 44623 70975
rect 44681 70929 44727 70975
rect 44785 70929 44831 70975
rect 44889 70929 44935 70975
rect 44993 70929 45039 70975
rect 45097 70929 45143 70975
rect 45201 70929 45247 70975
rect 45305 70929 45351 70975
rect 45409 70929 45455 70975
rect 45513 70929 45559 70975
rect 45617 70929 45663 70975
rect 45721 70929 45767 70975
rect 45825 70929 45871 70975
rect 45929 70929 45975 70975
rect 46033 70929 46079 70975
rect 46137 70929 46183 70975
rect 46241 70929 46287 70975
rect 46345 70929 46391 70975
rect 46449 70929 46495 70975
rect 46553 70929 46599 70975
rect 46657 70929 46703 70975
rect 46761 70929 46807 70975
rect 46865 70929 46911 70975
rect 46969 70929 47015 70975
rect 47073 70929 47119 70975
rect 47177 70929 47223 70975
rect 47281 70929 47327 70975
rect 47385 70929 47431 70975
rect 47489 70929 47535 70975
rect 47593 70929 47639 70975
rect 47697 70929 47743 70975
rect 47801 70929 47847 70975
rect 47905 70929 47951 70975
rect 48009 70929 48055 70975
rect 48113 70929 48159 70975
rect 48217 70929 48263 70975
rect 48321 70929 48367 70975
rect 48425 70929 48471 70975
rect 48529 70929 48575 70975
rect 48633 70929 48679 70975
rect 48737 70929 48783 70975
rect 48841 70929 48887 70975
rect 48945 70929 48991 70975
rect 49049 70929 49095 70975
rect 49153 70929 49199 70975
rect 49257 70929 49303 70975
rect 49361 70929 49407 70975
rect 49465 70929 49511 70975
rect 49569 70929 49615 70975
rect 49673 70929 49719 70975
rect 49777 70929 49823 70975
rect 49881 70929 49927 70975
rect 49985 70929 50031 70975
rect 50089 70929 50135 70975
rect 50193 70929 50239 70975
rect 50297 70929 50343 70975
rect 50401 70929 50447 70975
rect 50505 70929 50551 70975
rect 50609 70929 50655 70975
rect 50713 70929 50759 70975
rect 50817 70929 50863 70975
rect 50921 70929 50967 70975
rect 51025 70929 51071 70975
rect 51129 70929 51175 70975
rect 51233 70929 51279 70975
rect 51337 70929 51383 70975
rect 51441 70929 51487 70975
rect 51545 70929 51591 70975
rect 51649 70929 51695 70975
rect 51753 70929 51799 70975
rect 51857 70929 51903 70975
rect 51961 70929 52007 70975
rect 52065 70929 52111 70975
rect 52169 70929 52215 70975
rect 52273 70929 52319 70975
rect 52377 70929 52423 70975
rect 52481 70929 52527 70975
rect 52585 70929 52631 70975
rect 52689 70929 52735 70975
rect 52793 70929 52839 70975
rect 52897 70929 52943 70975
rect 53001 70929 53047 70975
rect 53105 70929 53151 70975
rect 53209 70929 53255 70975
rect 53313 70929 53359 70975
rect 53417 70929 53463 70975
rect 53521 70929 53567 70975
rect 53625 70929 53671 70975
rect 53729 70929 53775 70975
rect 53833 70929 53879 70975
rect 53937 70929 53983 70975
rect 54041 70929 54087 70975
rect 54145 70929 54191 70975
rect 54249 70929 54295 70975
rect 54353 70929 54399 70975
rect 54457 70929 54503 70975
rect 54561 70929 54607 70975
rect 54665 70929 54711 70975
rect 54769 70929 54815 70975
rect 54873 70929 54919 70975
rect 54977 70929 55023 70975
rect 55081 70929 55127 70975
rect 55185 70929 55231 70975
rect 55289 70929 55335 70975
rect 55393 70929 55439 70975
rect 55497 70929 55543 70975
rect 55601 70929 55647 70975
rect 55705 70929 55751 70975
rect 55809 70929 55855 70975
rect 55913 70929 55959 70975
rect 56017 70929 56063 70975
rect 56121 70929 56167 70975
rect 56225 70929 56271 70975
rect 56329 70929 56375 70975
rect 56433 70929 56479 70975
rect 56537 70929 56583 70975
rect 56641 70929 56687 70975
rect 56745 70929 56791 70975
rect 56849 70929 56895 70975
rect 56953 70929 56999 70975
rect 57057 70929 57103 70975
rect 57161 70929 57207 70975
rect 57265 70929 57311 70975
rect 57369 70929 57415 70975
rect 57473 70929 57519 70975
rect 57577 70929 57623 70975
rect 57681 70929 57727 70975
rect 57785 70929 57831 70975
rect 57889 70929 57935 70975
rect 57993 70929 58039 70975
rect 58097 70929 58143 70975
rect 58201 70929 58247 70975
rect 58305 70929 58351 70975
rect 58409 70929 58455 70975
rect 58513 70929 58559 70975
rect 58617 70929 58663 70975
rect 58721 70929 58767 70975
rect 58825 70929 58871 70975
rect 58929 70929 58975 70975
rect 59033 70929 59079 70975
rect 59137 70929 59183 70975
rect 59241 70929 59287 70975
rect 59345 70929 59391 70975
rect 59449 70929 59495 70975
rect 59553 70929 59599 70975
rect 59657 70929 59703 70975
rect 59761 70929 59807 70975
rect 59865 70929 59911 70975
rect 59969 70929 60015 70975
rect 60073 70929 60119 70975
rect 60177 70929 60223 70975
rect 60281 70929 60327 70975
rect 60385 70929 60431 70975
rect 60489 70929 60535 70975
rect 60593 70929 60639 70975
rect 60697 70929 60743 70975
rect 60801 70929 60847 70975
rect 60905 70929 60951 70975
rect 61009 70929 61055 70975
rect 61113 70929 61159 70975
rect 61217 70929 61263 70975
rect 61321 70929 61367 70975
rect 61425 70929 61471 70975
rect 61529 70929 61575 70975
rect 61633 70929 61679 70975
rect 61737 70929 61783 70975
rect 61841 70929 61887 70975
rect 61945 70929 61991 70975
rect 62049 70929 62095 70975
rect 62153 70929 62199 70975
rect 62257 70929 62303 70975
rect 62361 70929 62407 70975
rect 62465 70929 62511 70975
rect 62569 70929 62615 70975
rect 62673 70929 62719 70975
rect 62777 70929 62823 70975
rect 62881 70929 62927 70975
rect 62985 70929 63031 70975
rect 63089 70929 63135 70975
rect 63193 70929 63239 70975
rect 63297 70929 63343 70975
rect 63401 70929 63447 70975
rect 63505 70929 63551 70975
rect 63609 70929 63655 70975
rect 63713 70929 63759 70975
rect 63817 70929 63863 70975
rect 63921 70929 63967 70975
rect 64025 70929 64071 70975
rect 64129 70929 64175 70975
rect 64233 70929 64279 70975
rect 64337 70929 64383 70975
rect 64441 70929 64487 70975
rect 64545 70929 64591 70975
rect 64649 70929 64695 70975
rect 64753 70929 64799 70975
rect 64857 70929 64903 70975
rect 64961 70929 65007 70975
rect 65065 70929 65111 70975
rect 65169 70929 65215 70975
rect 65273 70929 65319 70975
rect 65377 70929 65423 70975
rect 65481 70929 65527 70975
rect 65585 70929 65631 70975
rect 65689 70929 65735 70975
rect 65793 70929 65839 70975
rect 65897 70929 65943 70975
rect 66001 70929 66047 70975
rect 66105 70929 66151 70975
rect 66209 70929 66255 70975
rect 66313 70929 66359 70975
rect 66417 70929 66463 70975
rect 66521 70929 66567 70975
rect 66625 70929 66671 70975
rect 66729 70929 66775 70975
rect 66833 70929 66879 70975
rect 66937 70929 66983 70975
rect 67041 70929 67087 70975
rect 67145 70929 67191 70975
rect 67249 70929 67295 70975
rect 67353 70929 67399 70975
rect 67457 70929 67503 70975
rect 67561 70929 67607 70975
rect 67665 70929 67711 70975
rect 67769 70929 67815 70975
rect 67873 70929 67919 70975
rect 67977 70929 68023 70975
rect 68081 70929 68127 70975
rect 68185 70929 68231 70975
rect 68289 70929 68335 70975
rect 68393 70929 68439 70975
rect 68497 70929 68543 70975
rect 68601 70929 68647 70975
rect 68705 70929 68751 70975
rect 68809 70929 68855 70975
rect 68913 70929 68959 70975
rect 69017 70929 69063 70975
rect 69121 70929 69167 70975
rect 69225 70929 69271 70975
rect 69329 70929 69375 70975
rect 69433 70929 69479 70975
rect 69537 70929 69583 70975
rect 69641 70929 69687 70975
rect 69745 70929 69791 70975
rect 69849 70929 69895 70975
rect 13119 70825 13165 70871
rect 13223 70825 13269 70871
rect 13377 70825 13423 70871
rect 13481 70825 13527 70871
rect 13585 70825 13631 70871
rect 13689 70825 13735 70871
rect 13793 70825 13839 70871
rect 13897 70825 13943 70871
rect 14001 70825 14047 70871
rect 14105 70825 14151 70871
rect 14209 70825 14255 70871
rect 14313 70825 14359 70871
rect 14417 70825 14463 70871
rect 14521 70825 14567 70871
rect 14625 70825 14671 70871
rect 14729 70825 14775 70871
rect 14833 70825 14879 70871
rect 14937 70825 14983 70871
rect 15041 70825 15087 70871
rect 15145 70825 15191 70871
rect 15249 70825 15295 70871
rect 15353 70825 15399 70871
rect 15457 70825 15503 70871
rect 15561 70825 15607 70871
rect 15665 70825 15711 70871
rect 15769 70825 15815 70871
rect 15873 70825 15919 70871
rect 15977 70825 16023 70871
rect 16081 70825 16127 70871
rect 16185 70825 16231 70871
rect 16289 70825 16335 70871
rect 16393 70825 16439 70871
rect 16497 70825 16543 70871
rect 16601 70825 16647 70871
rect 16705 70825 16751 70871
rect 16809 70825 16855 70871
rect 16913 70825 16959 70871
rect 17017 70825 17063 70871
rect 17121 70825 17167 70871
rect 17225 70825 17271 70871
rect 17329 70825 17375 70871
rect 17433 70825 17479 70871
rect 17537 70825 17583 70871
rect 17641 70825 17687 70871
rect 17745 70825 17791 70871
rect 17849 70825 17895 70871
rect 17953 70825 17999 70871
rect 18057 70825 18103 70871
rect 18161 70825 18207 70871
rect 18265 70825 18311 70871
rect 18369 70825 18415 70871
rect 18473 70825 18519 70871
rect 18577 70825 18623 70871
rect 18681 70825 18727 70871
rect 18785 70825 18831 70871
rect 18889 70825 18935 70871
rect 18993 70825 19039 70871
rect 19097 70825 19143 70871
rect 19201 70825 19247 70871
rect 19305 70825 19351 70871
rect 19409 70825 19455 70871
rect 19513 70825 19559 70871
rect 19617 70825 19663 70871
rect 19721 70825 19767 70871
rect 19825 70825 19871 70871
rect 19929 70825 19975 70871
rect 20033 70825 20079 70871
rect 20137 70825 20183 70871
rect 20241 70825 20287 70871
rect 20345 70825 20391 70871
rect 20449 70825 20495 70871
rect 20553 70825 20599 70871
rect 20657 70825 20703 70871
rect 20761 70825 20807 70871
rect 20865 70825 20911 70871
rect 20969 70825 21015 70871
rect 21073 70825 21119 70871
rect 21177 70825 21223 70871
rect 21281 70825 21327 70871
rect 21385 70825 21431 70871
rect 21489 70825 21535 70871
rect 21593 70825 21639 70871
rect 21697 70825 21743 70871
rect 21801 70825 21847 70871
rect 21905 70825 21951 70871
rect 22009 70825 22055 70871
rect 22113 70825 22159 70871
rect 22217 70825 22263 70871
rect 22321 70825 22367 70871
rect 22425 70825 22471 70871
rect 22529 70825 22575 70871
rect 22633 70825 22679 70871
rect 22737 70825 22783 70871
rect 22841 70825 22887 70871
rect 22945 70825 22991 70871
rect 23049 70825 23095 70871
rect 23153 70825 23199 70871
rect 23257 70825 23303 70871
rect 23361 70825 23407 70871
rect 23465 70825 23511 70871
rect 23569 70825 23615 70871
rect 23673 70825 23719 70871
rect 23777 70825 23823 70871
rect 23881 70825 23927 70871
rect 23985 70825 24031 70871
rect 24089 70825 24135 70871
rect 24193 70825 24239 70871
rect 24297 70825 24343 70871
rect 24401 70825 24447 70871
rect 24505 70825 24551 70871
rect 24609 70825 24655 70871
rect 24713 70825 24759 70871
rect 24817 70825 24863 70871
rect 24921 70825 24967 70871
rect 25025 70825 25071 70871
rect 25129 70825 25175 70871
rect 25233 70825 25279 70871
rect 25337 70825 25383 70871
rect 25441 70825 25487 70871
rect 25545 70825 25591 70871
rect 25649 70825 25695 70871
rect 25753 70825 25799 70871
rect 25857 70825 25903 70871
rect 25961 70825 26007 70871
rect 26065 70825 26111 70871
rect 26169 70825 26215 70871
rect 26273 70825 26319 70871
rect 26377 70825 26423 70871
rect 26481 70825 26527 70871
rect 26585 70825 26631 70871
rect 26689 70825 26735 70871
rect 26793 70825 26839 70871
rect 26897 70825 26943 70871
rect 27001 70825 27047 70871
rect 27105 70825 27151 70871
rect 27209 70825 27255 70871
rect 27313 70825 27359 70871
rect 27417 70825 27463 70871
rect 27521 70825 27567 70871
rect 27625 70825 27671 70871
rect 27729 70825 27775 70871
rect 27833 70825 27879 70871
rect 27937 70825 27983 70871
rect 28041 70825 28087 70871
rect 28145 70825 28191 70871
rect 28249 70825 28295 70871
rect 28353 70825 28399 70871
rect 28457 70825 28503 70871
rect 28561 70825 28607 70871
rect 28665 70825 28711 70871
rect 28769 70825 28815 70871
rect 28873 70825 28919 70871
rect 28977 70825 29023 70871
rect 29081 70825 29127 70871
rect 29185 70825 29231 70871
rect 29289 70825 29335 70871
rect 29393 70825 29439 70871
rect 29497 70825 29543 70871
rect 29601 70825 29647 70871
rect 29705 70825 29751 70871
rect 29809 70825 29855 70871
rect 29913 70825 29959 70871
rect 30017 70825 30063 70871
rect 30121 70825 30167 70871
rect 30225 70825 30271 70871
rect 30329 70825 30375 70871
rect 30433 70825 30479 70871
rect 30537 70825 30583 70871
rect 30641 70825 30687 70871
rect 30745 70825 30791 70871
rect 30849 70825 30895 70871
rect 30953 70825 30999 70871
rect 31057 70825 31103 70871
rect 31161 70825 31207 70871
rect 31265 70825 31311 70871
rect 31369 70825 31415 70871
rect 31473 70825 31519 70871
rect 31577 70825 31623 70871
rect 31681 70825 31727 70871
rect 31785 70825 31831 70871
rect 31889 70825 31935 70871
rect 31993 70825 32039 70871
rect 32097 70825 32143 70871
rect 32201 70825 32247 70871
rect 32305 70825 32351 70871
rect 32409 70825 32455 70871
rect 32513 70825 32559 70871
rect 32617 70825 32663 70871
rect 32721 70825 32767 70871
rect 32825 70825 32871 70871
rect 32929 70825 32975 70871
rect 33033 70825 33079 70871
rect 33137 70825 33183 70871
rect 33241 70825 33287 70871
rect 33345 70825 33391 70871
rect 33449 70825 33495 70871
rect 33553 70825 33599 70871
rect 33657 70825 33703 70871
rect 33761 70825 33807 70871
rect 33865 70825 33911 70871
rect 33969 70825 34015 70871
rect 34073 70825 34119 70871
rect 34177 70825 34223 70871
rect 34281 70825 34327 70871
rect 34385 70825 34431 70871
rect 34489 70825 34535 70871
rect 34593 70825 34639 70871
rect 34697 70825 34743 70871
rect 34801 70825 34847 70871
rect 34905 70825 34951 70871
rect 35009 70825 35055 70871
rect 35113 70825 35159 70871
rect 35217 70825 35263 70871
rect 35321 70825 35367 70871
rect 35425 70825 35471 70871
rect 35529 70825 35575 70871
rect 35633 70825 35679 70871
rect 35737 70825 35783 70871
rect 35841 70825 35887 70871
rect 35945 70825 35991 70871
rect 36049 70825 36095 70871
rect 36153 70825 36199 70871
rect 36257 70825 36303 70871
rect 36361 70825 36407 70871
rect 36465 70825 36511 70871
rect 36569 70825 36615 70871
rect 36673 70825 36719 70871
rect 36777 70825 36823 70871
rect 36881 70825 36927 70871
rect 36985 70825 37031 70871
rect 37089 70825 37135 70871
rect 37193 70825 37239 70871
rect 37297 70825 37343 70871
rect 37401 70825 37447 70871
rect 37505 70825 37551 70871
rect 37609 70825 37655 70871
rect 37713 70825 37759 70871
rect 37817 70825 37863 70871
rect 37921 70825 37967 70871
rect 38025 70825 38071 70871
rect 38129 70825 38175 70871
rect 38233 70825 38279 70871
rect 38337 70825 38383 70871
rect 38441 70825 38487 70871
rect 38545 70825 38591 70871
rect 38649 70825 38695 70871
rect 38753 70825 38799 70871
rect 38857 70825 38903 70871
rect 38961 70825 39007 70871
rect 39065 70825 39111 70871
rect 39169 70825 39215 70871
rect 39273 70825 39319 70871
rect 39377 70825 39423 70871
rect 39481 70825 39527 70871
rect 39585 70825 39631 70871
rect 39689 70825 39735 70871
rect 39793 70825 39839 70871
rect 39897 70825 39943 70871
rect 40001 70825 40047 70871
rect 40105 70825 40151 70871
rect 40209 70825 40255 70871
rect 40313 70825 40359 70871
rect 40417 70825 40463 70871
rect 40521 70825 40567 70871
rect 40625 70825 40671 70871
rect 40729 70825 40775 70871
rect 40833 70825 40879 70871
rect 40937 70825 40983 70871
rect 41041 70825 41087 70871
rect 41145 70825 41191 70871
rect 41249 70825 41295 70871
rect 41353 70825 41399 70871
rect 41457 70825 41503 70871
rect 41561 70825 41607 70871
rect 41665 70825 41711 70871
rect 41769 70825 41815 70871
rect 41873 70825 41919 70871
rect 41977 70825 42023 70871
rect 42081 70825 42127 70871
rect 42185 70825 42231 70871
rect 42289 70825 42335 70871
rect 42393 70825 42439 70871
rect 42497 70825 42543 70871
rect 42601 70825 42647 70871
rect 42705 70825 42751 70871
rect 42809 70825 42855 70871
rect 42913 70825 42959 70871
rect 43017 70825 43063 70871
rect 43121 70825 43167 70871
rect 43225 70825 43271 70871
rect 43329 70825 43375 70871
rect 43433 70825 43479 70871
rect 43537 70825 43583 70871
rect 43641 70825 43687 70871
rect 43745 70825 43791 70871
rect 43849 70825 43895 70871
rect 43953 70825 43999 70871
rect 44057 70825 44103 70871
rect 44161 70825 44207 70871
rect 44265 70825 44311 70871
rect 44369 70825 44415 70871
rect 44473 70825 44519 70871
rect 44577 70825 44623 70871
rect 44681 70825 44727 70871
rect 44785 70825 44831 70871
rect 44889 70825 44935 70871
rect 44993 70825 45039 70871
rect 45097 70825 45143 70871
rect 45201 70825 45247 70871
rect 45305 70825 45351 70871
rect 45409 70825 45455 70871
rect 45513 70825 45559 70871
rect 45617 70825 45663 70871
rect 45721 70825 45767 70871
rect 45825 70825 45871 70871
rect 45929 70825 45975 70871
rect 46033 70825 46079 70871
rect 46137 70825 46183 70871
rect 46241 70825 46287 70871
rect 46345 70825 46391 70871
rect 46449 70825 46495 70871
rect 46553 70825 46599 70871
rect 46657 70825 46703 70871
rect 46761 70825 46807 70871
rect 46865 70825 46911 70871
rect 46969 70825 47015 70871
rect 47073 70825 47119 70871
rect 47177 70825 47223 70871
rect 47281 70825 47327 70871
rect 47385 70825 47431 70871
rect 47489 70825 47535 70871
rect 47593 70825 47639 70871
rect 47697 70825 47743 70871
rect 47801 70825 47847 70871
rect 47905 70825 47951 70871
rect 48009 70825 48055 70871
rect 48113 70825 48159 70871
rect 48217 70825 48263 70871
rect 48321 70825 48367 70871
rect 48425 70825 48471 70871
rect 48529 70825 48575 70871
rect 48633 70825 48679 70871
rect 48737 70825 48783 70871
rect 48841 70825 48887 70871
rect 48945 70825 48991 70871
rect 49049 70825 49095 70871
rect 49153 70825 49199 70871
rect 49257 70825 49303 70871
rect 49361 70825 49407 70871
rect 49465 70825 49511 70871
rect 49569 70825 49615 70871
rect 49673 70825 49719 70871
rect 49777 70825 49823 70871
rect 49881 70825 49927 70871
rect 49985 70825 50031 70871
rect 50089 70825 50135 70871
rect 50193 70825 50239 70871
rect 50297 70825 50343 70871
rect 50401 70825 50447 70871
rect 50505 70825 50551 70871
rect 50609 70825 50655 70871
rect 50713 70825 50759 70871
rect 50817 70825 50863 70871
rect 50921 70825 50967 70871
rect 51025 70825 51071 70871
rect 51129 70825 51175 70871
rect 51233 70825 51279 70871
rect 51337 70825 51383 70871
rect 51441 70825 51487 70871
rect 51545 70825 51591 70871
rect 51649 70825 51695 70871
rect 51753 70825 51799 70871
rect 51857 70825 51903 70871
rect 51961 70825 52007 70871
rect 52065 70825 52111 70871
rect 52169 70825 52215 70871
rect 52273 70825 52319 70871
rect 52377 70825 52423 70871
rect 52481 70825 52527 70871
rect 52585 70825 52631 70871
rect 52689 70825 52735 70871
rect 52793 70825 52839 70871
rect 52897 70825 52943 70871
rect 53001 70825 53047 70871
rect 53105 70825 53151 70871
rect 53209 70825 53255 70871
rect 53313 70825 53359 70871
rect 53417 70825 53463 70871
rect 53521 70825 53567 70871
rect 53625 70825 53671 70871
rect 53729 70825 53775 70871
rect 53833 70825 53879 70871
rect 53937 70825 53983 70871
rect 54041 70825 54087 70871
rect 54145 70825 54191 70871
rect 54249 70825 54295 70871
rect 54353 70825 54399 70871
rect 54457 70825 54503 70871
rect 54561 70825 54607 70871
rect 54665 70825 54711 70871
rect 54769 70825 54815 70871
rect 54873 70825 54919 70871
rect 54977 70825 55023 70871
rect 55081 70825 55127 70871
rect 55185 70825 55231 70871
rect 55289 70825 55335 70871
rect 55393 70825 55439 70871
rect 55497 70825 55543 70871
rect 55601 70825 55647 70871
rect 55705 70825 55751 70871
rect 55809 70825 55855 70871
rect 55913 70825 55959 70871
rect 56017 70825 56063 70871
rect 56121 70825 56167 70871
rect 56225 70825 56271 70871
rect 56329 70825 56375 70871
rect 56433 70825 56479 70871
rect 56537 70825 56583 70871
rect 56641 70825 56687 70871
rect 56745 70825 56791 70871
rect 56849 70825 56895 70871
rect 56953 70825 56999 70871
rect 57057 70825 57103 70871
rect 57161 70825 57207 70871
rect 57265 70825 57311 70871
rect 57369 70825 57415 70871
rect 57473 70825 57519 70871
rect 57577 70825 57623 70871
rect 57681 70825 57727 70871
rect 57785 70825 57831 70871
rect 57889 70825 57935 70871
rect 57993 70825 58039 70871
rect 58097 70825 58143 70871
rect 58201 70825 58247 70871
rect 58305 70825 58351 70871
rect 58409 70825 58455 70871
rect 58513 70825 58559 70871
rect 58617 70825 58663 70871
rect 58721 70825 58767 70871
rect 58825 70825 58871 70871
rect 58929 70825 58975 70871
rect 59033 70825 59079 70871
rect 59137 70825 59183 70871
rect 59241 70825 59287 70871
rect 59345 70825 59391 70871
rect 59449 70825 59495 70871
rect 59553 70825 59599 70871
rect 59657 70825 59703 70871
rect 59761 70825 59807 70871
rect 59865 70825 59911 70871
rect 59969 70825 60015 70871
rect 60073 70825 60119 70871
rect 60177 70825 60223 70871
rect 60281 70825 60327 70871
rect 60385 70825 60431 70871
rect 60489 70825 60535 70871
rect 60593 70825 60639 70871
rect 60697 70825 60743 70871
rect 60801 70825 60847 70871
rect 60905 70825 60951 70871
rect 61009 70825 61055 70871
rect 61113 70825 61159 70871
rect 61217 70825 61263 70871
rect 61321 70825 61367 70871
rect 61425 70825 61471 70871
rect 61529 70825 61575 70871
rect 61633 70825 61679 70871
rect 61737 70825 61783 70871
rect 61841 70825 61887 70871
rect 61945 70825 61991 70871
rect 62049 70825 62095 70871
rect 62153 70825 62199 70871
rect 62257 70825 62303 70871
rect 62361 70825 62407 70871
rect 62465 70825 62511 70871
rect 62569 70825 62615 70871
rect 62673 70825 62719 70871
rect 62777 70825 62823 70871
rect 62881 70825 62927 70871
rect 62985 70825 63031 70871
rect 63089 70825 63135 70871
rect 63193 70825 63239 70871
rect 63297 70825 63343 70871
rect 63401 70825 63447 70871
rect 63505 70825 63551 70871
rect 63609 70825 63655 70871
rect 63713 70825 63759 70871
rect 63817 70825 63863 70871
rect 63921 70825 63967 70871
rect 64025 70825 64071 70871
rect 64129 70825 64175 70871
rect 64233 70825 64279 70871
rect 64337 70825 64383 70871
rect 64441 70825 64487 70871
rect 64545 70825 64591 70871
rect 64649 70825 64695 70871
rect 64753 70825 64799 70871
rect 64857 70825 64903 70871
rect 64961 70825 65007 70871
rect 65065 70825 65111 70871
rect 65169 70825 65215 70871
rect 65273 70825 65319 70871
rect 65377 70825 65423 70871
rect 65481 70825 65527 70871
rect 65585 70825 65631 70871
rect 65689 70825 65735 70871
rect 65793 70825 65839 70871
rect 65897 70825 65943 70871
rect 66001 70825 66047 70871
rect 66105 70825 66151 70871
rect 66209 70825 66255 70871
rect 66313 70825 66359 70871
rect 66417 70825 66463 70871
rect 66521 70825 66567 70871
rect 66625 70825 66671 70871
rect 66729 70825 66775 70871
rect 66833 70825 66879 70871
rect 66937 70825 66983 70871
rect 67041 70825 67087 70871
rect 67145 70825 67191 70871
rect 67249 70825 67295 70871
rect 67353 70825 67399 70871
rect 67457 70825 67503 70871
rect 67561 70825 67607 70871
rect 67665 70825 67711 70871
rect 67769 70825 67815 70871
rect 67873 70825 67919 70871
rect 67977 70825 68023 70871
rect 68081 70825 68127 70871
rect 68185 70825 68231 70871
rect 68289 70825 68335 70871
rect 68393 70825 68439 70871
rect 68497 70825 68543 70871
rect 68601 70825 68647 70871
rect 68705 70825 68751 70871
rect 68809 70825 68855 70871
rect 68913 70825 68959 70871
rect 69017 70825 69063 70871
rect 69121 70825 69167 70871
rect 69225 70825 69271 70871
rect 69329 70825 69375 70871
rect 69433 70825 69479 70871
rect 69537 70825 69583 70871
rect 69641 70825 69687 70871
rect 69745 70825 69791 70871
rect 69849 70825 69895 70871
rect 13119 70721 13165 70767
rect 13223 70721 13269 70767
rect 13119 70617 13165 70663
rect 13223 70617 13269 70663
rect 13119 70513 13165 70559
rect 13223 70513 13269 70559
rect 13119 70409 13165 70455
rect 13223 70409 13269 70455
rect 13119 70305 13165 70351
rect 13223 70305 13269 70351
rect 13119 70201 13165 70247
rect 13223 70201 13269 70247
rect 13119 70097 13165 70143
rect 13223 70097 13269 70143
rect 13119 69993 13165 70039
rect 13223 69993 13269 70039
rect 13119 69889 13165 69935
rect 13223 69889 13269 69935
rect 13119 69785 13165 69831
rect 13223 69785 13269 69831
rect 69796 70674 69842 70720
rect 69900 70674 69946 70720
rect 69796 70570 69842 70616
rect 69900 70570 69946 70616
rect 69796 70466 69842 70512
rect 69900 70466 69946 70512
rect 69796 70362 69842 70408
rect 69900 70362 69946 70408
rect 69796 70258 69842 70304
rect 69900 70258 69946 70304
rect 69796 70154 69842 70200
rect 69900 70154 69946 70200
rect 69796 70050 69842 70096
rect 69900 70050 69946 70096
rect 69796 69900 69842 69946
rect 69900 69900 69946 69946
rect 70004 69900 70050 69946
rect 70108 69900 70154 69946
rect 70212 69900 70258 69946
rect 70316 69900 70362 69946
rect 70420 69900 70466 69946
rect 70524 69900 70570 69946
rect 70628 69900 70674 69946
rect 70824 69862 70870 69908
rect 70928 69862 70974 69908
rect 69796 69796 69842 69842
rect 69900 69796 69946 69842
rect 70004 69796 70050 69842
rect 70108 69796 70154 69842
rect 70212 69796 70258 69842
rect 70316 69796 70362 69842
rect 70420 69796 70466 69842
rect 70524 69796 70570 69842
rect 70628 69796 70674 69842
rect 13119 69681 13165 69727
rect 13223 69681 13269 69727
rect 13119 69577 13165 69623
rect 13223 69577 13269 69623
rect 13119 69473 13165 69519
rect 13223 69473 13269 69519
rect 13119 69369 13165 69415
rect 13223 69369 13269 69415
rect 13119 69265 13165 69311
rect 13223 69265 13269 69311
rect 13119 69161 13165 69207
rect 13223 69161 13269 69207
rect 13119 69057 13165 69103
rect 13223 69057 13269 69103
rect 13119 68953 13165 68999
rect 13223 68953 13269 68999
rect 13119 68849 13165 68895
rect 13223 68849 13269 68895
rect 13119 68745 13165 68791
rect 13223 68745 13269 68791
rect 13119 68641 13165 68687
rect 13223 68641 13269 68687
rect 13119 68537 13165 68583
rect 13223 68537 13269 68583
rect 13119 68433 13165 68479
rect 13223 68433 13269 68479
rect 13119 68329 13165 68375
rect 13223 68329 13269 68375
rect 13119 68225 13165 68271
rect 13223 68225 13269 68271
rect 13119 68121 13165 68167
rect 13223 68121 13269 68167
rect 13119 68017 13165 68063
rect 13223 68017 13269 68063
rect 13119 67913 13165 67959
rect 13223 67913 13269 67959
rect 13119 67809 13165 67855
rect 13223 67809 13269 67855
rect 13119 67705 13165 67751
rect 13223 67705 13269 67751
rect 13119 67601 13165 67647
rect 13223 67601 13269 67647
rect 13119 67497 13165 67543
rect 13223 67497 13269 67543
rect 13119 67393 13165 67439
rect 13223 67393 13269 67439
rect 13119 67289 13165 67335
rect 13223 67289 13269 67335
rect 13119 67185 13165 67231
rect 13223 67185 13269 67231
rect 13119 67081 13165 67127
rect 13223 67081 13269 67127
rect 13119 66977 13165 67023
rect 13223 66977 13269 67023
rect 13119 66873 13165 66919
rect 13223 66873 13269 66919
rect 13119 66769 13165 66815
rect 13223 66769 13269 66815
rect 13119 66665 13165 66711
rect 13223 66665 13269 66711
rect 13119 66561 13165 66607
rect 13223 66561 13269 66607
rect 13119 66457 13165 66503
rect 13223 66457 13269 66503
rect 13119 66353 13165 66399
rect 13223 66353 13269 66399
rect 13119 66249 13165 66295
rect 13223 66249 13269 66295
rect 13119 66145 13165 66191
rect 13223 66145 13269 66191
rect 13119 66041 13165 66087
rect 13223 66041 13269 66087
rect 13119 65937 13165 65983
rect 13223 65937 13269 65983
rect 13119 65833 13165 65879
rect 13223 65833 13269 65879
rect 13119 65729 13165 65775
rect 13223 65729 13269 65775
rect 13119 65625 13165 65671
rect 13223 65625 13269 65671
rect 13119 65521 13165 65567
rect 13223 65521 13269 65567
rect 13119 65417 13165 65463
rect 13223 65417 13269 65463
rect 13119 65313 13165 65359
rect 13223 65313 13269 65359
rect 13119 65209 13165 65255
rect 13223 65209 13269 65255
rect 13119 65105 13165 65151
rect 13223 65105 13269 65151
rect 13119 65001 13165 65047
rect 13223 65001 13269 65047
rect 13119 64897 13165 64943
rect 13223 64897 13269 64943
rect 13119 64793 13165 64839
rect 13223 64793 13269 64839
rect 13119 64689 13165 64735
rect 13223 64689 13269 64735
rect 13119 64585 13165 64631
rect 13223 64585 13269 64631
rect 13119 64481 13165 64527
rect 13223 64481 13269 64527
rect 13119 64377 13165 64423
rect 13223 64377 13269 64423
rect 13119 64273 13165 64319
rect 13223 64273 13269 64319
rect 13119 64169 13165 64215
rect 13223 64169 13269 64215
rect 13119 64065 13165 64111
rect 13223 64065 13269 64111
rect 13119 63961 13165 64007
rect 13223 63961 13269 64007
rect 13119 63857 13165 63903
rect 13223 63857 13269 63903
rect 13119 63753 13165 63799
rect 13223 63753 13269 63799
rect 13119 63649 13165 63695
rect 13223 63649 13269 63695
rect 13119 63545 13165 63591
rect 13223 63545 13269 63591
rect 13119 63441 13165 63487
rect 13223 63441 13269 63487
rect 13119 63337 13165 63383
rect 13223 63337 13269 63383
rect 13119 63233 13165 63279
rect 13223 63233 13269 63279
rect 13119 63129 13165 63175
rect 13223 63129 13269 63175
rect 13119 63025 13165 63071
rect 13223 63025 13269 63071
rect 13119 62921 13165 62967
rect 13223 62921 13269 62967
rect 13119 62817 13165 62863
rect 13223 62817 13269 62863
rect 13119 62713 13165 62759
rect 13223 62713 13269 62759
rect 13119 62609 13165 62655
rect 13223 62609 13269 62655
rect 13119 62505 13165 62551
rect 13223 62505 13269 62551
rect 13119 62401 13165 62447
rect 13223 62401 13269 62447
rect 13119 62297 13165 62343
rect 13223 62297 13269 62343
rect 13119 62193 13165 62239
rect 13223 62193 13269 62239
rect 13119 62089 13165 62135
rect 13223 62089 13269 62135
rect 13119 61985 13165 62031
rect 13223 61985 13269 62031
rect 13119 61881 13165 61927
rect 13223 61881 13269 61927
rect 13119 61777 13165 61823
rect 13223 61777 13269 61823
rect 13119 61673 13165 61719
rect 13223 61673 13269 61719
rect 13119 61569 13165 61615
rect 13223 61569 13269 61615
rect 13119 61465 13165 61511
rect 13223 61465 13269 61511
rect 13119 61361 13165 61407
rect 13223 61361 13269 61407
rect 13119 61257 13165 61303
rect 13223 61257 13269 61303
rect 13119 61153 13165 61199
rect 13223 61153 13269 61199
rect 13119 61049 13165 61095
rect 13223 61049 13269 61095
rect 13119 60945 13165 60991
rect 13223 60945 13269 60991
rect 13119 60841 13165 60887
rect 13223 60841 13269 60887
rect 13119 60737 13165 60783
rect 13223 60737 13269 60783
rect 13119 60633 13165 60679
rect 13223 60633 13269 60679
rect 13119 60529 13165 60575
rect 13223 60529 13269 60575
rect 13119 60425 13165 60471
rect 13223 60425 13269 60471
rect 13119 60321 13165 60367
rect 13223 60321 13269 60367
rect 13119 60217 13165 60263
rect 13223 60217 13269 60263
rect 13119 60113 13165 60159
rect 13223 60113 13269 60159
rect 13119 60009 13165 60055
rect 13223 60009 13269 60055
rect 13119 59905 13165 59951
rect 13223 59905 13269 59951
rect 13119 59801 13165 59847
rect 13223 59801 13269 59847
rect 13119 59697 13165 59743
rect 13223 59697 13269 59743
rect 13119 59593 13165 59639
rect 13223 59593 13269 59639
rect 13119 59489 13165 59535
rect 13223 59489 13269 59535
rect 13119 59385 13165 59431
rect 13223 59385 13269 59431
rect 13119 59281 13165 59327
rect 13223 59281 13269 59327
rect 13119 59177 13165 59223
rect 13223 59177 13269 59223
rect 13119 59073 13165 59119
rect 13223 59073 13269 59119
rect 13119 58969 13165 59015
rect 13223 58969 13269 59015
rect 13119 58865 13165 58911
rect 13223 58865 13269 58911
rect 13119 58761 13165 58807
rect 13223 58761 13269 58807
rect 13119 58657 13165 58703
rect 13223 58657 13269 58703
rect 13119 58553 13165 58599
rect 13223 58553 13269 58599
rect 13119 58449 13165 58495
rect 13223 58449 13269 58495
rect 13119 58345 13165 58391
rect 13223 58345 13269 58391
rect 13119 58241 13165 58287
rect 13223 58241 13269 58287
rect 13119 58137 13165 58183
rect 13223 58137 13269 58183
rect 13119 58033 13165 58079
rect 13223 58033 13269 58079
rect 13119 57929 13165 57975
rect 13223 57929 13269 57975
rect 13119 57825 13165 57871
rect 13223 57825 13269 57871
rect 13119 57721 13165 57767
rect 13223 57721 13269 57767
rect 13119 57617 13165 57663
rect 13223 57617 13269 57663
rect 13119 57513 13165 57559
rect 13223 57513 13269 57559
rect 13119 57409 13165 57455
rect 13223 57409 13269 57455
rect 13119 57305 13165 57351
rect 13223 57305 13269 57351
rect 13119 57201 13165 57247
rect 13223 57201 13269 57247
rect 13119 57097 13165 57143
rect 13223 57097 13269 57143
rect 13119 56993 13165 57039
rect 13223 56993 13269 57039
rect 13119 56889 13165 56935
rect 13223 56889 13269 56935
rect 13119 56785 13165 56831
rect 13223 56785 13269 56831
rect 13119 56681 13165 56727
rect 13223 56681 13269 56727
rect 13119 56577 13165 56623
rect 13223 56577 13269 56623
rect 13119 56473 13165 56519
rect 13223 56473 13269 56519
rect 13119 56369 13165 56415
rect 13223 56369 13269 56415
rect 13119 56265 13165 56311
rect 13223 56265 13269 56311
rect 13119 56161 13165 56207
rect 13223 56161 13269 56207
rect 13119 56057 13165 56103
rect 13223 56057 13269 56103
rect 13119 55953 13165 55999
rect 13223 55953 13269 55999
rect 13119 55849 13165 55895
rect 13223 55849 13269 55895
rect 13119 55745 13165 55791
rect 13223 55745 13269 55791
rect 13119 55641 13165 55687
rect 13223 55641 13269 55687
rect 13119 55537 13165 55583
rect 13223 55537 13269 55583
rect 13119 55433 13165 55479
rect 13223 55433 13269 55479
rect 13119 55329 13165 55375
rect 13223 55329 13269 55375
rect 13119 55225 13165 55271
rect 13223 55225 13269 55271
rect 13119 55121 13165 55167
rect 13223 55121 13269 55167
rect 13119 55017 13165 55063
rect 13223 55017 13269 55063
rect 13119 54913 13165 54959
rect 13223 54913 13269 54959
rect 13119 54809 13165 54855
rect 13223 54809 13269 54855
rect 13119 54705 13165 54751
rect 13223 54705 13269 54751
rect 13119 54601 13165 54647
rect 13223 54601 13269 54647
rect 13119 54497 13165 54543
rect 13223 54497 13269 54543
rect 13119 54393 13165 54439
rect 13223 54393 13269 54439
rect 13119 54289 13165 54335
rect 13223 54289 13269 54335
rect 13119 54185 13165 54231
rect 13223 54185 13269 54231
rect 13119 54081 13165 54127
rect 13223 54081 13269 54127
rect 13119 53977 13165 54023
rect 13223 53977 13269 54023
rect 13119 53873 13165 53919
rect 13223 53873 13269 53919
rect 13119 53769 13165 53815
rect 13223 53769 13269 53815
rect 13119 53665 13165 53711
rect 13223 53665 13269 53711
rect 13119 53561 13165 53607
rect 13223 53561 13269 53607
rect 13119 53457 13165 53503
rect 13223 53457 13269 53503
rect 13119 53353 13165 53399
rect 13223 53353 13269 53399
rect 13119 53249 13165 53295
rect 13223 53249 13269 53295
rect 13119 53145 13165 53191
rect 13223 53145 13269 53191
rect 13119 53041 13165 53087
rect 13223 53041 13269 53087
rect 13119 52937 13165 52983
rect 13223 52937 13269 52983
rect 13119 52833 13165 52879
rect 13223 52833 13269 52879
rect 13119 52729 13165 52775
rect 13223 52729 13269 52775
rect 13119 52625 13165 52671
rect 13223 52625 13269 52671
rect 13119 52521 13165 52567
rect 13223 52521 13269 52567
rect 13119 52417 13165 52463
rect 13223 52417 13269 52463
rect 13119 52313 13165 52359
rect 13223 52313 13269 52359
rect 13119 52209 13165 52255
rect 13223 52209 13269 52255
rect 13119 52105 13165 52151
rect 13223 52105 13269 52151
rect 13119 52001 13165 52047
rect 13223 52001 13269 52047
rect 13119 51897 13165 51943
rect 13223 51897 13269 51943
rect 13119 51793 13165 51839
rect 13223 51793 13269 51839
rect 13119 51689 13165 51735
rect 13223 51689 13269 51735
rect 13119 51585 13165 51631
rect 13223 51585 13269 51631
rect 13119 51481 13165 51527
rect 13223 51481 13269 51527
rect 13119 51377 13165 51423
rect 13223 51377 13269 51423
rect 13119 51273 13165 51319
rect 13223 51273 13269 51319
rect 13119 51169 13165 51215
rect 13223 51169 13269 51215
rect 13119 51065 13165 51111
rect 13223 51065 13269 51111
rect 13119 50961 13165 51007
rect 13223 50961 13269 51007
rect 13119 50857 13165 50903
rect 13223 50857 13269 50903
rect 13119 50753 13165 50799
rect 13223 50753 13269 50799
rect 13119 50649 13165 50695
rect 13223 50649 13269 50695
rect 13119 50545 13165 50591
rect 13223 50545 13269 50591
rect 13119 50441 13165 50487
rect 13223 50441 13269 50487
rect 13119 50337 13165 50383
rect 13223 50337 13269 50383
rect 13119 50233 13165 50279
rect 13223 50233 13269 50279
rect 13119 50129 13165 50175
rect 13223 50129 13269 50175
rect 13119 50025 13165 50071
rect 13223 50025 13269 50071
rect 13119 49921 13165 49967
rect 13223 49921 13269 49967
rect 13119 49817 13165 49863
rect 13223 49817 13269 49863
rect 13119 49713 13165 49759
rect 13223 49713 13269 49759
rect 13119 49609 13165 49655
rect 13223 49609 13269 49655
rect 13119 49505 13165 49551
rect 13223 49505 13269 49551
rect 13119 49401 13165 49447
rect 13223 49401 13269 49447
rect 13119 49297 13165 49343
rect 13223 49297 13269 49343
rect 13119 49193 13165 49239
rect 13223 49193 13269 49239
rect 13119 49089 13165 49135
rect 13223 49089 13269 49135
rect 13119 48985 13165 49031
rect 13223 48985 13269 49031
rect 13119 48881 13165 48927
rect 13223 48881 13269 48927
rect 13119 48777 13165 48823
rect 13223 48777 13269 48823
rect 13119 48673 13165 48719
rect 13223 48673 13269 48719
rect 13119 48569 13165 48615
rect 13223 48569 13269 48615
rect 13119 48465 13165 48511
rect 13223 48465 13269 48511
rect 13119 48361 13165 48407
rect 13223 48361 13269 48407
rect 13119 48257 13165 48303
rect 13223 48257 13269 48303
rect 13119 48153 13165 48199
rect 13223 48153 13269 48199
rect 13119 48049 13165 48095
rect 13223 48049 13269 48095
rect 13119 47945 13165 47991
rect 13223 47945 13269 47991
rect 13119 47841 13165 47887
rect 13223 47841 13269 47887
rect 13119 47737 13165 47783
rect 13223 47737 13269 47783
rect 13119 47633 13165 47679
rect 13223 47633 13269 47679
rect 13119 47529 13165 47575
rect 13223 47529 13269 47575
rect 13119 47425 13165 47471
rect 13223 47425 13269 47471
rect 13119 47321 13165 47367
rect 13223 47321 13269 47367
rect 13119 47217 13165 47263
rect 13223 47217 13269 47263
rect 13119 47113 13165 47159
rect 13223 47113 13269 47159
rect 13119 47009 13165 47055
rect 13223 47009 13269 47055
rect 13119 46905 13165 46951
rect 13223 46905 13269 46951
rect 13119 46801 13165 46847
rect 13223 46801 13269 46847
rect 13119 46697 13165 46743
rect 13223 46697 13269 46743
rect 13119 46593 13165 46639
rect 13223 46593 13269 46639
rect 13119 46489 13165 46535
rect 13223 46489 13269 46535
rect 13119 46385 13165 46431
rect 13223 46385 13269 46431
rect 13119 46281 13165 46327
rect 13223 46281 13269 46327
rect 13119 46177 13165 46223
rect 13223 46177 13269 46223
rect 13119 46073 13165 46119
rect 13223 46073 13269 46119
rect 13119 45969 13165 46015
rect 13223 45969 13269 46015
rect 13119 45865 13165 45911
rect 13223 45865 13269 45911
rect 13119 45761 13165 45807
rect 13223 45761 13269 45807
rect 13119 45657 13165 45703
rect 13223 45657 13269 45703
rect 13119 45553 13165 45599
rect 13223 45553 13269 45599
rect 13119 45449 13165 45495
rect 13223 45449 13269 45495
rect 13119 45345 13165 45391
rect 13223 45345 13269 45391
rect 13119 45241 13165 45287
rect 13223 45241 13269 45287
rect 13119 45137 13165 45183
rect 13223 45137 13269 45183
rect 13119 45033 13165 45079
rect 13223 45033 13269 45079
rect 70824 69758 70870 69804
rect 70928 69758 70974 69804
rect 70824 69654 70870 69700
rect 70928 69654 70974 69700
rect 70824 69550 70870 69596
rect 70928 69550 70974 69596
rect 70824 69446 70870 69492
rect 70928 69446 70974 69492
rect 70824 69342 70870 69388
rect 70928 69342 70974 69388
rect 70824 69238 70870 69284
rect 70928 69238 70974 69284
rect 70824 69134 70870 69180
rect 70928 69134 70974 69180
rect 70824 69030 70870 69076
rect 70928 69030 70974 69076
rect 70824 68926 70870 68972
rect 70928 68926 70974 68972
rect 70824 68822 70870 68868
rect 70928 68822 70974 68868
rect 70824 68718 70870 68764
rect 70928 68718 70974 68764
rect 70824 68614 70870 68660
rect 70928 68614 70974 68660
rect 70824 68510 70870 68556
rect 70928 68510 70974 68556
rect 70824 68406 70870 68452
rect 70928 68406 70974 68452
rect 70824 68302 70870 68348
rect 70928 68302 70974 68348
rect 70824 68198 70870 68244
rect 70928 68198 70974 68244
rect 70824 68094 70870 68140
rect 70928 68094 70974 68140
rect 70824 67990 70870 68036
rect 70928 67990 70974 68036
rect 70824 67886 70870 67932
rect 70928 67886 70974 67932
rect 70824 67782 70870 67828
rect 70928 67782 70974 67828
rect 70824 67678 70870 67724
rect 70928 67678 70974 67724
rect 70824 67574 70870 67620
rect 70928 67574 70974 67620
rect 70824 67470 70870 67516
rect 70928 67470 70974 67516
rect 70824 67366 70870 67412
rect 70928 67366 70974 67412
rect 70824 67262 70870 67308
rect 70928 67262 70974 67308
rect 70824 67158 70870 67204
rect 70928 67158 70974 67204
rect 70824 67054 70870 67100
rect 70928 67054 70974 67100
rect 70824 66950 70870 66996
rect 70928 66950 70974 66996
rect 70824 66846 70870 66892
rect 70928 66846 70974 66892
rect 70824 66742 70870 66788
rect 70928 66742 70974 66788
rect 70824 66638 70870 66684
rect 70928 66638 70974 66684
rect 70824 66534 70870 66580
rect 70928 66534 70974 66580
rect 70824 66430 70870 66476
rect 70928 66430 70974 66476
rect 70824 66326 70870 66372
rect 70928 66326 70974 66372
rect 70824 66222 70870 66268
rect 70928 66222 70974 66268
rect 70824 66118 70870 66164
rect 70928 66118 70974 66164
rect 70824 66014 70870 66060
rect 70928 66014 70974 66060
rect 70824 65910 70870 65956
rect 70928 65910 70974 65956
rect 70824 65806 70870 65852
rect 70928 65806 70974 65852
rect 70824 65702 70870 65748
rect 70928 65702 70974 65748
rect 70824 65598 70870 65644
rect 70928 65598 70974 65644
rect 70824 65494 70870 65540
rect 70928 65494 70974 65540
rect 70824 65390 70870 65436
rect 70928 65390 70974 65436
rect 70824 65286 70870 65332
rect 70928 65286 70974 65332
rect 70824 65182 70870 65228
rect 70928 65182 70974 65228
rect 70824 65078 70870 65124
rect 70928 65078 70974 65124
rect 70824 64974 70870 65020
rect 70928 64974 70974 65020
rect 70824 64870 70870 64916
rect 70928 64870 70974 64916
rect 70824 64766 70870 64812
rect 70928 64766 70974 64812
rect 70824 64662 70870 64708
rect 70928 64662 70974 64708
rect 70824 64558 70870 64604
rect 70928 64558 70974 64604
rect 70824 64454 70870 64500
rect 70928 64454 70974 64500
rect 70824 64350 70870 64396
rect 70928 64350 70974 64396
rect 70824 64246 70870 64292
rect 70928 64246 70974 64292
rect 70824 64142 70870 64188
rect 70928 64142 70974 64188
rect 70824 64038 70870 64084
rect 70928 64038 70974 64084
rect 70824 63934 70870 63980
rect 70928 63934 70974 63980
rect 70824 63830 70870 63876
rect 70928 63830 70974 63876
rect 70824 63726 70870 63772
rect 70928 63726 70974 63772
rect 70824 63622 70870 63668
rect 70928 63622 70974 63668
rect 70824 63518 70870 63564
rect 70928 63518 70974 63564
rect 70824 63414 70870 63460
rect 70928 63414 70974 63460
rect 70824 63310 70870 63356
rect 70928 63310 70974 63356
rect 70824 63206 70870 63252
rect 70928 63206 70974 63252
rect 70824 63102 70870 63148
rect 70928 63102 70974 63148
rect 70824 62998 70870 63044
rect 70928 62998 70974 63044
rect 70824 62894 70870 62940
rect 70928 62894 70974 62940
rect 70824 62790 70870 62836
rect 70928 62790 70974 62836
rect 70824 62686 70870 62732
rect 70928 62686 70974 62732
rect 70824 62582 70870 62628
rect 70928 62582 70974 62628
rect 70824 62478 70870 62524
rect 70928 62478 70974 62524
rect 70824 62374 70870 62420
rect 70928 62374 70974 62420
rect 70824 62270 70870 62316
rect 70928 62270 70974 62316
rect 70824 62166 70870 62212
rect 70928 62166 70974 62212
rect 70824 62062 70870 62108
rect 70928 62062 70974 62108
rect 70824 61958 70870 62004
rect 70928 61958 70974 62004
rect 70824 61854 70870 61900
rect 70928 61854 70974 61900
rect 70824 61750 70870 61796
rect 70928 61750 70974 61796
rect 70824 61646 70870 61692
rect 70928 61646 70974 61692
rect 70824 61542 70870 61588
rect 70928 61542 70974 61588
rect 70824 61438 70870 61484
rect 70928 61438 70974 61484
rect 70824 61334 70870 61380
rect 70928 61334 70974 61380
rect 70824 61230 70870 61276
rect 70928 61230 70974 61276
rect 70824 61126 70870 61172
rect 70928 61126 70974 61172
rect 70824 61022 70870 61068
rect 70928 61022 70974 61068
rect 70824 60918 70870 60964
rect 70928 60918 70974 60964
rect 70824 60814 70870 60860
rect 70928 60814 70974 60860
rect 70824 60710 70870 60756
rect 70928 60710 70974 60756
rect 70824 60606 70870 60652
rect 70928 60606 70974 60652
rect 70824 60502 70870 60548
rect 70928 60502 70974 60548
rect 70824 60398 70870 60444
rect 70928 60398 70974 60444
rect 70824 60294 70870 60340
rect 70928 60294 70974 60340
rect 70824 60190 70870 60236
rect 70928 60190 70974 60236
rect 70824 60086 70870 60132
rect 70928 60086 70974 60132
rect 70824 59982 70870 60028
rect 70928 59982 70974 60028
rect 70824 59878 70870 59924
rect 70928 59878 70974 59924
rect 70824 59774 70870 59820
rect 70928 59774 70974 59820
rect 70824 59670 70870 59716
rect 70928 59670 70974 59716
rect 70824 59566 70870 59612
rect 70928 59566 70974 59612
rect 70824 59462 70870 59508
rect 70928 59462 70974 59508
rect 70824 59358 70870 59404
rect 70928 59358 70974 59404
rect 70824 59254 70870 59300
rect 70928 59254 70974 59300
rect 70824 59150 70870 59196
rect 70928 59150 70974 59196
rect 70824 59046 70870 59092
rect 70928 59046 70974 59092
rect 70824 58942 70870 58988
rect 70928 58942 70974 58988
rect 70824 58838 70870 58884
rect 70928 58838 70974 58884
rect 70824 58734 70870 58780
rect 70928 58734 70974 58780
rect 70824 58630 70870 58676
rect 70928 58630 70974 58676
rect 70824 58526 70870 58572
rect 70928 58526 70974 58572
rect 70824 58422 70870 58468
rect 70928 58422 70974 58468
rect 70824 58318 70870 58364
rect 70928 58318 70974 58364
rect 70824 58214 70870 58260
rect 70928 58214 70974 58260
rect 70824 58110 70870 58156
rect 70928 58110 70974 58156
rect 70824 58006 70870 58052
rect 70928 58006 70974 58052
rect 70824 57902 70870 57948
rect 70928 57902 70974 57948
rect 70824 57798 70870 57844
rect 70928 57798 70974 57844
rect 70824 57694 70870 57740
rect 70928 57694 70974 57740
rect 70824 57590 70870 57636
rect 70928 57590 70974 57636
rect 70824 57486 70870 57532
rect 70928 57486 70974 57532
rect 70824 57382 70870 57428
rect 70928 57382 70974 57428
rect 70824 57278 70870 57324
rect 70928 57278 70974 57324
rect 70824 57174 70870 57220
rect 70928 57174 70974 57220
rect 70824 57070 70870 57116
rect 70928 57070 70974 57116
rect 70824 56966 70870 57012
rect 70928 56966 70974 57012
rect 70824 56862 70870 56908
rect 70928 56862 70974 56908
rect 70824 56758 70870 56804
rect 70928 56758 70974 56804
rect 70824 56654 70870 56700
rect 70928 56654 70974 56700
rect 70824 56550 70870 56596
rect 70928 56550 70974 56596
rect 70824 56446 70870 56492
rect 70928 56446 70974 56492
rect 70824 56342 70870 56388
rect 70928 56342 70974 56388
rect 70824 56238 70870 56284
rect 70928 56238 70974 56284
rect 70824 56134 70870 56180
rect 70928 56134 70974 56180
rect 70824 56030 70870 56076
rect 70928 56030 70974 56076
rect 70824 55926 70870 55972
rect 70928 55926 70974 55972
rect 70824 55822 70870 55868
rect 70928 55822 70974 55868
rect 70824 55718 70870 55764
rect 70928 55718 70974 55764
rect 70824 55614 70870 55660
rect 70928 55614 70974 55660
rect 70824 55510 70870 55556
rect 70928 55510 70974 55556
rect 70824 55406 70870 55452
rect 70928 55406 70974 55452
rect 70824 55302 70870 55348
rect 70928 55302 70974 55348
rect 70824 55198 70870 55244
rect 70928 55198 70974 55244
rect 70824 55094 70870 55140
rect 70928 55094 70974 55140
rect 70824 54990 70870 55036
rect 70928 54990 70974 55036
rect 70824 54886 70870 54932
rect 70928 54886 70974 54932
rect 70824 54782 70870 54828
rect 70928 54782 70974 54828
rect 70824 54678 70870 54724
rect 70928 54678 70974 54724
rect 70824 54574 70870 54620
rect 70928 54574 70974 54620
rect 70824 54470 70870 54516
rect 70928 54470 70974 54516
rect 70824 54366 70870 54412
rect 70928 54366 70974 54412
rect 70824 54262 70870 54308
rect 70928 54262 70974 54308
rect 70824 54158 70870 54204
rect 70928 54158 70974 54204
rect 70824 54054 70870 54100
rect 70928 54054 70974 54100
rect 70824 53950 70870 53996
rect 70928 53950 70974 53996
rect 70824 53846 70870 53892
rect 70928 53846 70974 53892
rect 70824 53742 70870 53788
rect 70928 53742 70974 53788
rect 70824 53638 70870 53684
rect 70928 53638 70974 53684
rect 70824 53534 70870 53580
rect 70928 53534 70974 53580
rect 70824 53430 70870 53476
rect 70928 53430 70974 53476
rect 70824 53326 70870 53372
rect 70928 53326 70974 53372
rect 70824 53222 70870 53268
rect 70928 53222 70974 53268
rect 70824 53118 70870 53164
rect 70928 53118 70974 53164
rect 70824 53014 70870 53060
rect 70928 53014 70974 53060
rect 70824 52910 70870 52956
rect 70928 52910 70974 52956
rect 70824 52806 70870 52852
rect 70928 52806 70974 52852
rect 70824 52702 70870 52748
rect 70928 52702 70974 52748
rect 70824 52598 70870 52644
rect 70928 52598 70974 52644
rect 70824 52494 70870 52540
rect 70928 52494 70974 52540
rect 70824 52390 70870 52436
rect 70928 52390 70974 52436
rect 70824 52286 70870 52332
rect 70928 52286 70974 52332
rect 70824 52182 70870 52228
rect 70928 52182 70974 52228
rect 70824 52078 70870 52124
rect 70928 52078 70974 52124
rect 70824 51974 70870 52020
rect 70928 51974 70974 52020
rect 70824 51870 70870 51916
rect 70928 51870 70974 51916
rect 70824 51766 70870 51812
rect 70928 51766 70974 51812
rect 70824 51662 70870 51708
rect 70928 51662 70974 51708
rect 70824 51558 70870 51604
rect 70928 51558 70974 51604
rect 70824 51454 70870 51500
rect 70928 51454 70974 51500
rect 70824 51350 70870 51396
rect 70928 51350 70974 51396
rect 70824 51246 70870 51292
rect 70928 51246 70974 51292
rect 70824 51142 70870 51188
rect 70928 51142 70974 51188
rect 70824 51038 70870 51084
rect 70928 51038 70974 51084
rect 70824 50934 70870 50980
rect 70928 50934 70974 50980
rect 70824 50830 70870 50876
rect 70928 50830 70974 50876
rect 70824 50726 70870 50772
rect 70928 50726 70974 50772
rect 70824 50622 70870 50668
rect 70928 50622 70974 50668
rect 70824 50518 70870 50564
rect 70928 50518 70974 50564
rect 70824 50414 70870 50460
rect 70928 50414 70974 50460
rect 70824 50310 70870 50356
rect 70928 50310 70974 50356
rect 70824 50206 70870 50252
rect 70928 50206 70974 50252
rect 70824 50102 70870 50148
rect 70928 50102 70974 50148
rect 70824 49998 70870 50044
rect 70928 49998 70974 50044
rect 70824 49894 70870 49940
rect 70928 49894 70974 49940
rect 70824 49790 70870 49836
rect 70928 49790 70974 49836
rect 70824 49686 70870 49732
rect 70928 49686 70974 49732
rect 70824 49582 70870 49628
rect 70928 49582 70974 49628
rect 70824 49478 70870 49524
rect 70928 49478 70974 49524
rect 70824 49374 70870 49420
rect 70928 49374 70974 49420
rect 70824 49270 70870 49316
rect 70928 49270 70974 49316
rect 70824 49166 70870 49212
rect 70928 49166 70974 49212
rect 70824 49062 70870 49108
rect 70928 49062 70974 49108
rect 70824 48958 70870 49004
rect 70928 48958 70974 49004
rect 70824 48854 70870 48900
rect 70928 48854 70974 48900
rect 70824 48750 70870 48796
rect 70928 48750 70974 48796
rect 70824 48646 70870 48692
rect 70928 48646 70974 48692
rect 70824 48542 70870 48588
rect 70928 48542 70974 48588
rect 70824 48438 70870 48484
rect 70928 48438 70974 48484
rect 70824 48334 70870 48380
rect 70928 48334 70974 48380
rect 70824 48230 70870 48276
rect 70928 48230 70974 48276
rect 70824 48126 70870 48172
rect 70928 48126 70974 48172
rect 70824 48022 70870 48068
rect 70928 48022 70974 48068
rect 70824 47918 70870 47964
rect 70928 47918 70974 47964
rect 70824 47814 70870 47860
rect 70928 47814 70974 47860
rect 70824 47710 70870 47756
rect 70928 47710 70974 47756
rect 70824 47606 70870 47652
rect 70928 47606 70974 47652
rect 70824 47502 70870 47548
rect 70928 47502 70974 47548
rect 70824 47398 70870 47444
rect 70928 47398 70974 47444
rect 70824 47294 70870 47340
rect 70928 47294 70974 47340
rect 70824 47190 70870 47236
rect 70928 47190 70974 47236
rect 70824 47086 70870 47132
rect 70928 47086 70974 47132
rect 70824 46982 70870 47028
rect 70928 46982 70974 47028
rect 70824 46878 70870 46924
rect 70928 46878 70974 46924
rect 70824 46774 70870 46820
rect 70928 46774 70974 46820
rect 70824 46670 70870 46716
rect 70928 46670 70974 46716
rect 70824 46566 70870 46612
rect 70928 46566 70974 46612
rect 70824 46462 70870 46508
rect 70928 46462 70974 46508
rect 70824 46358 70870 46404
rect 70928 46358 70974 46404
rect 70824 46254 70870 46300
rect 70928 46254 70974 46300
rect 70824 46150 70870 46196
rect 70928 46150 70974 46196
rect 70824 46046 70870 46092
rect 70928 46046 70974 46092
rect 70824 45942 70870 45988
rect 70928 45942 70974 45988
rect 70824 45838 70870 45884
rect 70928 45838 70974 45884
rect 70824 45734 70870 45780
rect 70928 45734 70974 45780
rect 70824 45630 70870 45676
rect 70928 45630 70974 45676
rect 70824 45526 70870 45572
rect 70928 45526 70974 45572
rect 70824 45422 70870 45468
rect 70928 45422 70974 45468
rect 70824 45318 70870 45364
rect 70928 45318 70974 45364
rect 70824 45214 70870 45260
rect 70928 45214 70974 45260
rect 70824 45110 70870 45156
rect 70928 45110 70974 45156
rect 70824 45006 70870 45052
rect 70928 45006 70974 45052
rect 70824 44902 70870 44948
rect 70928 44902 70974 44948
rect 13254 44778 13300 44824
rect 70824 44798 70870 44844
rect 70928 44798 70974 44844
rect 13386 44646 13432 44692
rect 70824 44694 70870 44740
rect 70928 44694 70974 44740
rect 70824 44590 70870 44636
rect 70928 44590 70974 44636
rect 13518 44514 13564 44560
rect 70824 44486 70870 44532
rect 70928 44486 70974 44532
rect 13650 44382 13696 44428
rect 70824 44382 70870 44428
rect 70928 44382 70974 44428
rect 13782 44250 13828 44296
rect 70824 44278 70870 44324
rect 70928 44278 70974 44324
rect 13914 44118 13960 44164
rect 70824 44174 70870 44220
rect 70928 44174 70974 44220
rect 70824 44070 70870 44116
rect 70928 44070 70974 44116
rect 14046 43986 14092 44032
rect 70824 43966 70870 44012
rect 70928 43966 70974 44012
rect 14178 43854 14224 43900
rect 70824 43862 70870 43908
rect 70928 43862 70974 43908
rect 14310 43722 14356 43768
rect 70824 43758 70870 43804
rect 70928 43758 70974 43804
rect 70824 43654 70870 43700
rect 70928 43654 70974 43700
rect 14442 43590 14488 43636
rect 70824 43550 70870 43596
rect 70928 43550 70974 43596
rect 14574 43458 14620 43504
rect 70824 43446 70870 43492
rect 70928 43446 70974 43492
rect 14706 43326 14752 43372
rect 70824 43342 70870 43388
rect 70928 43342 70974 43388
rect 14838 43194 14884 43240
rect 70824 43238 70870 43284
rect 70928 43238 70974 43284
rect 70824 43134 70870 43180
rect 70928 43134 70974 43180
rect 14970 43062 15016 43108
rect 70824 43030 70870 43076
rect 70928 43030 70974 43076
rect 15102 42930 15148 42976
rect 70824 42926 70870 42972
rect 70928 42926 70974 42972
rect 15234 42798 15280 42844
rect 70824 42822 70870 42868
rect 70928 42822 70974 42868
rect 15366 42666 15412 42712
rect 70824 42718 70870 42764
rect 70928 42718 70974 42764
rect 70824 42614 70870 42660
rect 70928 42614 70974 42660
rect 15498 42534 15544 42580
rect 70824 42510 70870 42556
rect 70928 42510 70974 42556
rect 15630 42402 15676 42448
rect 70824 42406 70870 42452
rect 70928 42406 70974 42452
rect 15762 42270 15808 42316
rect 70824 42302 70870 42348
rect 70928 42302 70974 42348
rect 15894 42138 15940 42184
rect 70824 42198 70870 42244
rect 70928 42198 70974 42244
rect 70824 42094 70870 42140
rect 70928 42094 70974 42140
rect 16026 42006 16072 42052
rect 70824 41990 70870 42036
rect 70928 41990 70974 42036
rect 16158 41874 16204 41920
rect 70824 41886 70870 41932
rect 70928 41886 70974 41932
rect 16290 41742 16336 41788
rect 70824 41782 70870 41828
rect 70928 41782 70974 41828
rect 70824 41678 70870 41724
rect 70928 41678 70974 41724
rect 16422 41610 16468 41656
rect 70824 41574 70870 41620
rect 70928 41574 70974 41620
rect 16554 41478 16600 41524
rect 70824 41470 70870 41516
rect 70928 41470 70974 41516
rect 16686 41346 16732 41392
rect 70824 41366 70870 41412
rect 70928 41366 70974 41412
rect 16818 41214 16864 41260
rect 70824 41262 70870 41308
rect 70928 41262 70974 41308
rect 70824 41158 70870 41204
rect 70928 41158 70974 41204
rect 16950 41082 16996 41128
rect 70824 41054 70870 41100
rect 70928 41054 70974 41100
rect 17082 40950 17128 40996
rect 70824 40950 70870 40996
rect 70928 40950 70974 40996
rect 17214 40818 17260 40864
rect 70824 40846 70870 40892
rect 70928 40846 70974 40892
rect 70824 40742 70870 40788
rect 70928 40742 70974 40788
rect 17346 40686 17392 40732
rect 70824 40638 70870 40684
rect 70928 40638 70974 40684
rect 17478 40554 17524 40600
rect 70824 40534 70870 40580
rect 70928 40534 70974 40580
rect 17610 40422 17656 40468
rect 70824 40430 70870 40476
rect 70928 40430 70974 40476
rect 17742 40290 17788 40336
rect 70824 40326 70870 40372
rect 70928 40326 70974 40372
rect 17874 40158 17920 40204
rect 70824 40222 70870 40268
rect 70928 40222 70974 40268
rect 70824 40118 70870 40164
rect 70928 40118 70974 40164
rect 18006 40026 18052 40072
rect 70824 40014 70870 40060
rect 70928 40014 70974 40060
rect 18138 39894 18184 39940
rect 70824 39910 70870 39956
rect 70928 39910 70974 39956
rect 18270 39762 18316 39808
rect 70824 39806 70870 39852
rect 70928 39806 70974 39852
rect 70824 39702 70870 39748
rect 70928 39702 70974 39748
rect 18402 39630 18448 39676
rect 70824 39598 70870 39644
rect 70928 39598 70974 39644
rect 18534 39498 18580 39544
rect 70824 39494 70870 39540
rect 70928 39494 70974 39540
rect 18666 39366 18712 39412
rect 70824 39390 70870 39436
rect 70928 39390 70974 39436
rect 18798 39234 18844 39280
rect 70824 39286 70870 39332
rect 70928 39286 70974 39332
rect 18930 39102 18976 39148
rect 70824 39182 70870 39228
rect 70928 39182 70974 39228
rect 70824 39078 70870 39124
rect 70928 39078 70974 39124
rect 19062 38970 19108 39016
rect 70824 38974 70870 39020
rect 70928 38974 70974 39020
rect 19194 38838 19240 38884
rect 70824 38870 70870 38916
rect 70928 38870 70974 38916
rect 70824 38766 70870 38812
rect 70928 38766 70974 38812
rect 19326 38706 19372 38752
rect 70824 38662 70870 38708
rect 70928 38662 70974 38708
rect 19458 38574 19504 38620
rect 70824 38558 70870 38604
rect 70928 38558 70974 38604
rect 19590 38442 19636 38488
rect 70824 38454 70870 38500
rect 70928 38454 70974 38500
rect 19722 38310 19768 38356
rect 70824 38350 70870 38396
rect 70928 38350 70974 38396
rect 19854 38178 19900 38224
rect 70824 38246 70870 38292
rect 70928 38246 70974 38292
rect 70824 38142 70870 38188
rect 70928 38142 70974 38188
rect 19986 38046 20032 38092
rect 70824 38038 70870 38084
rect 70928 38038 70974 38084
rect 20118 37914 20164 37960
rect 70824 37934 70870 37980
rect 70928 37934 70974 37980
rect 20250 37782 20296 37828
rect 70824 37830 70870 37876
rect 70928 37830 70974 37876
rect 70824 37726 70870 37772
rect 70928 37726 70974 37772
rect 20382 37650 20428 37696
rect 70824 37622 70870 37668
rect 70928 37622 70974 37668
rect 20514 37518 20560 37564
rect 70824 37518 70870 37564
rect 70928 37518 70974 37564
rect 20646 37386 20692 37432
rect 70824 37414 70870 37460
rect 70928 37414 70974 37460
rect 20778 37254 20824 37300
rect 70824 37310 70870 37356
rect 70928 37310 70974 37356
rect 70824 37206 70870 37252
rect 70928 37206 70974 37252
rect 20910 37122 20956 37168
rect 70824 37102 70870 37148
rect 70928 37102 70974 37148
rect 21042 36990 21088 37036
rect 70824 36998 70870 37044
rect 70928 36998 70974 37044
rect 21174 36858 21220 36904
rect 70824 36894 70870 36940
rect 70928 36894 70974 36940
rect 21306 36726 21352 36772
rect 70824 36790 70870 36836
rect 70928 36790 70974 36836
rect 70824 36686 70870 36732
rect 70928 36686 70974 36732
rect 21438 36594 21484 36640
rect 70824 36582 70870 36628
rect 70928 36582 70974 36628
rect 21570 36462 21616 36508
rect 70824 36478 70870 36524
rect 70928 36478 70974 36524
rect 21702 36330 21748 36376
rect 70824 36374 70870 36420
rect 70928 36374 70974 36420
rect 21834 36198 21880 36244
rect 70824 36270 70870 36316
rect 70928 36270 70974 36316
rect 70824 36166 70870 36212
rect 70928 36166 70974 36212
rect 21966 36066 22012 36112
rect 70824 36062 70870 36108
rect 70928 36062 70974 36108
rect 22098 35934 22144 35980
rect 70824 35958 70870 36004
rect 70928 35958 70974 36004
rect 22230 35802 22276 35848
rect 70824 35854 70870 35900
rect 70928 35854 70974 35900
rect 70824 35750 70870 35796
rect 70928 35750 70974 35796
rect 22362 35670 22408 35716
rect 70824 35646 70870 35692
rect 70928 35646 70974 35692
rect 22494 35538 22540 35584
rect 70824 35542 70870 35588
rect 70928 35542 70974 35588
rect 22626 35406 22672 35452
rect 70824 35438 70870 35484
rect 70928 35438 70974 35484
rect 22758 35274 22804 35320
rect 70824 35334 70870 35380
rect 70928 35334 70974 35380
rect 70824 35230 70870 35276
rect 70928 35230 70974 35276
rect 22890 35142 22936 35188
rect 70824 35126 70870 35172
rect 70928 35126 70974 35172
rect 23022 35010 23068 35056
rect 70824 35022 70870 35068
rect 70928 35022 70974 35068
rect 23154 34878 23200 34924
rect 70824 34918 70870 34964
rect 70928 34918 70974 34964
rect 70824 34814 70870 34860
rect 70928 34814 70974 34860
rect 23286 34746 23332 34792
rect 70824 34710 70870 34756
rect 70928 34710 70974 34756
rect 23418 34614 23464 34660
rect 70824 34606 70870 34652
rect 70928 34606 70974 34652
rect 23550 34482 23596 34528
rect 70824 34502 70870 34548
rect 70928 34502 70974 34548
rect 23682 34350 23728 34396
rect 70824 34398 70870 34444
rect 70928 34398 70974 34444
rect 70824 34294 70870 34340
rect 70928 34294 70974 34340
rect 23814 34218 23860 34264
rect 70824 34190 70870 34236
rect 70928 34190 70974 34236
rect 23946 34086 23992 34132
rect 70824 34086 70870 34132
rect 70928 34086 70974 34132
rect 24078 33954 24124 34000
rect 70824 33982 70870 34028
rect 70928 33982 70974 34028
rect 24210 33822 24256 33868
rect 70824 33878 70870 33924
rect 70928 33878 70974 33924
rect 70824 33774 70870 33820
rect 70928 33774 70974 33820
rect 24342 33690 24388 33736
rect 70824 33670 70870 33716
rect 70928 33670 70974 33716
rect 24474 33558 24520 33604
rect 70824 33566 70870 33612
rect 70928 33566 70974 33612
rect 24606 33426 24652 33472
rect 70824 33462 70870 33508
rect 70928 33462 70974 33508
rect 24738 33294 24784 33340
rect 70824 33358 70870 33404
rect 70928 33358 70974 33404
rect 70824 33254 70870 33300
rect 70928 33254 70974 33300
rect 24870 33162 24916 33208
rect 70824 33150 70870 33196
rect 70928 33150 70974 33196
rect 25002 33030 25048 33076
rect 70824 33046 70870 33092
rect 70928 33046 70974 33092
rect 25134 32898 25180 32944
rect 70824 32942 70870 32988
rect 70928 32942 70974 32988
rect 70824 32838 70870 32884
rect 70928 32838 70974 32884
rect 25266 32766 25312 32812
rect 70824 32734 70870 32780
rect 70928 32734 70974 32780
rect 25398 32634 25444 32680
rect 70824 32630 70870 32676
rect 70928 32630 70974 32676
rect 25530 32502 25576 32548
rect 70824 32526 70870 32572
rect 70928 32526 70974 32572
rect 70824 32422 70870 32468
rect 70928 32422 70974 32468
rect 25662 32370 25708 32416
rect 25794 32238 25840 32284
rect 70824 32318 70870 32364
rect 70928 32318 70974 32364
rect 70824 32214 70870 32260
rect 70928 32214 70974 32260
rect 25926 32106 25972 32152
rect 70824 32110 70870 32156
rect 70928 32110 70974 32156
rect 26058 31974 26104 32020
rect 70824 32006 70870 32052
rect 70928 32006 70974 32052
rect 26190 31842 26236 31888
rect 70824 31902 70870 31948
rect 70928 31902 70974 31948
rect 70824 31798 70870 31844
rect 70928 31798 70974 31844
rect 26322 31710 26368 31756
rect 70824 31694 70870 31740
rect 70928 31694 70974 31740
rect 26454 31578 26500 31624
rect 70824 31590 70870 31636
rect 70928 31590 70974 31636
rect 26586 31446 26632 31492
rect 70824 31486 70870 31532
rect 70928 31486 70974 31532
rect 70824 31382 70870 31428
rect 70928 31382 70974 31428
rect 26718 31314 26764 31360
rect 70824 31278 70870 31324
rect 70928 31278 70974 31324
rect 26850 31182 26896 31228
rect 70824 31174 70870 31220
rect 70928 31174 70974 31220
rect 26982 31050 27028 31096
rect 70824 31070 70870 31116
rect 70928 31070 70974 31116
rect 27114 30918 27160 30964
rect 70824 30966 70870 31012
rect 70928 30966 70974 31012
rect 70824 30862 70870 30908
rect 70928 30862 70974 30908
rect 27246 30786 27292 30832
rect 70824 30758 70870 30804
rect 70928 30758 70974 30804
rect 27378 30654 27424 30700
rect 70824 30654 70870 30700
rect 70928 30654 70974 30700
rect 27510 30522 27556 30568
rect 70824 30550 70870 30596
rect 70928 30550 70974 30596
rect 70824 30446 70870 30492
rect 70928 30446 70974 30492
rect 27642 30390 27688 30436
rect 70824 30342 70870 30388
rect 70928 30342 70974 30388
rect 27774 30258 27820 30304
rect 70824 30238 70870 30284
rect 70928 30238 70974 30284
rect 27906 30126 27952 30172
rect 70824 30134 70870 30180
rect 70928 30134 70974 30180
rect 28038 29994 28084 30040
rect 70824 30030 70870 30076
rect 70928 30030 70974 30076
rect 28170 29862 28216 29908
rect 70824 29926 70870 29972
rect 70928 29926 70974 29972
rect 70824 29822 70870 29868
rect 70928 29822 70974 29868
rect 28302 29730 28348 29776
rect 70824 29718 70870 29764
rect 70928 29718 70974 29764
rect 28434 29598 28480 29644
rect 70824 29614 70870 29660
rect 70928 29614 70974 29660
rect 28566 29466 28612 29512
rect 70824 29510 70870 29556
rect 70928 29510 70974 29556
rect 70824 29406 70870 29452
rect 70928 29406 70974 29452
rect 28698 29334 28744 29380
rect 70824 29302 70870 29348
rect 70928 29302 70974 29348
rect 28830 29202 28876 29248
rect 70824 29198 70870 29244
rect 70928 29198 70974 29244
rect 28962 29070 29008 29116
rect 70824 29094 70870 29140
rect 70928 29094 70974 29140
rect 29094 28938 29140 28984
rect 70824 28990 70870 29036
rect 70928 28990 70974 29036
rect 70824 28886 70870 28932
rect 70928 28886 70974 28932
rect 29226 28806 29272 28852
rect 70824 28782 70870 28828
rect 70928 28782 70974 28828
rect 29358 28674 29404 28720
rect 70824 28678 70870 28724
rect 70928 28678 70974 28724
rect 29490 28542 29536 28588
rect 70824 28574 70870 28620
rect 70928 28574 70974 28620
rect 29622 28410 29668 28456
rect 70824 28470 70870 28516
rect 70928 28470 70974 28516
rect 70824 28366 70870 28412
rect 70928 28366 70974 28412
rect 29754 28278 29800 28324
rect 70824 28262 70870 28308
rect 70928 28262 70974 28308
rect 29886 28146 29932 28192
rect 70824 28158 70870 28204
rect 70928 28158 70974 28204
rect 30018 28014 30064 28060
rect 70824 28054 70870 28100
rect 70928 28054 70974 28100
rect 30150 27882 30196 27928
rect 70824 27950 70870 27996
rect 70928 27950 70974 27996
rect 70824 27846 70870 27892
rect 70928 27846 70974 27892
rect 30282 27750 30328 27796
rect 70824 27742 70870 27788
rect 70928 27742 70974 27788
rect 30414 27618 30460 27664
rect 70824 27638 70870 27684
rect 70928 27638 70974 27684
rect 30546 27486 30592 27532
rect 70824 27534 70870 27580
rect 70928 27534 70974 27580
rect 70824 27430 70870 27476
rect 70928 27430 70974 27476
rect 30678 27354 30724 27400
rect 70824 27326 70870 27372
rect 70928 27326 70974 27372
rect 30810 27222 30856 27268
rect 70824 27222 70870 27268
rect 70928 27222 70974 27268
rect 30942 27090 30988 27136
rect 70824 27118 70870 27164
rect 70928 27118 70974 27164
rect 31074 26958 31120 27004
rect 70824 27014 70870 27060
rect 70928 27014 70974 27060
rect 70824 26910 70870 26956
rect 70928 26910 70974 26956
rect 31206 26826 31252 26872
rect 70824 26806 70870 26852
rect 70928 26806 70974 26852
rect 31338 26694 31384 26740
rect 70824 26702 70870 26748
rect 70928 26702 70974 26748
rect 31470 26562 31516 26608
rect 70824 26598 70870 26644
rect 70928 26598 70974 26644
rect 31602 26430 31648 26476
rect 70824 26494 70870 26540
rect 70928 26494 70974 26540
rect 70824 26390 70870 26436
rect 70928 26390 70974 26436
rect 31734 26298 31780 26344
rect 70824 26286 70870 26332
rect 70928 26286 70974 26332
rect 31866 26166 31912 26212
rect 70824 26182 70870 26228
rect 70928 26182 70974 26228
rect 31998 26034 32044 26080
rect 70824 26078 70870 26124
rect 70928 26078 70974 26124
rect 70824 25974 70870 26020
rect 70928 25974 70974 26020
rect 32130 25902 32176 25948
rect 70824 25870 70870 25916
rect 70928 25870 70974 25916
rect 32262 25770 32308 25816
rect 70824 25766 70870 25812
rect 70928 25766 70974 25812
rect 32394 25638 32440 25684
rect 70824 25662 70870 25708
rect 70928 25662 70974 25708
rect 32526 25506 32572 25552
rect 70824 25558 70870 25604
rect 70928 25558 70974 25604
rect 32658 25374 32704 25420
rect 70824 25454 70870 25500
rect 70928 25454 70974 25500
rect 70824 25350 70870 25396
rect 70928 25350 70974 25396
rect 32790 25242 32836 25288
rect 70824 25246 70870 25292
rect 70928 25246 70974 25292
rect 32922 25110 32968 25156
rect 70824 25142 70870 25188
rect 70928 25142 70974 25188
rect 33054 24978 33100 25024
rect 70824 25038 70870 25084
rect 70928 25038 70974 25084
rect 70824 24934 70870 24980
rect 70928 24934 70974 24980
rect 33186 24846 33232 24892
rect 70824 24830 70870 24876
rect 70928 24830 70974 24876
rect 33318 24714 33364 24760
rect 70824 24726 70870 24772
rect 70928 24726 70974 24772
rect 33450 24582 33496 24628
rect 70824 24622 70870 24668
rect 70928 24622 70974 24668
rect 70824 24518 70870 24564
rect 70928 24518 70974 24564
rect 33582 24450 33628 24496
rect 70824 24414 70870 24460
rect 70928 24414 70974 24460
rect 33714 24318 33760 24364
rect 70824 24310 70870 24356
rect 70928 24310 70974 24356
rect 33846 24186 33892 24232
rect 70824 24206 70870 24252
rect 70928 24206 70974 24252
rect 33978 24054 34024 24100
rect 70824 24102 70870 24148
rect 70928 24102 70974 24148
rect 34110 23922 34156 23968
rect 70824 23998 70870 24044
rect 70928 23998 70974 24044
rect 70824 23894 70870 23940
rect 70928 23894 70974 23940
rect 34242 23790 34288 23836
rect 70824 23790 70870 23836
rect 70928 23790 70974 23836
rect 34374 23658 34420 23704
rect 70824 23686 70870 23732
rect 70928 23686 70974 23732
rect 34506 23526 34552 23572
rect 70824 23582 70870 23628
rect 70928 23582 70974 23628
rect 70824 23478 70870 23524
rect 70928 23478 70974 23524
rect 34638 23394 34684 23440
rect 70824 23374 70870 23420
rect 70928 23374 70974 23420
rect 34770 23262 34816 23308
rect 70824 23270 70870 23316
rect 70928 23270 70974 23316
rect 34902 23130 34948 23176
rect 70824 23166 70870 23212
rect 70928 23166 70974 23212
rect 35034 22998 35080 23044
rect 70824 23062 70870 23108
rect 70928 23062 70974 23108
rect 70824 22958 70870 23004
rect 70928 22958 70974 23004
rect 35166 22866 35212 22912
rect 70824 22854 70870 22900
rect 70928 22854 70974 22900
rect 35298 22734 35344 22780
rect 70824 22750 70870 22796
rect 70928 22750 70974 22796
rect 35430 22602 35476 22648
rect 70824 22646 70870 22692
rect 70928 22646 70974 22692
rect 70824 22542 70870 22588
rect 70928 22542 70974 22588
rect 35562 22470 35608 22516
rect 70824 22438 70870 22484
rect 70928 22438 70974 22484
rect 35694 22338 35740 22384
rect 70824 22334 70870 22380
rect 70928 22334 70974 22380
rect 35826 22206 35872 22252
rect 70824 22230 70870 22276
rect 70928 22230 70974 22276
rect 70824 22126 70870 22172
rect 70928 22126 70974 22172
rect 35958 22074 36004 22120
rect 70824 22022 70870 22068
rect 70928 22022 70974 22068
rect 36090 21942 36136 21988
rect 70824 21918 70870 21964
rect 70928 21918 70974 21964
rect 36222 21810 36268 21856
rect 70824 21814 70870 21860
rect 70928 21814 70974 21860
rect 36354 21678 36400 21724
rect 70824 21710 70870 21756
rect 70928 21710 70974 21756
rect 36486 21546 36532 21592
rect 70824 21606 70870 21652
rect 70928 21606 70974 21652
rect 70824 21502 70870 21548
rect 70928 21502 70974 21548
rect 36618 21414 36664 21460
rect 70824 21398 70870 21444
rect 70928 21398 70974 21444
rect 36750 21282 36796 21328
rect 70824 21294 70870 21340
rect 70928 21294 70974 21340
rect 36882 21150 36928 21196
rect 70824 21190 70870 21236
rect 70928 21190 70974 21236
rect 70824 21086 70870 21132
rect 70928 21086 70974 21132
rect 37014 21018 37060 21064
rect 70824 20982 70870 21028
rect 70928 20982 70974 21028
rect 37146 20886 37192 20932
rect 70824 20878 70870 20924
rect 70928 20878 70974 20924
rect 37278 20754 37324 20800
rect 70824 20774 70870 20820
rect 70928 20774 70974 20820
rect 37410 20622 37456 20668
rect 70824 20670 70870 20716
rect 70928 20670 70974 20716
rect 70824 20566 70870 20612
rect 70928 20566 70974 20612
rect 37542 20490 37588 20536
rect 70824 20462 70870 20508
rect 70928 20462 70974 20508
rect 37674 20358 37720 20404
rect 70824 20358 70870 20404
rect 70928 20358 70974 20404
rect 37806 20226 37852 20272
rect 70824 20254 70870 20300
rect 70928 20254 70974 20300
rect 37938 20094 37984 20140
rect 70824 20150 70870 20196
rect 70928 20150 70974 20196
rect 70824 20046 70870 20092
rect 70928 20046 70974 20092
rect 38070 19962 38116 20008
rect 70824 19942 70870 19988
rect 70928 19942 70974 19988
rect 38202 19830 38248 19876
rect 70824 19838 70870 19884
rect 70928 19838 70974 19884
rect 38334 19698 38380 19744
rect 70824 19734 70870 19780
rect 70928 19734 70974 19780
rect 38466 19566 38512 19612
rect 70824 19630 70870 19676
rect 70928 19630 70974 19676
rect 70824 19526 70870 19572
rect 70928 19526 70974 19572
rect 38598 19434 38644 19480
rect 70824 19422 70870 19468
rect 70928 19422 70974 19468
rect 38730 19302 38776 19348
rect 70824 19318 70870 19364
rect 70928 19318 70974 19364
rect 38862 19170 38908 19216
rect 70824 19214 70870 19260
rect 70928 19214 70974 19260
rect 38994 19038 39040 19084
rect 70824 19110 70870 19156
rect 70928 19110 70974 19156
rect 70824 19006 70870 19052
rect 70928 19006 70974 19052
rect 39126 18906 39172 18952
rect 70824 18902 70870 18948
rect 70928 18902 70974 18948
rect 39258 18774 39304 18820
rect 70824 18798 70870 18844
rect 70928 18798 70974 18844
rect 39390 18642 39436 18688
rect 70824 18694 70870 18740
rect 70928 18694 70974 18740
rect 39522 18510 39568 18556
rect 70824 18590 70870 18636
rect 70928 18590 70974 18636
rect 70824 18486 70870 18532
rect 70928 18486 70974 18532
rect 39654 18378 39700 18424
rect 70824 18382 70870 18428
rect 70928 18382 70974 18428
rect 39786 18246 39832 18292
rect 70824 18278 70870 18324
rect 70928 18278 70974 18324
rect 39918 18114 39964 18160
rect 70824 18174 70870 18220
rect 70928 18174 70974 18220
rect 70824 18070 70870 18116
rect 70928 18070 70974 18116
rect 40050 17982 40096 18028
rect 70824 17966 70870 18012
rect 70928 17966 70974 18012
rect 40182 17850 40228 17896
rect 70824 17862 70870 17908
rect 70928 17862 70974 17908
rect 40314 17718 40360 17764
rect 70824 17758 70870 17804
rect 70928 17758 70974 17804
rect 70824 17654 70870 17700
rect 70928 17654 70974 17700
rect 40446 17586 40492 17632
rect 70824 17550 70870 17596
rect 70928 17550 70974 17596
rect 40578 17454 40624 17500
rect 70824 17446 70870 17492
rect 70928 17446 70974 17492
rect 40710 17322 40756 17368
rect 70824 17342 70870 17388
rect 70928 17342 70974 17388
rect 70824 17238 70870 17284
rect 70928 17238 70974 17284
rect 40842 17190 40888 17236
rect 40974 17058 41020 17104
rect 70824 17134 70870 17180
rect 70928 17134 70974 17180
rect 70824 17030 70870 17076
rect 70928 17030 70974 17076
rect 41106 16926 41152 16972
rect 70824 16926 70870 16972
rect 70928 16926 70974 16972
rect 41238 16794 41284 16840
rect 70824 16822 70870 16868
rect 70928 16822 70974 16868
rect 41370 16662 41416 16708
rect 70824 16718 70870 16764
rect 70928 16718 70974 16764
rect 70824 16614 70870 16660
rect 70928 16614 70974 16660
rect 41502 16530 41548 16576
rect 70824 16510 70870 16556
rect 70928 16510 70974 16556
rect 41634 16398 41680 16444
rect 70824 16406 70870 16452
rect 70928 16406 70974 16452
rect 41766 16266 41812 16312
rect 70824 16302 70870 16348
rect 70928 16302 70974 16348
rect 41898 16134 41944 16180
rect 70824 16198 70870 16244
rect 70928 16198 70974 16244
rect 70824 16094 70870 16140
rect 70928 16094 70974 16140
rect 42030 16002 42076 16048
rect 70824 15990 70870 16036
rect 70928 15990 70974 16036
rect 42162 15870 42208 15916
rect 70824 15886 70870 15932
rect 70928 15886 70974 15932
rect 42294 15738 42340 15784
rect 70824 15782 70870 15828
rect 70928 15782 70974 15828
rect 70824 15678 70870 15724
rect 70928 15678 70974 15724
rect 42426 15606 42472 15652
rect 70824 15574 70870 15620
rect 70928 15574 70974 15620
rect 42558 15474 42604 15520
rect 70824 15470 70870 15516
rect 70928 15470 70974 15516
rect 42690 15342 42736 15388
rect 70824 15366 70870 15412
rect 70928 15366 70974 15412
rect 70824 15262 70870 15308
rect 70928 15262 70974 15308
rect 42822 15210 42868 15256
rect 70824 15158 70870 15204
rect 70928 15158 70974 15204
rect 42954 15078 43000 15124
rect 70824 15054 70870 15100
rect 70928 15054 70974 15100
rect 43086 14946 43132 14992
rect 70824 14950 70870 14996
rect 70928 14950 70974 14996
rect 43218 14814 43264 14860
rect 70824 14846 70870 14892
rect 70928 14846 70974 14892
rect 43350 14682 43396 14728
rect 70824 14742 70870 14788
rect 70928 14742 70974 14788
rect 70824 14638 70870 14684
rect 70928 14638 70974 14684
rect 43482 14550 43528 14596
rect 70824 14534 70870 14580
rect 70928 14534 70974 14580
rect 43614 14418 43660 14464
rect 70824 14430 70870 14476
rect 70928 14430 70974 14476
rect 43746 14286 43792 14332
rect 70824 14326 70870 14372
rect 70928 14326 70974 14372
rect 70824 14222 70870 14268
rect 70928 14222 70974 14268
rect 43878 14154 43924 14200
rect 70824 14118 70870 14164
rect 70928 14118 70974 14164
rect 44010 14022 44056 14068
rect 70824 14014 70870 14060
rect 70928 14014 70974 14060
rect 44142 13890 44188 13936
rect 70824 13910 70870 13956
rect 70928 13910 70974 13956
rect 44274 13758 44320 13804
rect 70824 13806 70870 13852
rect 70928 13806 70974 13852
rect 70824 13702 70870 13748
rect 70928 13702 70974 13748
rect 44406 13626 44452 13672
rect 70824 13598 70870 13644
rect 70928 13598 70974 13644
rect 44538 13494 44584 13540
rect 70824 13494 70870 13540
rect 70928 13494 70974 13540
rect 44670 13362 44716 13408
rect 70824 13390 70870 13436
rect 70928 13390 70974 13436
rect 44850 13210 44896 13256
rect 45088 13223 45134 13269
rect 45192 13223 45238 13269
rect 45296 13223 45342 13269
rect 45400 13223 45446 13269
rect 45504 13223 45550 13269
rect 45608 13223 45654 13269
rect 45712 13223 45758 13269
rect 45816 13223 45862 13269
rect 45920 13223 45966 13269
rect 46024 13223 46070 13269
rect 46128 13223 46174 13269
rect 46232 13223 46278 13269
rect 46336 13223 46382 13269
rect 46440 13223 46486 13269
rect 46544 13223 46590 13269
rect 46648 13223 46694 13269
rect 46752 13223 46798 13269
rect 46856 13223 46902 13269
rect 46960 13223 47006 13269
rect 47064 13223 47110 13269
rect 47168 13223 47214 13269
rect 47272 13223 47318 13269
rect 47376 13223 47422 13269
rect 47480 13223 47526 13269
rect 47584 13223 47630 13269
rect 47688 13223 47734 13269
rect 47792 13223 47838 13269
rect 47896 13223 47942 13269
rect 48000 13223 48046 13269
rect 48104 13223 48150 13269
rect 48208 13223 48254 13269
rect 48312 13223 48358 13269
rect 48416 13223 48462 13269
rect 48520 13223 48566 13269
rect 48624 13223 48670 13269
rect 48728 13223 48774 13269
rect 48832 13223 48878 13269
rect 48936 13223 48982 13269
rect 49040 13223 49086 13269
rect 49144 13223 49190 13269
rect 49248 13223 49294 13269
rect 49352 13223 49398 13269
rect 49456 13223 49502 13269
rect 49560 13223 49606 13269
rect 49664 13223 49710 13269
rect 49768 13223 49814 13269
rect 49872 13223 49918 13269
rect 49976 13223 50022 13269
rect 50080 13223 50126 13269
rect 50184 13223 50230 13269
rect 50288 13223 50334 13269
rect 50392 13223 50438 13269
rect 50496 13223 50542 13269
rect 50600 13223 50646 13269
rect 50704 13223 50750 13269
rect 50808 13223 50854 13269
rect 50912 13223 50958 13269
rect 51016 13223 51062 13269
rect 51120 13223 51166 13269
rect 51224 13223 51270 13269
rect 51328 13223 51374 13269
rect 51432 13223 51478 13269
rect 51536 13223 51582 13269
rect 51640 13223 51686 13269
rect 51744 13223 51790 13269
rect 51848 13223 51894 13269
rect 51952 13223 51998 13269
rect 52056 13223 52102 13269
rect 52160 13223 52206 13269
rect 52264 13223 52310 13269
rect 52368 13223 52414 13269
rect 52472 13223 52518 13269
rect 52576 13223 52622 13269
rect 52680 13223 52726 13269
rect 52784 13223 52830 13269
rect 52888 13223 52934 13269
rect 52992 13223 53038 13269
rect 53096 13223 53142 13269
rect 53200 13223 53246 13269
rect 53304 13223 53350 13269
rect 53408 13223 53454 13269
rect 53512 13223 53558 13269
rect 53616 13223 53662 13269
rect 53720 13223 53766 13269
rect 53824 13223 53870 13269
rect 53928 13223 53974 13269
rect 54032 13223 54078 13269
rect 54136 13223 54182 13269
rect 54240 13223 54286 13269
rect 54344 13223 54390 13269
rect 54448 13223 54494 13269
rect 54552 13223 54598 13269
rect 54656 13223 54702 13269
rect 54760 13223 54806 13269
rect 54864 13223 54910 13269
rect 54968 13223 55014 13269
rect 55072 13223 55118 13269
rect 55176 13223 55222 13269
rect 55280 13223 55326 13269
rect 55384 13223 55430 13269
rect 55488 13223 55534 13269
rect 55592 13223 55638 13269
rect 55696 13223 55742 13269
rect 55800 13223 55846 13269
rect 55904 13223 55950 13269
rect 56008 13223 56054 13269
rect 56112 13223 56158 13269
rect 56216 13223 56262 13269
rect 56320 13223 56366 13269
rect 56424 13223 56470 13269
rect 56528 13223 56574 13269
rect 56632 13223 56678 13269
rect 56736 13223 56782 13269
rect 56840 13223 56886 13269
rect 56944 13223 56990 13269
rect 57048 13223 57094 13269
rect 57152 13223 57198 13269
rect 57256 13223 57302 13269
rect 57360 13223 57406 13269
rect 57464 13223 57510 13269
rect 57568 13223 57614 13269
rect 57672 13223 57718 13269
rect 57776 13223 57822 13269
rect 57880 13223 57926 13269
rect 57984 13223 58030 13269
rect 58088 13223 58134 13269
rect 58192 13223 58238 13269
rect 58296 13223 58342 13269
rect 58400 13223 58446 13269
rect 58504 13223 58550 13269
rect 58608 13223 58654 13269
rect 58712 13223 58758 13269
rect 58816 13223 58862 13269
rect 58920 13223 58966 13269
rect 59024 13223 59070 13269
rect 59128 13223 59174 13269
rect 59232 13223 59278 13269
rect 59336 13223 59382 13269
rect 59440 13223 59486 13269
rect 59544 13223 59590 13269
rect 59648 13223 59694 13269
rect 59752 13223 59798 13269
rect 59856 13223 59902 13269
rect 59960 13223 60006 13269
rect 60064 13223 60110 13269
rect 60168 13223 60214 13269
rect 60272 13223 60318 13269
rect 60376 13223 60422 13269
rect 60480 13223 60526 13269
rect 60584 13223 60630 13269
rect 60688 13223 60734 13269
rect 60792 13223 60838 13269
rect 60896 13223 60942 13269
rect 61000 13223 61046 13269
rect 61104 13223 61150 13269
rect 61208 13223 61254 13269
rect 61312 13223 61358 13269
rect 61416 13223 61462 13269
rect 61520 13223 61566 13269
rect 61624 13223 61670 13269
rect 61728 13223 61774 13269
rect 61832 13223 61878 13269
rect 61936 13223 61982 13269
rect 62040 13223 62086 13269
rect 62144 13223 62190 13269
rect 62248 13223 62294 13269
rect 62352 13223 62398 13269
rect 62456 13223 62502 13269
rect 62560 13223 62606 13269
rect 62664 13223 62710 13269
rect 62768 13223 62814 13269
rect 62872 13223 62918 13269
rect 62976 13223 63022 13269
rect 63080 13223 63126 13269
rect 63184 13223 63230 13269
rect 63288 13223 63334 13269
rect 63392 13223 63438 13269
rect 63496 13223 63542 13269
rect 63600 13223 63646 13269
rect 63704 13223 63750 13269
rect 63808 13223 63854 13269
rect 63912 13223 63958 13269
rect 64016 13223 64062 13269
rect 64120 13223 64166 13269
rect 64224 13223 64270 13269
rect 64328 13223 64374 13269
rect 64432 13223 64478 13269
rect 64536 13223 64582 13269
rect 64640 13223 64686 13269
rect 64744 13223 64790 13269
rect 64848 13223 64894 13269
rect 64952 13223 64998 13269
rect 65056 13223 65102 13269
rect 65160 13223 65206 13269
rect 65264 13223 65310 13269
rect 65368 13223 65414 13269
rect 65472 13223 65518 13269
rect 65576 13223 65622 13269
rect 65680 13223 65726 13269
rect 65784 13223 65830 13269
rect 65888 13223 65934 13269
rect 65992 13223 66038 13269
rect 66096 13223 66142 13269
rect 66200 13223 66246 13269
rect 66304 13223 66350 13269
rect 66408 13223 66454 13269
rect 66512 13223 66558 13269
rect 66616 13223 66662 13269
rect 66720 13223 66766 13269
rect 66824 13223 66870 13269
rect 66928 13223 66974 13269
rect 67032 13223 67078 13269
rect 67136 13223 67182 13269
rect 67240 13223 67286 13269
rect 67344 13223 67390 13269
rect 67448 13223 67494 13269
rect 67552 13223 67598 13269
rect 67656 13223 67702 13269
rect 67760 13223 67806 13269
rect 67864 13223 67910 13269
rect 67968 13223 68014 13269
rect 68072 13223 68118 13269
rect 68176 13223 68222 13269
rect 68280 13223 68326 13269
rect 68384 13223 68430 13269
rect 68488 13223 68534 13269
rect 68592 13223 68638 13269
rect 68696 13223 68742 13269
rect 68800 13223 68846 13269
rect 68904 13223 68950 13269
rect 69008 13223 69054 13269
rect 69112 13223 69158 13269
rect 69216 13223 69262 13269
rect 69320 13223 69366 13269
rect 69424 13223 69470 13269
rect 69528 13223 69574 13269
rect 69632 13223 69678 13269
rect 69736 13223 69782 13269
rect 69840 13223 69886 13269
rect 69944 13223 69990 13269
rect 70048 13223 70094 13269
rect 70152 13223 70198 13269
rect 70256 13223 70302 13269
rect 70360 13223 70406 13269
rect 70464 13223 70510 13269
rect 70568 13223 70614 13269
rect 70672 13223 70718 13269
rect 70776 13223 70822 13269
rect 70880 13223 70926 13269
rect 45088 13119 45134 13165
rect 45192 13119 45238 13165
rect 45296 13119 45342 13165
rect 45400 13119 45446 13165
rect 45504 13119 45550 13165
rect 45608 13119 45654 13165
rect 45712 13119 45758 13165
rect 45816 13119 45862 13165
rect 45920 13119 45966 13165
rect 46024 13119 46070 13165
rect 46128 13119 46174 13165
rect 46232 13119 46278 13165
rect 46336 13119 46382 13165
rect 46440 13119 46486 13165
rect 46544 13119 46590 13165
rect 46648 13119 46694 13165
rect 46752 13119 46798 13165
rect 46856 13119 46902 13165
rect 46960 13119 47006 13165
rect 47064 13119 47110 13165
rect 47168 13119 47214 13165
rect 47272 13119 47318 13165
rect 47376 13119 47422 13165
rect 47480 13119 47526 13165
rect 47584 13119 47630 13165
rect 47688 13119 47734 13165
rect 47792 13119 47838 13165
rect 47896 13119 47942 13165
rect 48000 13119 48046 13165
rect 48104 13119 48150 13165
rect 48208 13119 48254 13165
rect 48312 13119 48358 13165
rect 48416 13119 48462 13165
rect 48520 13119 48566 13165
rect 48624 13119 48670 13165
rect 48728 13119 48774 13165
rect 48832 13119 48878 13165
rect 48936 13119 48982 13165
rect 49040 13119 49086 13165
rect 49144 13119 49190 13165
rect 49248 13119 49294 13165
rect 49352 13119 49398 13165
rect 49456 13119 49502 13165
rect 49560 13119 49606 13165
rect 49664 13119 49710 13165
rect 49768 13119 49814 13165
rect 49872 13119 49918 13165
rect 49976 13119 50022 13165
rect 50080 13119 50126 13165
rect 50184 13119 50230 13165
rect 50288 13119 50334 13165
rect 50392 13119 50438 13165
rect 50496 13119 50542 13165
rect 50600 13119 50646 13165
rect 50704 13119 50750 13165
rect 50808 13119 50854 13165
rect 50912 13119 50958 13165
rect 51016 13119 51062 13165
rect 51120 13119 51166 13165
rect 51224 13119 51270 13165
rect 51328 13119 51374 13165
rect 51432 13119 51478 13165
rect 51536 13119 51582 13165
rect 51640 13119 51686 13165
rect 51744 13119 51790 13165
rect 51848 13119 51894 13165
rect 51952 13119 51998 13165
rect 52056 13119 52102 13165
rect 52160 13119 52206 13165
rect 52264 13119 52310 13165
rect 52368 13119 52414 13165
rect 52472 13119 52518 13165
rect 52576 13119 52622 13165
rect 52680 13119 52726 13165
rect 52784 13119 52830 13165
rect 52888 13119 52934 13165
rect 52992 13119 53038 13165
rect 53096 13119 53142 13165
rect 53200 13119 53246 13165
rect 53304 13119 53350 13165
rect 53408 13119 53454 13165
rect 53512 13119 53558 13165
rect 53616 13119 53662 13165
rect 53720 13119 53766 13165
rect 53824 13119 53870 13165
rect 53928 13119 53974 13165
rect 54032 13119 54078 13165
rect 54136 13119 54182 13165
rect 54240 13119 54286 13165
rect 54344 13119 54390 13165
rect 54448 13119 54494 13165
rect 54552 13119 54598 13165
rect 54656 13119 54702 13165
rect 54760 13119 54806 13165
rect 54864 13119 54910 13165
rect 54968 13119 55014 13165
rect 55072 13119 55118 13165
rect 55176 13119 55222 13165
rect 55280 13119 55326 13165
rect 55384 13119 55430 13165
rect 55488 13119 55534 13165
rect 55592 13119 55638 13165
rect 55696 13119 55742 13165
rect 55800 13119 55846 13165
rect 55904 13119 55950 13165
rect 56008 13119 56054 13165
rect 56112 13119 56158 13165
rect 56216 13119 56262 13165
rect 56320 13119 56366 13165
rect 56424 13119 56470 13165
rect 56528 13119 56574 13165
rect 56632 13119 56678 13165
rect 56736 13119 56782 13165
rect 56840 13119 56886 13165
rect 56944 13119 56990 13165
rect 57048 13119 57094 13165
rect 57152 13119 57198 13165
rect 57256 13119 57302 13165
rect 57360 13119 57406 13165
rect 57464 13119 57510 13165
rect 57568 13119 57614 13165
rect 57672 13119 57718 13165
rect 57776 13119 57822 13165
rect 57880 13119 57926 13165
rect 57984 13119 58030 13165
rect 58088 13119 58134 13165
rect 58192 13119 58238 13165
rect 58296 13119 58342 13165
rect 58400 13119 58446 13165
rect 58504 13119 58550 13165
rect 58608 13119 58654 13165
rect 58712 13119 58758 13165
rect 58816 13119 58862 13165
rect 58920 13119 58966 13165
rect 59024 13119 59070 13165
rect 59128 13119 59174 13165
rect 59232 13119 59278 13165
rect 59336 13119 59382 13165
rect 59440 13119 59486 13165
rect 59544 13119 59590 13165
rect 59648 13119 59694 13165
rect 59752 13119 59798 13165
rect 59856 13119 59902 13165
rect 59960 13119 60006 13165
rect 60064 13119 60110 13165
rect 60168 13119 60214 13165
rect 60272 13119 60318 13165
rect 60376 13119 60422 13165
rect 60480 13119 60526 13165
rect 60584 13119 60630 13165
rect 60688 13119 60734 13165
rect 60792 13119 60838 13165
rect 60896 13119 60942 13165
rect 61000 13119 61046 13165
rect 61104 13119 61150 13165
rect 61208 13119 61254 13165
rect 61312 13119 61358 13165
rect 61416 13119 61462 13165
rect 61520 13119 61566 13165
rect 61624 13119 61670 13165
rect 61728 13119 61774 13165
rect 61832 13119 61878 13165
rect 61936 13119 61982 13165
rect 62040 13119 62086 13165
rect 62144 13119 62190 13165
rect 62248 13119 62294 13165
rect 62352 13119 62398 13165
rect 62456 13119 62502 13165
rect 62560 13119 62606 13165
rect 62664 13119 62710 13165
rect 62768 13119 62814 13165
rect 62872 13119 62918 13165
rect 62976 13119 63022 13165
rect 63080 13119 63126 13165
rect 63184 13119 63230 13165
rect 63288 13119 63334 13165
rect 63392 13119 63438 13165
rect 63496 13119 63542 13165
rect 63600 13119 63646 13165
rect 63704 13119 63750 13165
rect 63808 13119 63854 13165
rect 63912 13119 63958 13165
rect 64016 13119 64062 13165
rect 64120 13119 64166 13165
rect 64224 13119 64270 13165
rect 64328 13119 64374 13165
rect 64432 13119 64478 13165
rect 64536 13119 64582 13165
rect 64640 13119 64686 13165
rect 64744 13119 64790 13165
rect 64848 13119 64894 13165
rect 64952 13119 64998 13165
rect 65056 13119 65102 13165
rect 65160 13119 65206 13165
rect 65264 13119 65310 13165
rect 65368 13119 65414 13165
rect 65472 13119 65518 13165
rect 65576 13119 65622 13165
rect 65680 13119 65726 13165
rect 65784 13119 65830 13165
rect 65888 13119 65934 13165
rect 65992 13119 66038 13165
rect 66096 13119 66142 13165
rect 66200 13119 66246 13165
rect 66304 13119 66350 13165
rect 66408 13119 66454 13165
rect 66512 13119 66558 13165
rect 66616 13119 66662 13165
rect 66720 13119 66766 13165
rect 66824 13119 66870 13165
rect 66928 13119 66974 13165
rect 67032 13119 67078 13165
rect 67136 13119 67182 13165
rect 67240 13119 67286 13165
rect 67344 13119 67390 13165
rect 67448 13119 67494 13165
rect 67552 13119 67598 13165
rect 67656 13119 67702 13165
rect 67760 13119 67806 13165
rect 67864 13119 67910 13165
rect 67968 13119 68014 13165
rect 68072 13119 68118 13165
rect 68176 13119 68222 13165
rect 68280 13119 68326 13165
rect 68384 13119 68430 13165
rect 68488 13119 68534 13165
rect 68592 13119 68638 13165
rect 68696 13119 68742 13165
rect 68800 13119 68846 13165
rect 68904 13119 68950 13165
rect 69008 13119 69054 13165
rect 69112 13119 69158 13165
rect 69216 13119 69262 13165
rect 69320 13119 69366 13165
rect 69424 13119 69470 13165
rect 69528 13119 69574 13165
rect 69632 13119 69678 13165
rect 69736 13119 69782 13165
rect 69840 13119 69886 13165
rect 69944 13119 69990 13165
rect 70048 13119 70094 13165
rect 70152 13119 70198 13165
rect 70256 13119 70302 13165
rect 70360 13119 70406 13165
rect 70464 13119 70510 13165
rect 70568 13119 70614 13165
rect 70672 13119 70718 13165
rect 70776 13119 70822 13165
rect 70880 13119 70926 13165
<< metal1 >>
rect 13108 70975 69957 71000
rect 13108 70929 13119 70975
rect 13165 70929 13223 70975
rect 13269 70929 13377 70975
rect 13423 70929 13481 70975
rect 13527 70929 13585 70975
rect 13631 70929 13689 70975
rect 13735 70929 13793 70975
rect 13839 70929 13897 70975
rect 13943 70929 14001 70975
rect 14047 70929 14105 70975
rect 14151 70929 14209 70975
rect 14255 70929 14313 70975
rect 14359 70929 14417 70975
rect 14463 70929 14521 70975
rect 14567 70929 14625 70975
rect 14671 70929 14729 70975
rect 14775 70929 14833 70975
rect 14879 70929 14937 70975
rect 14983 70929 15041 70975
rect 15087 70929 15145 70975
rect 15191 70929 15249 70975
rect 15295 70929 15353 70975
rect 15399 70929 15457 70975
rect 15503 70929 15561 70975
rect 15607 70929 15665 70975
rect 15711 70929 15769 70975
rect 15815 70929 15873 70975
rect 15919 70929 15977 70975
rect 16023 70929 16081 70975
rect 16127 70929 16185 70975
rect 16231 70929 16289 70975
rect 16335 70929 16393 70975
rect 16439 70929 16497 70975
rect 16543 70929 16601 70975
rect 16647 70929 16705 70975
rect 16751 70929 16809 70975
rect 16855 70929 16913 70975
rect 16959 70929 17017 70975
rect 17063 70929 17121 70975
rect 17167 70929 17225 70975
rect 17271 70929 17329 70975
rect 17375 70929 17433 70975
rect 17479 70929 17537 70975
rect 17583 70929 17641 70975
rect 17687 70929 17745 70975
rect 17791 70929 17849 70975
rect 17895 70929 17953 70975
rect 17999 70929 18057 70975
rect 18103 70929 18161 70975
rect 18207 70929 18265 70975
rect 18311 70929 18369 70975
rect 18415 70929 18473 70975
rect 18519 70929 18577 70975
rect 18623 70929 18681 70975
rect 18727 70929 18785 70975
rect 18831 70929 18889 70975
rect 18935 70929 18993 70975
rect 19039 70929 19097 70975
rect 19143 70929 19201 70975
rect 19247 70929 19305 70975
rect 19351 70929 19409 70975
rect 19455 70929 19513 70975
rect 19559 70929 19617 70975
rect 19663 70929 19721 70975
rect 19767 70929 19825 70975
rect 19871 70929 19929 70975
rect 19975 70929 20033 70975
rect 20079 70929 20137 70975
rect 20183 70929 20241 70975
rect 20287 70929 20345 70975
rect 20391 70929 20449 70975
rect 20495 70929 20553 70975
rect 20599 70929 20657 70975
rect 20703 70929 20761 70975
rect 20807 70929 20865 70975
rect 20911 70929 20969 70975
rect 21015 70929 21073 70975
rect 21119 70929 21177 70975
rect 21223 70929 21281 70975
rect 21327 70929 21385 70975
rect 21431 70929 21489 70975
rect 21535 70929 21593 70975
rect 21639 70929 21697 70975
rect 21743 70929 21801 70975
rect 21847 70929 21905 70975
rect 21951 70929 22009 70975
rect 22055 70929 22113 70975
rect 22159 70929 22217 70975
rect 22263 70929 22321 70975
rect 22367 70929 22425 70975
rect 22471 70929 22529 70975
rect 22575 70929 22633 70975
rect 22679 70929 22737 70975
rect 22783 70929 22841 70975
rect 22887 70929 22945 70975
rect 22991 70929 23049 70975
rect 23095 70929 23153 70975
rect 23199 70929 23257 70975
rect 23303 70929 23361 70975
rect 23407 70929 23465 70975
rect 23511 70929 23569 70975
rect 23615 70929 23673 70975
rect 23719 70929 23777 70975
rect 23823 70929 23881 70975
rect 23927 70929 23985 70975
rect 24031 70929 24089 70975
rect 24135 70929 24193 70975
rect 24239 70929 24297 70975
rect 24343 70929 24401 70975
rect 24447 70929 24505 70975
rect 24551 70929 24609 70975
rect 24655 70929 24713 70975
rect 24759 70929 24817 70975
rect 24863 70929 24921 70975
rect 24967 70929 25025 70975
rect 25071 70929 25129 70975
rect 25175 70929 25233 70975
rect 25279 70929 25337 70975
rect 25383 70929 25441 70975
rect 25487 70929 25545 70975
rect 25591 70929 25649 70975
rect 25695 70929 25753 70975
rect 25799 70929 25857 70975
rect 25903 70929 25961 70975
rect 26007 70929 26065 70975
rect 26111 70929 26169 70975
rect 26215 70929 26273 70975
rect 26319 70929 26377 70975
rect 26423 70929 26481 70975
rect 26527 70929 26585 70975
rect 26631 70929 26689 70975
rect 26735 70929 26793 70975
rect 26839 70929 26897 70975
rect 26943 70929 27001 70975
rect 27047 70929 27105 70975
rect 27151 70929 27209 70975
rect 27255 70929 27313 70975
rect 27359 70929 27417 70975
rect 27463 70929 27521 70975
rect 27567 70929 27625 70975
rect 27671 70929 27729 70975
rect 27775 70929 27833 70975
rect 27879 70929 27937 70975
rect 27983 70929 28041 70975
rect 28087 70929 28145 70975
rect 28191 70929 28249 70975
rect 28295 70929 28353 70975
rect 28399 70929 28457 70975
rect 28503 70929 28561 70975
rect 28607 70929 28665 70975
rect 28711 70929 28769 70975
rect 28815 70929 28873 70975
rect 28919 70929 28977 70975
rect 29023 70929 29081 70975
rect 29127 70929 29185 70975
rect 29231 70929 29289 70975
rect 29335 70929 29393 70975
rect 29439 70929 29497 70975
rect 29543 70929 29601 70975
rect 29647 70929 29705 70975
rect 29751 70929 29809 70975
rect 29855 70929 29913 70975
rect 29959 70929 30017 70975
rect 30063 70929 30121 70975
rect 30167 70929 30225 70975
rect 30271 70929 30329 70975
rect 30375 70929 30433 70975
rect 30479 70929 30537 70975
rect 30583 70929 30641 70975
rect 30687 70929 30745 70975
rect 30791 70929 30849 70975
rect 30895 70929 30953 70975
rect 30999 70929 31057 70975
rect 31103 70929 31161 70975
rect 31207 70929 31265 70975
rect 31311 70929 31369 70975
rect 31415 70929 31473 70975
rect 31519 70929 31577 70975
rect 31623 70929 31681 70975
rect 31727 70929 31785 70975
rect 31831 70929 31889 70975
rect 31935 70929 31993 70975
rect 32039 70929 32097 70975
rect 32143 70929 32201 70975
rect 32247 70929 32305 70975
rect 32351 70929 32409 70975
rect 32455 70929 32513 70975
rect 32559 70929 32617 70975
rect 32663 70929 32721 70975
rect 32767 70929 32825 70975
rect 32871 70929 32929 70975
rect 32975 70929 33033 70975
rect 33079 70929 33137 70975
rect 33183 70929 33241 70975
rect 33287 70929 33345 70975
rect 33391 70929 33449 70975
rect 33495 70929 33553 70975
rect 33599 70929 33657 70975
rect 33703 70929 33761 70975
rect 33807 70929 33865 70975
rect 33911 70929 33969 70975
rect 34015 70929 34073 70975
rect 34119 70929 34177 70975
rect 34223 70929 34281 70975
rect 34327 70929 34385 70975
rect 34431 70929 34489 70975
rect 34535 70929 34593 70975
rect 34639 70929 34697 70975
rect 34743 70929 34801 70975
rect 34847 70929 34905 70975
rect 34951 70929 35009 70975
rect 35055 70929 35113 70975
rect 35159 70929 35217 70975
rect 35263 70929 35321 70975
rect 35367 70929 35425 70975
rect 35471 70929 35529 70975
rect 35575 70929 35633 70975
rect 35679 70929 35737 70975
rect 35783 70929 35841 70975
rect 35887 70929 35945 70975
rect 35991 70929 36049 70975
rect 36095 70929 36153 70975
rect 36199 70929 36257 70975
rect 36303 70929 36361 70975
rect 36407 70929 36465 70975
rect 36511 70929 36569 70975
rect 36615 70929 36673 70975
rect 36719 70929 36777 70975
rect 36823 70929 36881 70975
rect 36927 70929 36985 70975
rect 37031 70929 37089 70975
rect 37135 70929 37193 70975
rect 37239 70929 37297 70975
rect 37343 70929 37401 70975
rect 37447 70929 37505 70975
rect 37551 70929 37609 70975
rect 37655 70929 37713 70975
rect 37759 70929 37817 70975
rect 37863 70929 37921 70975
rect 37967 70929 38025 70975
rect 38071 70929 38129 70975
rect 38175 70929 38233 70975
rect 38279 70929 38337 70975
rect 38383 70929 38441 70975
rect 38487 70929 38545 70975
rect 38591 70929 38649 70975
rect 38695 70929 38753 70975
rect 38799 70929 38857 70975
rect 38903 70929 38961 70975
rect 39007 70929 39065 70975
rect 39111 70929 39169 70975
rect 39215 70929 39273 70975
rect 39319 70929 39377 70975
rect 39423 70929 39481 70975
rect 39527 70929 39585 70975
rect 39631 70929 39689 70975
rect 39735 70929 39793 70975
rect 39839 70929 39897 70975
rect 39943 70929 40001 70975
rect 40047 70929 40105 70975
rect 40151 70929 40209 70975
rect 40255 70929 40313 70975
rect 40359 70929 40417 70975
rect 40463 70929 40521 70975
rect 40567 70929 40625 70975
rect 40671 70929 40729 70975
rect 40775 70929 40833 70975
rect 40879 70929 40937 70975
rect 40983 70929 41041 70975
rect 41087 70929 41145 70975
rect 41191 70929 41249 70975
rect 41295 70929 41353 70975
rect 41399 70929 41457 70975
rect 41503 70929 41561 70975
rect 41607 70929 41665 70975
rect 41711 70929 41769 70975
rect 41815 70929 41873 70975
rect 41919 70929 41977 70975
rect 42023 70929 42081 70975
rect 42127 70929 42185 70975
rect 42231 70929 42289 70975
rect 42335 70929 42393 70975
rect 42439 70929 42497 70975
rect 42543 70929 42601 70975
rect 42647 70929 42705 70975
rect 42751 70929 42809 70975
rect 42855 70929 42913 70975
rect 42959 70929 43017 70975
rect 43063 70929 43121 70975
rect 43167 70929 43225 70975
rect 43271 70929 43329 70975
rect 43375 70929 43433 70975
rect 43479 70929 43537 70975
rect 43583 70929 43641 70975
rect 43687 70929 43745 70975
rect 43791 70929 43849 70975
rect 43895 70929 43953 70975
rect 43999 70929 44057 70975
rect 44103 70929 44161 70975
rect 44207 70929 44265 70975
rect 44311 70929 44369 70975
rect 44415 70929 44473 70975
rect 44519 70929 44577 70975
rect 44623 70929 44681 70975
rect 44727 70929 44785 70975
rect 44831 70929 44889 70975
rect 44935 70929 44993 70975
rect 45039 70929 45097 70975
rect 45143 70929 45201 70975
rect 45247 70929 45305 70975
rect 45351 70929 45409 70975
rect 45455 70929 45513 70975
rect 45559 70929 45617 70975
rect 45663 70929 45721 70975
rect 45767 70929 45825 70975
rect 45871 70929 45929 70975
rect 45975 70929 46033 70975
rect 46079 70929 46137 70975
rect 46183 70929 46241 70975
rect 46287 70929 46345 70975
rect 46391 70929 46449 70975
rect 46495 70929 46553 70975
rect 46599 70929 46657 70975
rect 46703 70929 46761 70975
rect 46807 70929 46865 70975
rect 46911 70929 46969 70975
rect 47015 70929 47073 70975
rect 47119 70929 47177 70975
rect 47223 70929 47281 70975
rect 47327 70929 47385 70975
rect 47431 70929 47489 70975
rect 47535 70929 47593 70975
rect 47639 70929 47697 70975
rect 47743 70929 47801 70975
rect 47847 70929 47905 70975
rect 47951 70929 48009 70975
rect 48055 70929 48113 70975
rect 48159 70929 48217 70975
rect 48263 70929 48321 70975
rect 48367 70929 48425 70975
rect 48471 70929 48529 70975
rect 48575 70929 48633 70975
rect 48679 70929 48737 70975
rect 48783 70929 48841 70975
rect 48887 70929 48945 70975
rect 48991 70929 49049 70975
rect 49095 70929 49153 70975
rect 49199 70929 49257 70975
rect 49303 70929 49361 70975
rect 49407 70929 49465 70975
rect 49511 70929 49569 70975
rect 49615 70929 49673 70975
rect 49719 70929 49777 70975
rect 49823 70929 49881 70975
rect 49927 70929 49985 70975
rect 50031 70929 50089 70975
rect 50135 70929 50193 70975
rect 50239 70929 50297 70975
rect 50343 70929 50401 70975
rect 50447 70929 50505 70975
rect 50551 70929 50609 70975
rect 50655 70929 50713 70975
rect 50759 70929 50817 70975
rect 50863 70929 50921 70975
rect 50967 70929 51025 70975
rect 51071 70929 51129 70975
rect 51175 70929 51233 70975
rect 51279 70929 51337 70975
rect 51383 70929 51441 70975
rect 51487 70929 51545 70975
rect 51591 70929 51649 70975
rect 51695 70929 51753 70975
rect 51799 70929 51857 70975
rect 51903 70929 51961 70975
rect 52007 70929 52065 70975
rect 52111 70929 52169 70975
rect 52215 70929 52273 70975
rect 52319 70929 52377 70975
rect 52423 70929 52481 70975
rect 52527 70929 52585 70975
rect 52631 70929 52689 70975
rect 52735 70929 52793 70975
rect 52839 70929 52897 70975
rect 52943 70929 53001 70975
rect 53047 70929 53105 70975
rect 53151 70929 53209 70975
rect 53255 70929 53313 70975
rect 53359 70929 53417 70975
rect 53463 70929 53521 70975
rect 53567 70929 53625 70975
rect 53671 70929 53729 70975
rect 53775 70929 53833 70975
rect 53879 70929 53937 70975
rect 53983 70929 54041 70975
rect 54087 70929 54145 70975
rect 54191 70929 54249 70975
rect 54295 70929 54353 70975
rect 54399 70929 54457 70975
rect 54503 70929 54561 70975
rect 54607 70929 54665 70975
rect 54711 70929 54769 70975
rect 54815 70929 54873 70975
rect 54919 70929 54977 70975
rect 55023 70929 55081 70975
rect 55127 70929 55185 70975
rect 55231 70929 55289 70975
rect 55335 70929 55393 70975
rect 55439 70929 55497 70975
rect 55543 70929 55601 70975
rect 55647 70929 55705 70975
rect 55751 70929 55809 70975
rect 55855 70929 55913 70975
rect 55959 70929 56017 70975
rect 56063 70929 56121 70975
rect 56167 70929 56225 70975
rect 56271 70929 56329 70975
rect 56375 70929 56433 70975
rect 56479 70929 56537 70975
rect 56583 70929 56641 70975
rect 56687 70929 56745 70975
rect 56791 70929 56849 70975
rect 56895 70929 56953 70975
rect 56999 70929 57057 70975
rect 57103 70929 57161 70975
rect 57207 70929 57265 70975
rect 57311 70929 57369 70975
rect 57415 70929 57473 70975
rect 57519 70929 57577 70975
rect 57623 70929 57681 70975
rect 57727 70929 57785 70975
rect 57831 70929 57889 70975
rect 57935 70929 57993 70975
rect 58039 70929 58097 70975
rect 58143 70929 58201 70975
rect 58247 70929 58305 70975
rect 58351 70929 58409 70975
rect 58455 70929 58513 70975
rect 58559 70929 58617 70975
rect 58663 70929 58721 70975
rect 58767 70929 58825 70975
rect 58871 70929 58929 70975
rect 58975 70929 59033 70975
rect 59079 70929 59137 70975
rect 59183 70929 59241 70975
rect 59287 70929 59345 70975
rect 59391 70929 59449 70975
rect 59495 70929 59553 70975
rect 59599 70929 59657 70975
rect 59703 70929 59761 70975
rect 59807 70929 59865 70975
rect 59911 70929 59969 70975
rect 60015 70929 60073 70975
rect 60119 70929 60177 70975
rect 60223 70929 60281 70975
rect 60327 70929 60385 70975
rect 60431 70929 60489 70975
rect 60535 70929 60593 70975
rect 60639 70929 60697 70975
rect 60743 70929 60801 70975
rect 60847 70929 60905 70975
rect 60951 70929 61009 70975
rect 61055 70929 61113 70975
rect 61159 70929 61217 70975
rect 61263 70929 61321 70975
rect 61367 70929 61425 70975
rect 61471 70929 61529 70975
rect 61575 70929 61633 70975
rect 61679 70929 61737 70975
rect 61783 70929 61841 70975
rect 61887 70929 61945 70975
rect 61991 70929 62049 70975
rect 62095 70929 62153 70975
rect 62199 70929 62257 70975
rect 62303 70929 62361 70975
rect 62407 70929 62465 70975
rect 62511 70929 62569 70975
rect 62615 70929 62673 70975
rect 62719 70929 62777 70975
rect 62823 70929 62881 70975
rect 62927 70929 62985 70975
rect 63031 70929 63089 70975
rect 63135 70929 63193 70975
rect 63239 70929 63297 70975
rect 63343 70929 63401 70975
rect 63447 70929 63505 70975
rect 63551 70929 63609 70975
rect 63655 70929 63713 70975
rect 63759 70929 63817 70975
rect 63863 70929 63921 70975
rect 63967 70929 64025 70975
rect 64071 70929 64129 70975
rect 64175 70929 64233 70975
rect 64279 70929 64337 70975
rect 64383 70929 64441 70975
rect 64487 70929 64545 70975
rect 64591 70929 64649 70975
rect 64695 70929 64753 70975
rect 64799 70929 64857 70975
rect 64903 70929 64961 70975
rect 65007 70929 65065 70975
rect 65111 70929 65169 70975
rect 65215 70929 65273 70975
rect 65319 70929 65377 70975
rect 65423 70929 65481 70975
rect 65527 70929 65585 70975
rect 65631 70929 65689 70975
rect 65735 70929 65793 70975
rect 65839 70929 65897 70975
rect 65943 70929 66001 70975
rect 66047 70929 66105 70975
rect 66151 70929 66209 70975
rect 66255 70929 66313 70975
rect 66359 70929 66417 70975
rect 66463 70929 66521 70975
rect 66567 70929 66625 70975
rect 66671 70929 66729 70975
rect 66775 70929 66833 70975
rect 66879 70929 66937 70975
rect 66983 70929 67041 70975
rect 67087 70929 67145 70975
rect 67191 70929 67249 70975
rect 67295 70929 67353 70975
rect 67399 70929 67457 70975
rect 67503 70929 67561 70975
rect 67607 70929 67665 70975
rect 67711 70929 67769 70975
rect 67815 70929 67873 70975
rect 67919 70929 67977 70975
rect 68023 70929 68081 70975
rect 68127 70929 68185 70975
rect 68231 70929 68289 70975
rect 68335 70929 68393 70975
rect 68439 70929 68497 70975
rect 68543 70929 68601 70975
rect 68647 70929 68705 70975
rect 68751 70929 68809 70975
rect 68855 70929 68913 70975
rect 68959 70929 69017 70975
rect 69063 70929 69121 70975
rect 69167 70929 69225 70975
rect 69271 70929 69329 70975
rect 69375 70929 69433 70975
rect 69479 70929 69537 70975
rect 69583 70929 69641 70975
rect 69687 70929 69745 70975
rect 69791 70929 69849 70975
rect 69895 70929 69957 70975
rect 13108 70871 69957 70929
rect 13108 70825 13119 70871
rect 13165 70825 13223 70871
rect 13269 70825 13377 70871
rect 13423 70825 13481 70871
rect 13527 70825 13585 70871
rect 13631 70825 13689 70871
rect 13735 70825 13793 70871
rect 13839 70825 13897 70871
rect 13943 70825 14001 70871
rect 14047 70825 14105 70871
rect 14151 70825 14209 70871
rect 14255 70825 14313 70871
rect 14359 70825 14417 70871
rect 14463 70825 14521 70871
rect 14567 70825 14625 70871
rect 14671 70825 14729 70871
rect 14775 70825 14833 70871
rect 14879 70825 14937 70871
rect 14983 70825 15041 70871
rect 15087 70825 15145 70871
rect 15191 70825 15249 70871
rect 15295 70825 15353 70871
rect 15399 70825 15457 70871
rect 15503 70825 15561 70871
rect 15607 70825 15665 70871
rect 15711 70825 15769 70871
rect 15815 70825 15873 70871
rect 15919 70825 15977 70871
rect 16023 70825 16081 70871
rect 16127 70825 16185 70871
rect 16231 70825 16289 70871
rect 16335 70825 16393 70871
rect 16439 70825 16497 70871
rect 16543 70825 16601 70871
rect 16647 70825 16705 70871
rect 16751 70825 16809 70871
rect 16855 70825 16913 70871
rect 16959 70825 17017 70871
rect 17063 70825 17121 70871
rect 17167 70825 17225 70871
rect 17271 70825 17329 70871
rect 17375 70825 17433 70871
rect 17479 70825 17537 70871
rect 17583 70825 17641 70871
rect 17687 70825 17745 70871
rect 17791 70825 17849 70871
rect 17895 70825 17953 70871
rect 17999 70825 18057 70871
rect 18103 70825 18161 70871
rect 18207 70825 18265 70871
rect 18311 70825 18369 70871
rect 18415 70825 18473 70871
rect 18519 70825 18577 70871
rect 18623 70825 18681 70871
rect 18727 70825 18785 70871
rect 18831 70825 18889 70871
rect 18935 70825 18993 70871
rect 19039 70825 19097 70871
rect 19143 70825 19201 70871
rect 19247 70825 19305 70871
rect 19351 70825 19409 70871
rect 19455 70825 19513 70871
rect 19559 70825 19617 70871
rect 19663 70825 19721 70871
rect 19767 70825 19825 70871
rect 19871 70825 19929 70871
rect 19975 70825 20033 70871
rect 20079 70825 20137 70871
rect 20183 70825 20241 70871
rect 20287 70825 20345 70871
rect 20391 70825 20449 70871
rect 20495 70825 20553 70871
rect 20599 70825 20657 70871
rect 20703 70825 20761 70871
rect 20807 70825 20865 70871
rect 20911 70825 20969 70871
rect 21015 70825 21073 70871
rect 21119 70825 21177 70871
rect 21223 70825 21281 70871
rect 21327 70825 21385 70871
rect 21431 70825 21489 70871
rect 21535 70825 21593 70871
rect 21639 70825 21697 70871
rect 21743 70825 21801 70871
rect 21847 70825 21905 70871
rect 21951 70825 22009 70871
rect 22055 70825 22113 70871
rect 22159 70825 22217 70871
rect 22263 70825 22321 70871
rect 22367 70825 22425 70871
rect 22471 70825 22529 70871
rect 22575 70825 22633 70871
rect 22679 70825 22737 70871
rect 22783 70825 22841 70871
rect 22887 70825 22945 70871
rect 22991 70825 23049 70871
rect 23095 70825 23153 70871
rect 23199 70825 23257 70871
rect 23303 70825 23361 70871
rect 23407 70825 23465 70871
rect 23511 70825 23569 70871
rect 23615 70825 23673 70871
rect 23719 70825 23777 70871
rect 23823 70825 23881 70871
rect 23927 70825 23985 70871
rect 24031 70825 24089 70871
rect 24135 70825 24193 70871
rect 24239 70825 24297 70871
rect 24343 70825 24401 70871
rect 24447 70825 24505 70871
rect 24551 70825 24609 70871
rect 24655 70825 24713 70871
rect 24759 70825 24817 70871
rect 24863 70825 24921 70871
rect 24967 70825 25025 70871
rect 25071 70825 25129 70871
rect 25175 70825 25233 70871
rect 25279 70825 25337 70871
rect 25383 70825 25441 70871
rect 25487 70825 25545 70871
rect 25591 70825 25649 70871
rect 25695 70825 25753 70871
rect 25799 70825 25857 70871
rect 25903 70825 25961 70871
rect 26007 70825 26065 70871
rect 26111 70825 26169 70871
rect 26215 70825 26273 70871
rect 26319 70825 26377 70871
rect 26423 70825 26481 70871
rect 26527 70825 26585 70871
rect 26631 70825 26689 70871
rect 26735 70825 26793 70871
rect 26839 70825 26897 70871
rect 26943 70825 27001 70871
rect 27047 70825 27105 70871
rect 27151 70825 27209 70871
rect 27255 70825 27313 70871
rect 27359 70825 27417 70871
rect 27463 70825 27521 70871
rect 27567 70825 27625 70871
rect 27671 70825 27729 70871
rect 27775 70825 27833 70871
rect 27879 70825 27937 70871
rect 27983 70825 28041 70871
rect 28087 70825 28145 70871
rect 28191 70825 28249 70871
rect 28295 70825 28353 70871
rect 28399 70825 28457 70871
rect 28503 70825 28561 70871
rect 28607 70825 28665 70871
rect 28711 70825 28769 70871
rect 28815 70825 28873 70871
rect 28919 70825 28977 70871
rect 29023 70825 29081 70871
rect 29127 70825 29185 70871
rect 29231 70825 29289 70871
rect 29335 70825 29393 70871
rect 29439 70825 29497 70871
rect 29543 70825 29601 70871
rect 29647 70825 29705 70871
rect 29751 70825 29809 70871
rect 29855 70825 29913 70871
rect 29959 70825 30017 70871
rect 30063 70825 30121 70871
rect 30167 70825 30225 70871
rect 30271 70825 30329 70871
rect 30375 70825 30433 70871
rect 30479 70825 30537 70871
rect 30583 70825 30641 70871
rect 30687 70825 30745 70871
rect 30791 70825 30849 70871
rect 30895 70825 30953 70871
rect 30999 70825 31057 70871
rect 31103 70825 31161 70871
rect 31207 70825 31265 70871
rect 31311 70825 31369 70871
rect 31415 70825 31473 70871
rect 31519 70825 31577 70871
rect 31623 70825 31681 70871
rect 31727 70825 31785 70871
rect 31831 70825 31889 70871
rect 31935 70825 31993 70871
rect 32039 70825 32097 70871
rect 32143 70825 32201 70871
rect 32247 70825 32305 70871
rect 32351 70825 32409 70871
rect 32455 70825 32513 70871
rect 32559 70825 32617 70871
rect 32663 70825 32721 70871
rect 32767 70825 32825 70871
rect 32871 70825 32929 70871
rect 32975 70825 33033 70871
rect 33079 70825 33137 70871
rect 33183 70825 33241 70871
rect 33287 70825 33345 70871
rect 33391 70825 33449 70871
rect 33495 70825 33553 70871
rect 33599 70825 33657 70871
rect 33703 70825 33761 70871
rect 33807 70825 33865 70871
rect 33911 70825 33969 70871
rect 34015 70825 34073 70871
rect 34119 70825 34177 70871
rect 34223 70825 34281 70871
rect 34327 70825 34385 70871
rect 34431 70825 34489 70871
rect 34535 70825 34593 70871
rect 34639 70825 34697 70871
rect 34743 70825 34801 70871
rect 34847 70825 34905 70871
rect 34951 70825 35009 70871
rect 35055 70825 35113 70871
rect 35159 70825 35217 70871
rect 35263 70825 35321 70871
rect 35367 70825 35425 70871
rect 35471 70825 35529 70871
rect 35575 70825 35633 70871
rect 35679 70825 35737 70871
rect 35783 70825 35841 70871
rect 35887 70825 35945 70871
rect 35991 70825 36049 70871
rect 36095 70825 36153 70871
rect 36199 70825 36257 70871
rect 36303 70825 36361 70871
rect 36407 70825 36465 70871
rect 36511 70825 36569 70871
rect 36615 70825 36673 70871
rect 36719 70825 36777 70871
rect 36823 70825 36881 70871
rect 36927 70825 36985 70871
rect 37031 70825 37089 70871
rect 37135 70825 37193 70871
rect 37239 70825 37297 70871
rect 37343 70825 37401 70871
rect 37447 70825 37505 70871
rect 37551 70825 37609 70871
rect 37655 70825 37713 70871
rect 37759 70825 37817 70871
rect 37863 70825 37921 70871
rect 37967 70825 38025 70871
rect 38071 70825 38129 70871
rect 38175 70825 38233 70871
rect 38279 70825 38337 70871
rect 38383 70825 38441 70871
rect 38487 70825 38545 70871
rect 38591 70825 38649 70871
rect 38695 70825 38753 70871
rect 38799 70825 38857 70871
rect 38903 70825 38961 70871
rect 39007 70825 39065 70871
rect 39111 70825 39169 70871
rect 39215 70825 39273 70871
rect 39319 70825 39377 70871
rect 39423 70825 39481 70871
rect 39527 70825 39585 70871
rect 39631 70825 39689 70871
rect 39735 70825 39793 70871
rect 39839 70825 39897 70871
rect 39943 70825 40001 70871
rect 40047 70825 40105 70871
rect 40151 70825 40209 70871
rect 40255 70825 40313 70871
rect 40359 70825 40417 70871
rect 40463 70825 40521 70871
rect 40567 70825 40625 70871
rect 40671 70825 40729 70871
rect 40775 70825 40833 70871
rect 40879 70825 40937 70871
rect 40983 70825 41041 70871
rect 41087 70825 41145 70871
rect 41191 70825 41249 70871
rect 41295 70825 41353 70871
rect 41399 70825 41457 70871
rect 41503 70825 41561 70871
rect 41607 70825 41665 70871
rect 41711 70825 41769 70871
rect 41815 70825 41873 70871
rect 41919 70825 41977 70871
rect 42023 70825 42081 70871
rect 42127 70825 42185 70871
rect 42231 70825 42289 70871
rect 42335 70825 42393 70871
rect 42439 70825 42497 70871
rect 42543 70825 42601 70871
rect 42647 70825 42705 70871
rect 42751 70825 42809 70871
rect 42855 70825 42913 70871
rect 42959 70825 43017 70871
rect 43063 70825 43121 70871
rect 43167 70825 43225 70871
rect 43271 70825 43329 70871
rect 43375 70825 43433 70871
rect 43479 70825 43537 70871
rect 43583 70825 43641 70871
rect 43687 70825 43745 70871
rect 43791 70825 43849 70871
rect 43895 70825 43953 70871
rect 43999 70825 44057 70871
rect 44103 70825 44161 70871
rect 44207 70825 44265 70871
rect 44311 70825 44369 70871
rect 44415 70825 44473 70871
rect 44519 70825 44577 70871
rect 44623 70825 44681 70871
rect 44727 70825 44785 70871
rect 44831 70825 44889 70871
rect 44935 70825 44993 70871
rect 45039 70825 45097 70871
rect 45143 70825 45201 70871
rect 45247 70825 45305 70871
rect 45351 70825 45409 70871
rect 45455 70825 45513 70871
rect 45559 70825 45617 70871
rect 45663 70825 45721 70871
rect 45767 70825 45825 70871
rect 45871 70825 45929 70871
rect 45975 70825 46033 70871
rect 46079 70825 46137 70871
rect 46183 70825 46241 70871
rect 46287 70825 46345 70871
rect 46391 70825 46449 70871
rect 46495 70825 46553 70871
rect 46599 70825 46657 70871
rect 46703 70825 46761 70871
rect 46807 70825 46865 70871
rect 46911 70825 46969 70871
rect 47015 70825 47073 70871
rect 47119 70825 47177 70871
rect 47223 70825 47281 70871
rect 47327 70825 47385 70871
rect 47431 70825 47489 70871
rect 47535 70825 47593 70871
rect 47639 70825 47697 70871
rect 47743 70825 47801 70871
rect 47847 70825 47905 70871
rect 47951 70825 48009 70871
rect 48055 70825 48113 70871
rect 48159 70825 48217 70871
rect 48263 70825 48321 70871
rect 48367 70825 48425 70871
rect 48471 70825 48529 70871
rect 48575 70825 48633 70871
rect 48679 70825 48737 70871
rect 48783 70825 48841 70871
rect 48887 70825 48945 70871
rect 48991 70825 49049 70871
rect 49095 70825 49153 70871
rect 49199 70825 49257 70871
rect 49303 70825 49361 70871
rect 49407 70825 49465 70871
rect 49511 70825 49569 70871
rect 49615 70825 49673 70871
rect 49719 70825 49777 70871
rect 49823 70825 49881 70871
rect 49927 70825 49985 70871
rect 50031 70825 50089 70871
rect 50135 70825 50193 70871
rect 50239 70825 50297 70871
rect 50343 70825 50401 70871
rect 50447 70825 50505 70871
rect 50551 70825 50609 70871
rect 50655 70825 50713 70871
rect 50759 70825 50817 70871
rect 50863 70825 50921 70871
rect 50967 70825 51025 70871
rect 51071 70825 51129 70871
rect 51175 70825 51233 70871
rect 51279 70825 51337 70871
rect 51383 70825 51441 70871
rect 51487 70825 51545 70871
rect 51591 70825 51649 70871
rect 51695 70825 51753 70871
rect 51799 70825 51857 70871
rect 51903 70825 51961 70871
rect 52007 70825 52065 70871
rect 52111 70825 52169 70871
rect 52215 70825 52273 70871
rect 52319 70825 52377 70871
rect 52423 70825 52481 70871
rect 52527 70825 52585 70871
rect 52631 70825 52689 70871
rect 52735 70825 52793 70871
rect 52839 70825 52897 70871
rect 52943 70825 53001 70871
rect 53047 70825 53105 70871
rect 53151 70825 53209 70871
rect 53255 70825 53313 70871
rect 53359 70825 53417 70871
rect 53463 70825 53521 70871
rect 53567 70825 53625 70871
rect 53671 70825 53729 70871
rect 53775 70825 53833 70871
rect 53879 70825 53937 70871
rect 53983 70825 54041 70871
rect 54087 70825 54145 70871
rect 54191 70825 54249 70871
rect 54295 70825 54353 70871
rect 54399 70825 54457 70871
rect 54503 70825 54561 70871
rect 54607 70825 54665 70871
rect 54711 70825 54769 70871
rect 54815 70825 54873 70871
rect 54919 70825 54977 70871
rect 55023 70825 55081 70871
rect 55127 70825 55185 70871
rect 55231 70825 55289 70871
rect 55335 70825 55393 70871
rect 55439 70825 55497 70871
rect 55543 70825 55601 70871
rect 55647 70825 55705 70871
rect 55751 70825 55809 70871
rect 55855 70825 55913 70871
rect 55959 70825 56017 70871
rect 56063 70825 56121 70871
rect 56167 70825 56225 70871
rect 56271 70825 56329 70871
rect 56375 70825 56433 70871
rect 56479 70825 56537 70871
rect 56583 70825 56641 70871
rect 56687 70825 56745 70871
rect 56791 70825 56849 70871
rect 56895 70825 56953 70871
rect 56999 70825 57057 70871
rect 57103 70825 57161 70871
rect 57207 70825 57265 70871
rect 57311 70825 57369 70871
rect 57415 70825 57473 70871
rect 57519 70825 57577 70871
rect 57623 70825 57681 70871
rect 57727 70825 57785 70871
rect 57831 70825 57889 70871
rect 57935 70825 57993 70871
rect 58039 70825 58097 70871
rect 58143 70825 58201 70871
rect 58247 70825 58305 70871
rect 58351 70825 58409 70871
rect 58455 70825 58513 70871
rect 58559 70825 58617 70871
rect 58663 70825 58721 70871
rect 58767 70825 58825 70871
rect 58871 70825 58929 70871
rect 58975 70825 59033 70871
rect 59079 70825 59137 70871
rect 59183 70825 59241 70871
rect 59287 70825 59345 70871
rect 59391 70825 59449 70871
rect 59495 70825 59553 70871
rect 59599 70825 59657 70871
rect 59703 70825 59761 70871
rect 59807 70825 59865 70871
rect 59911 70825 59969 70871
rect 60015 70825 60073 70871
rect 60119 70825 60177 70871
rect 60223 70825 60281 70871
rect 60327 70825 60385 70871
rect 60431 70825 60489 70871
rect 60535 70825 60593 70871
rect 60639 70825 60697 70871
rect 60743 70825 60801 70871
rect 60847 70825 60905 70871
rect 60951 70825 61009 70871
rect 61055 70825 61113 70871
rect 61159 70825 61217 70871
rect 61263 70825 61321 70871
rect 61367 70825 61425 70871
rect 61471 70825 61529 70871
rect 61575 70825 61633 70871
rect 61679 70825 61737 70871
rect 61783 70825 61841 70871
rect 61887 70825 61945 70871
rect 61991 70825 62049 70871
rect 62095 70825 62153 70871
rect 62199 70825 62257 70871
rect 62303 70825 62361 70871
rect 62407 70825 62465 70871
rect 62511 70825 62569 70871
rect 62615 70825 62673 70871
rect 62719 70825 62777 70871
rect 62823 70825 62881 70871
rect 62927 70825 62985 70871
rect 63031 70825 63089 70871
rect 63135 70825 63193 70871
rect 63239 70825 63297 70871
rect 63343 70825 63401 70871
rect 63447 70825 63505 70871
rect 63551 70825 63609 70871
rect 63655 70825 63713 70871
rect 63759 70825 63817 70871
rect 63863 70825 63921 70871
rect 63967 70825 64025 70871
rect 64071 70825 64129 70871
rect 64175 70825 64233 70871
rect 64279 70825 64337 70871
rect 64383 70825 64441 70871
rect 64487 70825 64545 70871
rect 64591 70825 64649 70871
rect 64695 70825 64753 70871
rect 64799 70825 64857 70871
rect 64903 70825 64961 70871
rect 65007 70825 65065 70871
rect 65111 70825 65169 70871
rect 65215 70825 65273 70871
rect 65319 70825 65377 70871
rect 65423 70825 65481 70871
rect 65527 70825 65585 70871
rect 65631 70825 65689 70871
rect 65735 70825 65793 70871
rect 65839 70825 65897 70871
rect 65943 70825 66001 70871
rect 66047 70825 66105 70871
rect 66151 70825 66209 70871
rect 66255 70825 66313 70871
rect 66359 70825 66417 70871
rect 66463 70825 66521 70871
rect 66567 70825 66625 70871
rect 66671 70825 66729 70871
rect 66775 70825 66833 70871
rect 66879 70825 66937 70871
rect 66983 70825 67041 70871
rect 67087 70825 67145 70871
rect 67191 70825 67249 70871
rect 67295 70825 67353 70871
rect 67399 70825 67457 70871
rect 67503 70825 67561 70871
rect 67607 70825 67665 70871
rect 67711 70825 67769 70871
rect 67815 70825 67873 70871
rect 67919 70825 67977 70871
rect 68023 70825 68081 70871
rect 68127 70825 68185 70871
rect 68231 70825 68289 70871
rect 68335 70825 68393 70871
rect 68439 70825 68497 70871
rect 68543 70825 68601 70871
rect 68647 70825 68705 70871
rect 68751 70825 68809 70871
rect 68855 70825 68913 70871
rect 68959 70825 69017 70871
rect 69063 70825 69121 70871
rect 69167 70825 69225 70871
rect 69271 70825 69329 70871
rect 69375 70825 69433 70871
rect 69479 70825 69537 70871
rect 69583 70825 69641 70871
rect 69687 70825 69745 70871
rect 69791 70825 69849 70871
rect 69895 70825 69957 70871
rect 13108 70814 69957 70825
rect 13108 70767 13280 70814
rect 13108 70721 13119 70767
rect 13165 70721 13223 70767
rect 13269 70721 13280 70767
rect 13108 70663 13280 70721
rect 13108 70617 13119 70663
rect 13165 70617 13223 70663
rect 13269 70617 13280 70663
rect 13108 70559 13280 70617
rect 13108 70513 13119 70559
rect 13165 70513 13223 70559
rect 13269 70513 13280 70559
rect 13108 70455 13280 70513
rect 13108 70409 13119 70455
rect 13165 70409 13223 70455
rect 13269 70409 13280 70455
rect 13108 70351 13280 70409
rect 13108 70305 13119 70351
rect 13165 70305 13223 70351
rect 13269 70305 13280 70351
rect 13108 70247 13280 70305
rect 13108 70201 13119 70247
rect 13165 70201 13223 70247
rect 13269 70201 13280 70247
rect 13108 70143 13280 70201
rect 13108 70097 13119 70143
rect 13165 70097 13223 70143
rect 13269 70097 13280 70143
rect 13108 70039 13280 70097
rect 13108 69993 13119 70039
rect 13165 69993 13223 70039
rect 13269 69993 13280 70039
rect 13108 69935 13280 69993
rect 13108 69889 13119 69935
rect 13165 69889 13223 69935
rect 13269 69889 13280 69935
rect 13108 69831 13280 69889
rect 13108 69785 13119 69831
rect 13165 69785 13223 69831
rect 13269 69785 13280 69831
rect 69785 70720 69957 70814
rect 69785 70674 69796 70720
rect 69842 70674 69900 70720
rect 69946 70674 69957 70720
rect 69785 70616 69957 70674
rect 69785 70570 69796 70616
rect 69842 70570 69900 70616
rect 69946 70570 69957 70616
rect 69785 70512 69957 70570
rect 69785 70466 69796 70512
rect 69842 70466 69900 70512
rect 69946 70466 69957 70512
rect 69785 70408 69957 70466
rect 69785 70362 69796 70408
rect 69842 70362 69900 70408
rect 69946 70362 69957 70408
rect 69785 70304 69957 70362
rect 69785 70258 69796 70304
rect 69842 70258 69900 70304
rect 69946 70258 69957 70304
rect 69785 70200 69957 70258
rect 69785 70154 69796 70200
rect 69842 70154 69900 70200
rect 69946 70154 69957 70200
rect 69785 70096 69957 70154
rect 69785 70050 69796 70096
rect 69842 70050 69900 70096
rect 69946 70050 69957 70096
rect 69785 69957 69957 70050
rect 69785 69946 71000 69957
rect 69785 69900 69796 69946
rect 69842 69900 69900 69946
rect 69946 69900 70004 69946
rect 70050 69900 70108 69946
rect 70154 69900 70212 69946
rect 70258 69900 70316 69946
rect 70362 69900 70420 69946
rect 70466 69900 70524 69946
rect 70570 69900 70628 69946
rect 70674 69908 71000 69946
rect 70674 69900 70824 69908
rect 69785 69862 70824 69900
rect 70870 69862 70928 69908
rect 70974 69862 71000 69908
rect 69785 69842 71000 69862
rect 69785 69796 69796 69842
rect 69842 69796 69900 69842
rect 69946 69796 70004 69842
rect 70050 69796 70108 69842
rect 70154 69796 70212 69842
rect 70258 69796 70316 69842
rect 70362 69796 70420 69842
rect 70466 69796 70524 69842
rect 70570 69796 70628 69842
rect 70674 69804 71000 69842
rect 70674 69796 70824 69804
rect 69785 69785 70824 69796
rect 13108 69727 13280 69785
rect 13108 69681 13119 69727
rect 13165 69681 13223 69727
rect 13269 69681 13280 69727
rect 13108 69623 13280 69681
rect 13108 69577 13119 69623
rect 13165 69577 13223 69623
rect 13269 69577 13280 69623
rect 13108 69519 13280 69577
rect 13108 69473 13119 69519
rect 13165 69473 13223 69519
rect 13269 69473 13280 69519
rect 13108 69415 13280 69473
rect 13108 69369 13119 69415
rect 13165 69369 13223 69415
rect 13269 69369 13280 69415
rect 13108 69311 13280 69369
rect 13108 69265 13119 69311
rect 13165 69265 13223 69311
rect 13269 69265 13280 69311
rect 13108 69207 13280 69265
rect 13108 69161 13119 69207
rect 13165 69161 13223 69207
rect 13269 69161 13280 69207
rect 13108 69103 13280 69161
rect 13108 69057 13119 69103
rect 13165 69057 13223 69103
rect 13269 69057 13280 69103
rect 13108 68999 13280 69057
rect 13108 68953 13119 68999
rect 13165 68953 13223 68999
rect 13269 68953 13280 68999
rect 13108 68895 13280 68953
rect 13108 68849 13119 68895
rect 13165 68849 13223 68895
rect 13269 68849 13280 68895
rect 13108 68791 13280 68849
rect 13108 68745 13119 68791
rect 13165 68745 13223 68791
rect 13269 68745 13280 68791
rect 13108 68687 13280 68745
rect 13108 68641 13119 68687
rect 13165 68641 13223 68687
rect 13269 68641 13280 68687
rect 13108 68583 13280 68641
rect 13108 68537 13119 68583
rect 13165 68537 13223 68583
rect 13269 68537 13280 68583
rect 13108 68479 13280 68537
rect 13108 68433 13119 68479
rect 13165 68433 13223 68479
rect 13269 68433 13280 68479
rect 13108 68375 13280 68433
rect 13108 68329 13119 68375
rect 13165 68329 13223 68375
rect 13269 68329 13280 68375
rect 13108 68271 13280 68329
rect 13108 68225 13119 68271
rect 13165 68225 13223 68271
rect 13269 68225 13280 68271
rect 13108 68167 13280 68225
rect 13108 68121 13119 68167
rect 13165 68121 13223 68167
rect 13269 68121 13280 68167
rect 13108 68063 13280 68121
rect 13108 68017 13119 68063
rect 13165 68017 13223 68063
rect 13269 68017 13280 68063
rect 13108 67959 13280 68017
rect 13108 67913 13119 67959
rect 13165 67913 13223 67959
rect 13269 67913 13280 67959
rect 13108 67855 13280 67913
rect 13108 67809 13119 67855
rect 13165 67809 13223 67855
rect 13269 67809 13280 67855
rect 13108 67751 13280 67809
rect 13108 67705 13119 67751
rect 13165 67705 13223 67751
rect 13269 67705 13280 67751
rect 13108 67647 13280 67705
rect 13108 67601 13119 67647
rect 13165 67601 13223 67647
rect 13269 67601 13280 67647
rect 13108 67543 13280 67601
rect 13108 67497 13119 67543
rect 13165 67497 13223 67543
rect 13269 67497 13280 67543
rect 13108 67439 13280 67497
rect 13108 67393 13119 67439
rect 13165 67393 13223 67439
rect 13269 67393 13280 67439
rect 13108 67335 13280 67393
rect 13108 67289 13119 67335
rect 13165 67289 13223 67335
rect 13269 67289 13280 67335
rect 13108 67231 13280 67289
rect 13108 67185 13119 67231
rect 13165 67185 13223 67231
rect 13269 67185 13280 67231
rect 13108 67127 13280 67185
rect 13108 67081 13119 67127
rect 13165 67081 13223 67127
rect 13269 67081 13280 67127
rect 13108 67023 13280 67081
rect 13108 66977 13119 67023
rect 13165 66977 13223 67023
rect 13269 66977 13280 67023
rect 13108 66919 13280 66977
rect 13108 66873 13119 66919
rect 13165 66873 13223 66919
rect 13269 66873 13280 66919
rect 13108 66815 13280 66873
rect 13108 66769 13119 66815
rect 13165 66769 13223 66815
rect 13269 66769 13280 66815
rect 13108 66711 13280 66769
rect 13108 66665 13119 66711
rect 13165 66665 13223 66711
rect 13269 66665 13280 66711
rect 13108 66607 13280 66665
rect 13108 66561 13119 66607
rect 13165 66561 13223 66607
rect 13269 66561 13280 66607
rect 13108 66503 13280 66561
rect 13108 66457 13119 66503
rect 13165 66457 13223 66503
rect 13269 66457 13280 66503
rect 13108 66399 13280 66457
rect 13108 66353 13119 66399
rect 13165 66353 13223 66399
rect 13269 66353 13280 66399
rect 13108 66295 13280 66353
rect 13108 66249 13119 66295
rect 13165 66249 13223 66295
rect 13269 66249 13280 66295
rect 13108 66191 13280 66249
rect 13108 66145 13119 66191
rect 13165 66145 13223 66191
rect 13269 66145 13280 66191
rect 13108 66087 13280 66145
rect 13108 66041 13119 66087
rect 13165 66041 13223 66087
rect 13269 66041 13280 66087
rect 13108 65983 13280 66041
rect 13108 65937 13119 65983
rect 13165 65937 13223 65983
rect 13269 65937 13280 65983
rect 13108 65879 13280 65937
rect 13108 65833 13119 65879
rect 13165 65833 13223 65879
rect 13269 65833 13280 65879
rect 13108 65775 13280 65833
rect 13108 65729 13119 65775
rect 13165 65729 13223 65775
rect 13269 65729 13280 65775
rect 13108 65671 13280 65729
rect 13108 65625 13119 65671
rect 13165 65625 13223 65671
rect 13269 65625 13280 65671
rect 13108 65567 13280 65625
rect 13108 65521 13119 65567
rect 13165 65521 13223 65567
rect 13269 65521 13280 65567
rect 13108 65463 13280 65521
rect 13108 65417 13119 65463
rect 13165 65417 13223 65463
rect 13269 65417 13280 65463
rect 13108 65359 13280 65417
rect 13108 65313 13119 65359
rect 13165 65313 13223 65359
rect 13269 65313 13280 65359
rect 13108 65255 13280 65313
rect 13108 65209 13119 65255
rect 13165 65209 13223 65255
rect 13269 65209 13280 65255
rect 13108 65151 13280 65209
rect 13108 65105 13119 65151
rect 13165 65105 13223 65151
rect 13269 65105 13280 65151
rect 13108 65047 13280 65105
rect 13108 65001 13119 65047
rect 13165 65001 13223 65047
rect 13269 65001 13280 65047
rect 13108 64943 13280 65001
rect 13108 64897 13119 64943
rect 13165 64897 13223 64943
rect 13269 64897 13280 64943
rect 13108 64839 13280 64897
rect 13108 64793 13119 64839
rect 13165 64793 13223 64839
rect 13269 64793 13280 64839
rect 13108 64735 13280 64793
rect 13108 64689 13119 64735
rect 13165 64689 13223 64735
rect 13269 64689 13280 64735
rect 13108 64631 13280 64689
rect 13108 64585 13119 64631
rect 13165 64585 13223 64631
rect 13269 64585 13280 64631
rect 13108 64527 13280 64585
rect 13108 64481 13119 64527
rect 13165 64481 13223 64527
rect 13269 64481 13280 64527
rect 13108 64423 13280 64481
rect 13108 64377 13119 64423
rect 13165 64377 13223 64423
rect 13269 64377 13280 64423
rect 13108 64319 13280 64377
rect 13108 64273 13119 64319
rect 13165 64273 13223 64319
rect 13269 64273 13280 64319
rect 13108 64215 13280 64273
rect 13108 64169 13119 64215
rect 13165 64169 13223 64215
rect 13269 64169 13280 64215
rect 13108 64111 13280 64169
rect 13108 64065 13119 64111
rect 13165 64065 13223 64111
rect 13269 64065 13280 64111
rect 13108 64007 13280 64065
rect 13108 63961 13119 64007
rect 13165 63961 13223 64007
rect 13269 63961 13280 64007
rect 13108 63903 13280 63961
rect 13108 63857 13119 63903
rect 13165 63857 13223 63903
rect 13269 63857 13280 63903
rect 13108 63799 13280 63857
rect 13108 63753 13119 63799
rect 13165 63753 13223 63799
rect 13269 63753 13280 63799
rect 13108 63695 13280 63753
rect 13108 63649 13119 63695
rect 13165 63649 13223 63695
rect 13269 63649 13280 63695
rect 13108 63591 13280 63649
rect 13108 63545 13119 63591
rect 13165 63545 13223 63591
rect 13269 63545 13280 63591
rect 13108 63487 13280 63545
rect 13108 63441 13119 63487
rect 13165 63441 13223 63487
rect 13269 63441 13280 63487
rect 13108 63383 13280 63441
rect 13108 63337 13119 63383
rect 13165 63337 13223 63383
rect 13269 63337 13280 63383
rect 13108 63279 13280 63337
rect 13108 63233 13119 63279
rect 13165 63233 13223 63279
rect 13269 63233 13280 63279
rect 13108 63175 13280 63233
rect 13108 63129 13119 63175
rect 13165 63129 13223 63175
rect 13269 63129 13280 63175
rect 13108 63071 13280 63129
rect 13108 63025 13119 63071
rect 13165 63025 13223 63071
rect 13269 63025 13280 63071
rect 13108 62967 13280 63025
rect 13108 62921 13119 62967
rect 13165 62921 13223 62967
rect 13269 62921 13280 62967
rect 13108 62863 13280 62921
rect 13108 62817 13119 62863
rect 13165 62817 13223 62863
rect 13269 62817 13280 62863
rect 13108 62759 13280 62817
rect 13108 62713 13119 62759
rect 13165 62713 13223 62759
rect 13269 62713 13280 62759
rect 13108 62655 13280 62713
rect 13108 62609 13119 62655
rect 13165 62609 13223 62655
rect 13269 62609 13280 62655
rect 13108 62551 13280 62609
rect 13108 62505 13119 62551
rect 13165 62505 13223 62551
rect 13269 62505 13280 62551
rect 13108 62447 13280 62505
rect 13108 62401 13119 62447
rect 13165 62401 13223 62447
rect 13269 62401 13280 62447
rect 13108 62343 13280 62401
rect 13108 62297 13119 62343
rect 13165 62297 13223 62343
rect 13269 62297 13280 62343
rect 13108 62239 13280 62297
rect 13108 62193 13119 62239
rect 13165 62193 13223 62239
rect 13269 62193 13280 62239
rect 13108 62135 13280 62193
rect 13108 62089 13119 62135
rect 13165 62089 13223 62135
rect 13269 62089 13280 62135
rect 13108 62031 13280 62089
rect 13108 61985 13119 62031
rect 13165 61985 13223 62031
rect 13269 61985 13280 62031
rect 13108 61927 13280 61985
rect 13108 61881 13119 61927
rect 13165 61881 13223 61927
rect 13269 61881 13280 61927
rect 13108 61823 13280 61881
rect 13108 61777 13119 61823
rect 13165 61777 13223 61823
rect 13269 61777 13280 61823
rect 13108 61719 13280 61777
rect 13108 61673 13119 61719
rect 13165 61673 13223 61719
rect 13269 61673 13280 61719
rect 13108 61615 13280 61673
rect 13108 61569 13119 61615
rect 13165 61569 13223 61615
rect 13269 61569 13280 61615
rect 13108 61511 13280 61569
rect 13108 61465 13119 61511
rect 13165 61465 13223 61511
rect 13269 61465 13280 61511
rect 13108 61407 13280 61465
rect 13108 61361 13119 61407
rect 13165 61361 13223 61407
rect 13269 61361 13280 61407
rect 13108 61303 13280 61361
rect 13108 61257 13119 61303
rect 13165 61257 13223 61303
rect 13269 61257 13280 61303
rect 13108 61199 13280 61257
rect 13108 61153 13119 61199
rect 13165 61153 13223 61199
rect 13269 61153 13280 61199
rect 13108 61095 13280 61153
rect 13108 61049 13119 61095
rect 13165 61049 13223 61095
rect 13269 61049 13280 61095
rect 13108 60991 13280 61049
rect 13108 60945 13119 60991
rect 13165 60945 13223 60991
rect 13269 60945 13280 60991
rect 13108 60887 13280 60945
rect 13108 60841 13119 60887
rect 13165 60841 13223 60887
rect 13269 60841 13280 60887
rect 13108 60783 13280 60841
rect 13108 60737 13119 60783
rect 13165 60737 13223 60783
rect 13269 60737 13280 60783
rect 13108 60679 13280 60737
rect 13108 60633 13119 60679
rect 13165 60633 13223 60679
rect 13269 60633 13280 60679
rect 13108 60575 13280 60633
rect 13108 60529 13119 60575
rect 13165 60529 13223 60575
rect 13269 60529 13280 60575
rect 13108 60471 13280 60529
rect 13108 60425 13119 60471
rect 13165 60425 13223 60471
rect 13269 60425 13280 60471
rect 13108 60367 13280 60425
rect 13108 60321 13119 60367
rect 13165 60321 13223 60367
rect 13269 60321 13280 60367
rect 13108 60263 13280 60321
rect 13108 60217 13119 60263
rect 13165 60217 13223 60263
rect 13269 60217 13280 60263
rect 13108 60159 13280 60217
rect 13108 60113 13119 60159
rect 13165 60113 13223 60159
rect 13269 60113 13280 60159
rect 13108 60055 13280 60113
rect 13108 60009 13119 60055
rect 13165 60009 13223 60055
rect 13269 60009 13280 60055
rect 13108 59951 13280 60009
rect 13108 59905 13119 59951
rect 13165 59905 13223 59951
rect 13269 59905 13280 59951
rect 13108 59847 13280 59905
rect 13108 59801 13119 59847
rect 13165 59801 13223 59847
rect 13269 59801 13280 59847
rect 13108 59743 13280 59801
rect 13108 59697 13119 59743
rect 13165 59697 13223 59743
rect 13269 59697 13280 59743
rect 13108 59639 13280 59697
rect 13108 59593 13119 59639
rect 13165 59593 13223 59639
rect 13269 59593 13280 59639
rect 13108 59535 13280 59593
rect 13108 59489 13119 59535
rect 13165 59489 13223 59535
rect 13269 59489 13280 59535
rect 13108 59431 13280 59489
rect 13108 59385 13119 59431
rect 13165 59385 13223 59431
rect 13269 59385 13280 59431
rect 13108 59327 13280 59385
rect 13108 59281 13119 59327
rect 13165 59281 13223 59327
rect 13269 59281 13280 59327
rect 13108 59223 13280 59281
rect 13108 59177 13119 59223
rect 13165 59177 13223 59223
rect 13269 59177 13280 59223
rect 13108 59119 13280 59177
rect 13108 59073 13119 59119
rect 13165 59073 13223 59119
rect 13269 59073 13280 59119
rect 13108 59015 13280 59073
rect 13108 58969 13119 59015
rect 13165 58969 13223 59015
rect 13269 58969 13280 59015
rect 13108 58911 13280 58969
rect 13108 58865 13119 58911
rect 13165 58865 13223 58911
rect 13269 58865 13280 58911
rect 13108 58807 13280 58865
rect 13108 58761 13119 58807
rect 13165 58761 13223 58807
rect 13269 58761 13280 58807
rect 13108 58703 13280 58761
rect 13108 58657 13119 58703
rect 13165 58657 13223 58703
rect 13269 58657 13280 58703
rect 13108 58599 13280 58657
rect 13108 58553 13119 58599
rect 13165 58553 13223 58599
rect 13269 58553 13280 58599
rect 13108 58495 13280 58553
rect 13108 58449 13119 58495
rect 13165 58449 13223 58495
rect 13269 58449 13280 58495
rect 13108 58391 13280 58449
rect 13108 58345 13119 58391
rect 13165 58345 13223 58391
rect 13269 58345 13280 58391
rect 13108 58287 13280 58345
rect 13108 58241 13119 58287
rect 13165 58241 13223 58287
rect 13269 58241 13280 58287
rect 13108 58183 13280 58241
rect 13108 58137 13119 58183
rect 13165 58137 13223 58183
rect 13269 58137 13280 58183
rect 13108 58079 13280 58137
rect 13108 58033 13119 58079
rect 13165 58033 13223 58079
rect 13269 58033 13280 58079
rect 13108 57975 13280 58033
rect 13108 57929 13119 57975
rect 13165 57929 13223 57975
rect 13269 57929 13280 57975
rect 13108 57871 13280 57929
rect 13108 57825 13119 57871
rect 13165 57825 13223 57871
rect 13269 57825 13280 57871
rect 13108 57767 13280 57825
rect 13108 57721 13119 57767
rect 13165 57721 13223 57767
rect 13269 57721 13280 57767
rect 13108 57663 13280 57721
rect 13108 57617 13119 57663
rect 13165 57617 13223 57663
rect 13269 57617 13280 57663
rect 13108 57559 13280 57617
rect 13108 57513 13119 57559
rect 13165 57513 13223 57559
rect 13269 57513 13280 57559
rect 13108 57455 13280 57513
rect 13108 57409 13119 57455
rect 13165 57409 13223 57455
rect 13269 57409 13280 57455
rect 13108 57351 13280 57409
rect 13108 57305 13119 57351
rect 13165 57305 13223 57351
rect 13269 57305 13280 57351
rect 13108 57247 13280 57305
rect 13108 57201 13119 57247
rect 13165 57201 13223 57247
rect 13269 57201 13280 57247
rect 13108 57143 13280 57201
rect 13108 57097 13119 57143
rect 13165 57097 13223 57143
rect 13269 57097 13280 57143
rect 13108 57039 13280 57097
rect 13108 56993 13119 57039
rect 13165 56993 13223 57039
rect 13269 56993 13280 57039
rect 13108 56935 13280 56993
rect 13108 56889 13119 56935
rect 13165 56889 13223 56935
rect 13269 56889 13280 56935
rect 13108 56831 13280 56889
rect 13108 56785 13119 56831
rect 13165 56785 13223 56831
rect 13269 56785 13280 56831
rect 13108 56727 13280 56785
rect 13108 56681 13119 56727
rect 13165 56681 13223 56727
rect 13269 56681 13280 56727
rect 13108 56623 13280 56681
rect 13108 56577 13119 56623
rect 13165 56577 13223 56623
rect 13269 56577 13280 56623
rect 13108 56519 13280 56577
rect 13108 56473 13119 56519
rect 13165 56473 13223 56519
rect 13269 56473 13280 56519
rect 13108 56415 13280 56473
rect 13108 56369 13119 56415
rect 13165 56369 13223 56415
rect 13269 56369 13280 56415
rect 13108 56311 13280 56369
rect 13108 56265 13119 56311
rect 13165 56265 13223 56311
rect 13269 56265 13280 56311
rect 13108 56207 13280 56265
rect 13108 56161 13119 56207
rect 13165 56161 13223 56207
rect 13269 56161 13280 56207
rect 13108 56103 13280 56161
rect 13108 56057 13119 56103
rect 13165 56057 13223 56103
rect 13269 56057 13280 56103
rect 13108 55999 13280 56057
rect 13108 55953 13119 55999
rect 13165 55953 13223 55999
rect 13269 55953 13280 55999
rect 13108 55895 13280 55953
rect 13108 55849 13119 55895
rect 13165 55849 13223 55895
rect 13269 55849 13280 55895
rect 13108 55791 13280 55849
rect 13108 55745 13119 55791
rect 13165 55745 13223 55791
rect 13269 55745 13280 55791
rect 13108 55687 13280 55745
rect 13108 55641 13119 55687
rect 13165 55641 13223 55687
rect 13269 55641 13280 55687
rect 13108 55583 13280 55641
rect 13108 55537 13119 55583
rect 13165 55537 13223 55583
rect 13269 55537 13280 55583
rect 13108 55479 13280 55537
rect 13108 55433 13119 55479
rect 13165 55433 13223 55479
rect 13269 55433 13280 55479
rect 13108 55375 13280 55433
rect 13108 55329 13119 55375
rect 13165 55329 13223 55375
rect 13269 55329 13280 55375
rect 13108 55271 13280 55329
rect 13108 55225 13119 55271
rect 13165 55225 13223 55271
rect 13269 55225 13280 55271
rect 13108 55167 13280 55225
rect 13108 55121 13119 55167
rect 13165 55121 13223 55167
rect 13269 55121 13280 55167
rect 13108 55063 13280 55121
rect 13108 55017 13119 55063
rect 13165 55017 13223 55063
rect 13269 55017 13280 55063
rect 13108 54959 13280 55017
rect 13108 54913 13119 54959
rect 13165 54913 13223 54959
rect 13269 54913 13280 54959
rect 13108 54855 13280 54913
rect 13108 54809 13119 54855
rect 13165 54809 13223 54855
rect 13269 54809 13280 54855
rect 13108 54751 13280 54809
rect 13108 54705 13119 54751
rect 13165 54705 13223 54751
rect 13269 54705 13280 54751
rect 13108 54647 13280 54705
rect 13108 54601 13119 54647
rect 13165 54601 13223 54647
rect 13269 54601 13280 54647
rect 13108 54543 13280 54601
rect 13108 54497 13119 54543
rect 13165 54497 13223 54543
rect 13269 54497 13280 54543
rect 13108 54439 13280 54497
rect 13108 54393 13119 54439
rect 13165 54393 13223 54439
rect 13269 54393 13280 54439
rect 13108 54335 13280 54393
rect 13108 54289 13119 54335
rect 13165 54289 13223 54335
rect 13269 54289 13280 54335
rect 13108 54231 13280 54289
rect 13108 54185 13119 54231
rect 13165 54185 13223 54231
rect 13269 54185 13280 54231
rect 13108 54127 13280 54185
rect 13108 54081 13119 54127
rect 13165 54081 13223 54127
rect 13269 54081 13280 54127
rect 13108 54023 13280 54081
rect 13108 53977 13119 54023
rect 13165 53977 13223 54023
rect 13269 53977 13280 54023
rect 13108 53919 13280 53977
rect 13108 53873 13119 53919
rect 13165 53873 13223 53919
rect 13269 53873 13280 53919
rect 13108 53815 13280 53873
rect 13108 53769 13119 53815
rect 13165 53769 13223 53815
rect 13269 53769 13280 53815
rect 13108 53711 13280 53769
rect 13108 53665 13119 53711
rect 13165 53665 13223 53711
rect 13269 53665 13280 53711
rect 13108 53607 13280 53665
rect 13108 53561 13119 53607
rect 13165 53561 13223 53607
rect 13269 53561 13280 53607
rect 13108 53503 13280 53561
rect 13108 53457 13119 53503
rect 13165 53457 13223 53503
rect 13269 53457 13280 53503
rect 13108 53399 13280 53457
rect 13108 53353 13119 53399
rect 13165 53353 13223 53399
rect 13269 53353 13280 53399
rect 13108 53295 13280 53353
rect 13108 53249 13119 53295
rect 13165 53249 13223 53295
rect 13269 53249 13280 53295
rect 13108 53191 13280 53249
rect 13108 53145 13119 53191
rect 13165 53145 13223 53191
rect 13269 53145 13280 53191
rect 13108 53087 13280 53145
rect 13108 53041 13119 53087
rect 13165 53041 13223 53087
rect 13269 53041 13280 53087
rect 13108 52983 13280 53041
rect 13108 52937 13119 52983
rect 13165 52937 13223 52983
rect 13269 52937 13280 52983
rect 13108 52879 13280 52937
rect 13108 52833 13119 52879
rect 13165 52833 13223 52879
rect 13269 52833 13280 52879
rect 13108 52775 13280 52833
rect 13108 52729 13119 52775
rect 13165 52729 13223 52775
rect 13269 52729 13280 52775
rect 13108 52671 13280 52729
rect 13108 52625 13119 52671
rect 13165 52625 13223 52671
rect 13269 52625 13280 52671
rect 13108 52567 13280 52625
rect 13108 52521 13119 52567
rect 13165 52521 13223 52567
rect 13269 52521 13280 52567
rect 13108 52463 13280 52521
rect 13108 52417 13119 52463
rect 13165 52417 13223 52463
rect 13269 52417 13280 52463
rect 13108 52359 13280 52417
rect 13108 52313 13119 52359
rect 13165 52313 13223 52359
rect 13269 52313 13280 52359
rect 13108 52255 13280 52313
rect 13108 52209 13119 52255
rect 13165 52209 13223 52255
rect 13269 52209 13280 52255
rect 13108 52151 13280 52209
rect 13108 52105 13119 52151
rect 13165 52105 13223 52151
rect 13269 52105 13280 52151
rect 13108 52047 13280 52105
rect 13108 52001 13119 52047
rect 13165 52001 13223 52047
rect 13269 52001 13280 52047
rect 13108 51943 13280 52001
rect 13108 51897 13119 51943
rect 13165 51897 13223 51943
rect 13269 51897 13280 51943
rect 13108 51839 13280 51897
rect 13108 51793 13119 51839
rect 13165 51793 13223 51839
rect 13269 51793 13280 51839
rect 13108 51735 13280 51793
rect 13108 51689 13119 51735
rect 13165 51689 13223 51735
rect 13269 51689 13280 51735
rect 13108 51631 13280 51689
rect 13108 51585 13119 51631
rect 13165 51585 13223 51631
rect 13269 51585 13280 51631
rect 13108 51527 13280 51585
rect 13108 51481 13119 51527
rect 13165 51481 13223 51527
rect 13269 51481 13280 51527
rect 13108 51423 13280 51481
rect 13108 51377 13119 51423
rect 13165 51377 13223 51423
rect 13269 51377 13280 51423
rect 13108 51319 13280 51377
rect 13108 51273 13119 51319
rect 13165 51273 13223 51319
rect 13269 51273 13280 51319
rect 13108 51215 13280 51273
rect 13108 51169 13119 51215
rect 13165 51169 13223 51215
rect 13269 51169 13280 51215
rect 13108 51111 13280 51169
rect 13108 51065 13119 51111
rect 13165 51065 13223 51111
rect 13269 51065 13280 51111
rect 13108 51007 13280 51065
rect 13108 50961 13119 51007
rect 13165 50961 13223 51007
rect 13269 50961 13280 51007
rect 13108 50903 13280 50961
rect 13108 50857 13119 50903
rect 13165 50857 13223 50903
rect 13269 50857 13280 50903
rect 13108 50799 13280 50857
rect 13108 50753 13119 50799
rect 13165 50753 13223 50799
rect 13269 50753 13280 50799
rect 13108 50695 13280 50753
rect 13108 50649 13119 50695
rect 13165 50649 13223 50695
rect 13269 50649 13280 50695
rect 13108 50591 13280 50649
rect 13108 50545 13119 50591
rect 13165 50545 13223 50591
rect 13269 50545 13280 50591
rect 13108 50487 13280 50545
rect 13108 50441 13119 50487
rect 13165 50441 13223 50487
rect 13269 50441 13280 50487
rect 13108 50383 13280 50441
rect 13108 50337 13119 50383
rect 13165 50337 13223 50383
rect 13269 50337 13280 50383
rect 13108 50279 13280 50337
rect 13108 50233 13119 50279
rect 13165 50233 13223 50279
rect 13269 50233 13280 50279
rect 13108 50175 13280 50233
rect 13108 50129 13119 50175
rect 13165 50129 13223 50175
rect 13269 50129 13280 50175
rect 13108 50071 13280 50129
rect 13108 50025 13119 50071
rect 13165 50025 13223 50071
rect 13269 50025 13280 50071
rect 13108 49967 13280 50025
rect 13108 49921 13119 49967
rect 13165 49921 13223 49967
rect 13269 49921 13280 49967
rect 13108 49863 13280 49921
rect 13108 49817 13119 49863
rect 13165 49817 13223 49863
rect 13269 49817 13280 49863
rect 13108 49759 13280 49817
rect 13108 49713 13119 49759
rect 13165 49713 13223 49759
rect 13269 49713 13280 49759
rect 13108 49655 13280 49713
rect 13108 49609 13119 49655
rect 13165 49609 13223 49655
rect 13269 49609 13280 49655
rect 13108 49551 13280 49609
rect 13108 49505 13119 49551
rect 13165 49505 13223 49551
rect 13269 49505 13280 49551
rect 13108 49447 13280 49505
rect 13108 49401 13119 49447
rect 13165 49401 13223 49447
rect 13269 49401 13280 49447
rect 13108 49343 13280 49401
rect 13108 49297 13119 49343
rect 13165 49297 13223 49343
rect 13269 49297 13280 49343
rect 13108 49239 13280 49297
rect 13108 49193 13119 49239
rect 13165 49193 13223 49239
rect 13269 49193 13280 49239
rect 13108 49135 13280 49193
rect 13108 49089 13119 49135
rect 13165 49089 13223 49135
rect 13269 49089 13280 49135
rect 13108 49031 13280 49089
rect 13108 48985 13119 49031
rect 13165 48985 13223 49031
rect 13269 48985 13280 49031
rect 13108 48927 13280 48985
rect 13108 48881 13119 48927
rect 13165 48881 13223 48927
rect 13269 48881 13280 48927
rect 13108 48823 13280 48881
rect 13108 48777 13119 48823
rect 13165 48777 13223 48823
rect 13269 48777 13280 48823
rect 13108 48719 13280 48777
rect 13108 48673 13119 48719
rect 13165 48673 13223 48719
rect 13269 48673 13280 48719
rect 13108 48615 13280 48673
rect 13108 48569 13119 48615
rect 13165 48569 13223 48615
rect 13269 48569 13280 48615
rect 13108 48511 13280 48569
rect 13108 48465 13119 48511
rect 13165 48465 13223 48511
rect 13269 48465 13280 48511
rect 13108 48407 13280 48465
rect 13108 48361 13119 48407
rect 13165 48361 13223 48407
rect 13269 48361 13280 48407
rect 13108 48303 13280 48361
rect 13108 48257 13119 48303
rect 13165 48257 13223 48303
rect 13269 48257 13280 48303
rect 13108 48199 13280 48257
rect 13108 48153 13119 48199
rect 13165 48153 13223 48199
rect 13269 48153 13280 48199
rect 13108 48095 13280 48153
rect 13108 48049 13119 48095
rect 13165 48049 13223 48095
rect 13269 48049 13280 48095
rect 13108 47991 13280 48049
rect 13108 47945 13119 47991
rect 13165 47945 13223 47991
rect 13269 47945 13280 47991
rect 13108 47887 13280 47945
rect 13108 47841 13119 47887
rect 13165 47841 13223 47887
rect 13269 47841 13280 47887
rect 13108 47783 13280 47841
rect 13108 47737 13119 47783
rect 13165 47737 13223 47783
rect 13269 47737 13280 47783
rect 13108 47679 13280 47737
rect 13108 47633 13119 47679
rect 13165 47633 13223 47679
rect 13269 47633 13280 47679
rect 13108 47575 13280 47633
rect 13108 47529 13119 47575
rect 13165 47529 13223 47575
rect 13269 47529 13280 47575
rect 13108 47471 13280 47529
rect 13108 47425 13119 47471
rect 13165 47425 13223 47471
rect 13269 47425 13280 47471
rect 13108 47367 13280 47425
rect 13108 47321 13119 47367
rect 13165 47321 13223 47367
rect 13269 47321 13280 47367
rect 13108 47263 13280 47321
rect 13108 47217 13119 47263
rect 13165 47217 13223 47263
rect 13269 47217 13280 47263
rect 13108 47159 13280 47217
rect 13108 47113 13119 47159
rect 13165 47113 13223 47159
rect 13269 47113 13280 47159
rect 13108 47055 13280 47113
rect 13108 47009 13119 47055
rect 13165 47009 13223 47055
rect 13269 47009 13280 47055
rect 13108 46951 13280 47009
rect 13108 46905 13119 46951
rect 13165 46905 13223 46951
rect 13269 46905 13280 46951
rect 13108 46847 13280 46905
rect 13108 46801 13119 46847
rect 13165 46801 13223 46847
rect 13269 46801 13280 46847
rect 13108 46743 13280 46801
rect 13108 46697 13119 46743
rect 13165 46697 13223 46743
rect 13269 46697 13280 46743
rect 13108 46639 13280 46697
rect 13108 46593 13119 46639
rect 13165 46593 13223 46639
rect 13269 46593 13280 46639
rect 13108 46535 13280 46593
rect 13108 46489 13119 46535
rect 13165 46489 13223 46535
rect 13269 46489 13280 46535
rect 13108 46431 13280 46489
rect 13108 46385 13119 46431
rect 13165 46385 13223 46431
rect 13269 46385 13280 46431
rect 13108 46327 13280 46385
rect 13108 46281 13119 46327
rect 13165 46281 13223 46327
rect 13269 46281 13280 46327
rect 13108 46223 13280 46281
rect 13108 46177 13119 46223
rect 13165 46177 13223 46223
rect 13269 46177 13280 46223
rect 13108 46119 13280 46177
rect 13108 46073 13119 46119
rect 13165 46073 13223 46119
rect 13269 46073 13280 46119
rect 13108 46015 13280 46073
rect 13108 45969 13119 46015
rect 13165 45969 13223 46015
rect 13269 45969 13280 46015
rect 13108 45911 13280 45969
rect 13108 45865 13119 45911
rect 13165 45865 13223 45911
rect 13269 45865 13280 45911
rect 13108 45807 13280 45865
rect 13108 45761 13119 45807
rect 13165 45761 13223 45807
rect 13269 45761 13280 45807
rect 13108 45703 13280 45761
rect 13108 45657 13119 45703
rect 13165 45657 13223 45703
rect 13269 45657 13280 45703
rect 13108 45599 13280 45657
rect 13108 45553 13119 45599
rect 13165 45553 13223 45599
rect 13269 45553 13280 45599
rect 13108 45495 13280 45553
rect 13108 45449 13119 45495
rect 13165 45449 13223 45495
rect 13269 45449 13280 45495
rect 13108 45391 13280 45449
rect 13108 45345 13119 45391
rect 13165 45345 13223 45391
rect 13269 45345 13280 45391
rect 13108 45287 13280 45345
rect 13108 45241 13119 45287
rect 13165 45241 13223 45287
rect 13269 45241 13280 45287
rect 13108 45183 13280 45241
rect 13108 45137 13119 45183
rect 13165 45137 13223 45183
rect 13269 45137 13280 45183
rect 13108 45079 13280 45137
rect 13108 45033 13119 45079
rect 13165 45033 13223 45079
rect 13269 45033 13280 45079
rect 13108 44848 13280 45033
rect 70813 69758 70824 69785
rect 70870 69758 70928 69804
rect 70974 69758 71000 69804
rect 70813 69700 71000 69758
rect 70813 69654 70824 69700
rect 70870 69654 70928 69700
rect 70974 69654 71000 69700
rect 70813 69596 71000 69654
rect 70813 69550 70824 69596
rect 70870 69550 70928 69596
rect 70974 69550 71000 69596
rect 70813 69492 71000 69550
rect 70813 69446 70824 69492
rect 70870 69446 70928 69492
rect 70974 69446 71000 69492
rect 70813 69388 71000 69446
rect 70813 69342 70824 69388
rect 70870 69342 70928 69388
rect 70974 69342 71000 69388
rect 70813 69284 71000 69342
rect 70813 69238 70824 69284
rect 70870 69238 70928 69284
rect 70974 69238 71000 69284
rect 70813 69180 71000 69238
rect 70813 69134 70824 69180
rect 70870 69134 70928 69180
rect 70974 69134 71000 69180
rect 70813 69076 71000 69134
rect 70813 69030 70824 69076
rect 70870 69030 70928 69076
rect 70974 69030 71000 69076
rect 70813 68972 71000 69030
rect 70813 68926 70824 68972
rect 70870 68926 70928 68972
rect 70974 68926 71000 68972
rect 70813 68868 71000 68926
rect 70813 68822 70824 68868
rect 70870 68822 70928 68868
rect 70974 68822 71000 68868
rect 70813 68764 71000 68822
rect 70813 68718 70824 68764
rect 70870 68718 70928 68764
rect 70974 68718 71000 68764
rect 70813 68660 71000 68718
rect 70813 68614 70824 68660
rect 70870 68614 70928 68660
rect 70974 68614 71000 68660
rect 70813 68556 71000 68614
rect 70813 68510 70824 68556
rect 70870 68510 70928 68556
rect 70974 68510 71000 68556
rect 70813 68452 71000 68510
rect 70813 68406 70824 68452
rect 70870 68406 70928 68452
rect 70974 68406 71000 68452
rect 70813 68348 71000 68406
rect 70813 68302 70824 68348
rect 70870 68302 70928 68348
rect 70974 68302 71000 68348
rect 70813 68244 71000 68302
rect 70813 68198 70824 68244
rect 70870 68198 70928 68244
rect 70974 68198 71000 68244
rect 70813 68140 71000 68198
rect 70813 68094 70824 68140
rect 70870 68094 70928 68140
rect 70974 68094 71000 68140
rect 70813 68036 71000 68094
rect 70813 67990 70824 68036
rect 70870 67990 70928 68036
rect 70974 67990 71000 68036
rect 70813 67932 71000 67990
rect 70813 67886 70824 67932
rect 70870 67886 70928 67932
rect 70974 67886 71000 67932
rect 70813 67828 71000 67886
rect 70813 67782 70824 67828
rect 70870 67782 70928 67828
rect 70974 67782 71000 67828
rect 70813 67724 71000 67782
rect 70813 67678 70824 67724
rect 70870 67678 70928 67724
rect 70974 67678 71000 67724
rect 70813 67620 71000 67678
rect 70813 67574 70824 67620
rect 70870 67574 70928 67620
rect 70974 67574 71000 67620
rect 70813 67516 71000 67574
rect 70813 67470 70824 67516
rect 70870 67470 70928 67516
rect 70974 67470 71000 67516
rect 70813 67412 71000 67470
rect 70813 67366 70824 67412
rect 70870 67366 70928 67412
rect 70974 67366 71000 67412
rect 70813 67308 71000 67366
rect 70813 67262 70824 67308
rect 70870 67262 70928 67308
rect 70974 67262 71000 67308
rect 70813 67204 71000 67262
rect 70813 67158 70824 67204
rect 70870 67158 70928 67204
rect 70974 67158 71000 67204
rect 70813 67100 71000 67158
rect 70813 67054 70824 67100
rect 70870 67054 70928 67100
rect 70974 67054 71000 67100
rect 70813 66996 71000 67054
rect 70813 66950 70824 66996
rect 70870 66950 70928 66996
rect 70974 66950 71000 66996
rect 70813 66892 71000 66950
rect 70813 66846 70824 66892
rect 70870 66846 70928 66892
rect 70974 66846 71000 66892
rect 70813 66788 71000 66846
rect 70813 66742 70824 66788
rect 70870 66742 70928 66788
rect 70974 66742 71000 66788
rect 70813 66684 71000 66742
rect 70813 66638 70824 66684
rect 70870 66638 70928 66684
rect 70974 66638 71000 66684
rect 70813 66580 71000 66638
rect 70813 66534 70824 66580
rect 70870 66534 70928 66580
rect 70974 66534 71000 66580
rect 70813 66476 71000 66534
rect 70813 66430 70824 66476
rect 70870 66430 70928 66476
rect 70974 66430 71000 66476
rect 70813 66372 71000 66430
rect 70813 66326 70824 66372
rect 70870 66326 70928 66372
rect 70974 66326 71000 66372
rect 70813 66268 71000 66326
rect 70813 66222 70824 66268
rect 70870 66222 70928 66268
rect 70974 66222 71000 66268
rect 70813 66164 71000 66222
rect 70813 66118 70824 66164
rect 70870 66118 70928 66164
rect 70974 66118 71000 66164
rect 70813 66060 71000 66118
rect 70813 66014 70824 66060
rect 70870 66014 70928 66060
rect 70974 66014 71000 66060
rect 70813 65956 71000 66014
rect 70813 65910 70824 65956
rect 70870 65910 70928 65956
rect 70974 65910 71000 65956
rect 70813 65852 71000 65910
rect 70813 65806 70824 65852
rect 70870 65806 70928 65852
rect 70974 65806 71000 65852
rect 70813 65748 71000 65806
rect 70813 65702 70824 65748
rect 70870 65702 70928 65748
rect 70974 65702 71000 65748
rect 70813 65644 71000 65702
rect 70813 65598 70824 65644
rect 70870 65598 70928 65644
rect 70974 65598 71000 65644
rect 70813 65540 71000 65598
rect 70813 65494 70824 65540
rect 70870 65494 70928 65540
rect 70974 65494 71000 65540
rect 70813 65436 71000 65494
rect 70813 65390 70824 65436
rect 70870 65390 70928 65436
rect 70974 65390 71000 65436
rect 70813 65332 71000 65390
rect 70813 65286 70824 65332
rect 70870 65286 70928 65332
rect 70974 65286 71000 65332
rect 70813 65228 71000 65286
rect 70813 65182 70824 65228
rect 70870 65182 70928 65228
rect 70974 65182 71000 65228
rect 70813 65124 71000 65182
rect 70813 65078 70824 65124
rect 70870 65078 70928 65124
rect 70974 65078 71000 65124
rect 70813 65020 71000 65078
rect 70813 64974 70824 65020
rect 70870 64974 70928 65020
rect 70974 64974 71000 65020
rect 70813 64916 71000 64974
rect 70813 64870 70824 64916
rect 70870 64870 70928 64916
rect 70974 64870 71000 64916
rect 70813 64812 71000 64870
rect 70813 64766 70824 64812
rect 70870 64766 70928 64812
rect 70974 64766 71000 64812
rect 70813 64708 71000 64766
rect 70813 64662 70824 64708
rect 70870 64662 70928 64708
rect 70974 64662 71000 64708
rect 70813 64604 71000 64662
rect 70813 64558 70824 64604
rect 70870 64558 70928 64604
rect 70974 64558 71000 64604
rect 70813 64500 71000 64558
rect 70813 64454 70824 64500
rect 70870 64454 70928 64500
rect 70974 64454 71000 64500
rect 70813 64396 71000 64454
rect 70813 64350 70824 64396
rect 70870 64350 70928 64396
rect 70974 64350 71000 64396
rect 70813 64292 71000 64350
rect 70813 64246 70824 64292
rect 70870 64246 70928 64292
rect 70974 64246 71000 64292
rect 70813 64188 71000 64246
rect 70813 64142 70824 64188
rect 70870 64142 70928 64188
rect 70974 64142 71000 64188
rect 70813 64084 71000 64142
rect 70813 64038 70824 64084
rect 70870 64038 70928 64084
rect 70974 64038 71000 64084
rect 70813 63980 71000 64038
rect 70813 63934 70824 63980
rect 70870 63934 70928 63980
rect 70974 63934 71000 63980
rect 70813 63876 71000 63934
rect 70813 63830 70824 63876
rect 70870 63830 70928 63876
rect 70974 63830 71000 63876
rect 70813 63772 71000 63830
rect 70813 63726 70824 63772
rect 70870 63726 70928 63772
rect 70974 63726 71000 63772
rect 70813 63668 71000 63726
rect 70813 63622 70824 63668
rect 70870 63622 70928 63668
rect 70974 63622 71000 63668
rect 70813 63564 71000 63622
rect 70813 63518 70824 63564
rect 70870 63518 70928 63564
rect 70974 63518 71000 63564
rect 70813 63460 71000 63518
rect 70813 63414 70824 63460
rect 70870 63414 70928 63460
rect 70974 63414 71000 63460
rect 70813 63356 71000 63414
rect 70813 63310 70824 63356
rect 70870 63310 70928 63356
rect 70974 63310 71000 63356
rect 70813 63252 71000 63310
rect 70813 63206 70824 63252
rect 70870 63206 70928 63252
rect 70974 63206 71000 63252
rect 70813 63148 71000 63206
rect 70813 63102 70824 63148
rect 70870 63102 70928 63148
rect 70974 63102 71000 63148
rect 70813 63044 71000 63102
rect 70813 62998 70824 63044
rect 70870 62998 70928 63044
rect 70974 62998 71000 63044
rect 70813 62940 71000 62998
rect 70813 62894 70824 62940
rect 70870 62894 70928 62940
rect 70974 62894 71000 62940
rect 70813 62836 71000 62894
rect 70813 62790 70824 62836
rect 70870 62790 70928 62836
rect 70974 62790 71000 62836
rect 70813 62732 71000 62790
rect 70813 62686 70824 62732
rect 70870 62686 70928 62732
rect 70974 62686 71000 62732
rect 70813 62628 71000 62686
rect 70813 62582 70824 62628
rect 70870 62582 70928 62628
rect 70974 62582 71000 62628
rect 70813 62524 71000 62582
rect 70813 62478 70824 62524
rect 70870 62478 70928 62524
rect 70974 62478 71000 62524
rect 70813 62420 71000 62478
rect 70813 62374 70824 62420
rect 70870 62374 70928 62420
rect 70974 62374 71000 62420
rect 70813 62316 71000 62374
rect 70813 62270 70824 62316
rect 70870 62270 70928 62316
rect 70974 62270 71000 62316
rect 70813 62212 71000 62270
rect 70813 62166 70824 62212
rect 70870 62166 70928 62212
rect 70974 62166 71000 62212
rect 70813 62108 71000 62166
rect 70813 62062 70824 62108
rect 70870 62062 70928 62108
rect 70974 62062 71000 62108
rect 70813 62004 71000 62062
rect 70813 61958 70824 62004
rect 70870 61958 70928 62004
rect 70974 61958 71000 62004
rect 70813 61900 71000 61958
rect 70813 61854 70824 61900
rect 70870 61854 70928 61900
rect 70974 61854 71000 61900
rect 70813 61796 71000 61854
rect 70813 61750 70824 61796
rect 70870 61750 70928 61796
rect 70974 61750 71000 61796
rect 70813 61692 71000 61750
rect 70813 61646 70824 61692
rect 70870 61646 70928 61692
rect 70974 61646 71000 61692
rect 70813 61588 71000 61646
rect 70813 61542 70824 61588
rect 70870 61542 70928 61588
rect 70974 61542 71000 61588
rect 70813 61484 71000 61542
rect 70813 61438 70824 61484
rect 70870 61438 70928 61484
rect 70974 61438 71000 61484
rect 70813 61380 71000 61438
rect 70813 61334 70824 61380
rect 70870 61334 70928 61380
rect 70974 61334 71000 61380
rect 70813 61276 71000 61334
rect 70813 61230 70824 61276
rect 70870 61230 70928 61276
rect 70974 61230 71000 61276
rect 70813 61172 71000 61230
rect 70813 61126 70824 61172
rect 70870 61126 70928 61172
rect 70974 61126 71000 61172
rect 70813 61068 71000 61126
rect 70813 61022 70824 61068
rect 70870 61022 70928 61068
rect 70974 61022 71000 61068
rect 70813 60964 71000 61022
rect 70813 60918 70824 60964
rect 70870 60918 70928 60964
rect 70974 60918 71000 60964
rect 70813 60860 71000 60918
rect 70813 60814 70824 60860
rect 70870 60814 70928 60860
rect 70974 60814 71000 60860
rect 70813 60756 71000 60814
rect 70813 60710 70824 60756
rect 70870 60710 70928 60756
rect 70974 60710 71000 60756
rect 70813 60652 71000 60710
rect 70813 60606 70824 60652
rect 70870 60606 70928 60652
rect 70974 60606 71000 60652
rect 70813 60548 71000 60606
rect 70813 60502 70824 60548
rect 70870 60502 70928 60548
rect 70974 60502 71000 60548
rect 70813 60444 71000 60502
rect 70813 60398 70824 60444
rect 70870 60398 70928 60444
rect 70974 60398 71000 60444
rect 70813 60340 71000 60398
rect 70813 60294 70824 60340
rect 70870 60294 70928 60340
rect 70974 60294 71000 60340
rect 70813 60236 71000 60294
rect 70813 60190 70824 60236
rect 70870 60190 70928 60236
rect 70974 60190 71000 60236
rect 70813 60132 71000 60190
rect 70813 60086 70824 60132
rect 70870 60086 70928 60132
rect 70974 60086 71000 60132
rect 70813 60028 71000 60086
rect 70813 59982 70824 60028
rect 70870 59982 70928 60028
rect 70974 59982 71000 60028
rect 70813 59924 71000 59982
rect 70813 59878 70824 59924
rect 70870 59878 70928 59924
rect 70974 59878 71000 59924
rect 70813 59820 71000 59878
rect 70813 59774 70824 59820
rect 70870 59774 70928 59820
rect 70974 59774 71000 59820
rect 70813 59716 71000 59774
rect 70813 59670 70824 59716
rect 70870 59670 70928 59716
rect 70974 59670 71000 59716
rect 70813 59612 71000 59670
rect 70813 59566 70824 59612
rect 70870 59566 70928 59612
rect 70974 59566 71000 59612
rect 70813 59508 71000 59566
rect 70813 59462 70824 59508
rect 70870 59462 70928 59508
rect 70974 59462 71000 59508
rect 70813 59404 71000 59462
rect 70813 59358 70824 59404
rect 70870 59358 70928 59404
rect 70974 59358 71000 59404
rect 70813 59300 71000 59358
rect 70813 59254 70824 59300
rect 70870 59254 70928 59300
rect 70974 59254 71000 59300
rect 70813 59196 71000 59254
rect 70813 59150 70824 59196
rect 70870 59150 70928 59196
rect 70974 59150 71000 59196
rect 70813 59092 71000 59150
rect 70813 59046 70824 59092
rect 70870 59046 70928 59092
rect 70974 59046 71000 59092
rect 70813 58988 71000 59046
rect 70813 58942 70824 58988
rect 70870 58942 70928 58988
rect 70974 58942 71000 58988
rect 70813 58884 71000 58942
rect 70813 58838 70824 58884
rect 70870 58838 70928 58884
rect 70974 58838 71000 58884
rect 70813 58780 71000 58838
rect 70813 58734 70824 58780
rect 70870 58734 70928 58780
rect 70974 58734 71000 58780
rect 70813 58676 71000 58734
rect 70813 58630 70824 58676
rect 70870 58630 70928 58676
rect 70974 58630 71000 58676
rect 70813 58572 71000 58630
rect 70813 58526 70824 58572
rect 70870 58526 70928 58572
rect 70974 58526 71000 58572
rect 70813 58468 71000 58526
rect 70813 58422 70824 58468
rect 70870 58422 70928 58468
rect 70974 58422 71000 58468
rect 70813 58364 71000 58422
rect 70813 58318 70824 58364
rect 70870 58318 70928 58364
rect 70974 58318 71000 58364
rect 70813 58260 71000 58318
rect 70813 58214 70824 58260
rect 70870 58214 70928 58260
rect 70974 58214 71000 58260
rect 70813 58156 71000 58214
rect 70813 58110 70824 58156
rect 70870 58110 70928 58156
rect 70974 58110 71000 58156
rect 70813 58052 71000 58110
rect 70813 58006 70824 58052
rect 70870 58006 70928 58052
rect 70974 58006 71000 58052
rect 70813 57948 71000 58006
rect 70813 57902 70824 57948
rect 70870 57902 70928 57948
rect 70974 57902 71000 57948
rect 70813 57844 71000 57902
rect 70813 57798 70824 57844
rect 70870 57798 70928 57844
rect 70974 57798 71000 57844
rect 70813 57740 71000 57798
rect 70813 57694 70824 57740
rect 70870 57694 70928 57740
rect 70974 57694 71000 57740
rect 70813 57636 71000 57694
rect 70813 57590 70824 57636
rect 70870 57590 70928 57636
rect 70974 57590 71000 57636
rect 70813 57532 71000 57590
rect 70813 57486 70824 57532
rect 70870 57486 70928 57532
rect 70974 57486 71000 57532
rect 70813 57428 71000 57486
rect 70813 57382 70824 57428
rect 70870 57382 70928 57428
rect 70974 57382 71000 57428
rect 70813 57324 71000 57382
rect 70813 57278 70824 57324
rect 70870 57278 70928 57324
rect 70974 57278 71000 57324
rect 70813 57220 71000 57278
rect 70813 57174 70824 57220
rect 70870 57174 70928 57220
rect 70974 57174 71000 57220
rect 70813 57116 71000 57174
rect 70813 57070 70824 57116
rect 70870 57070 70928 57116
rect 70974 57070 71000 57116
rect 70813 57012 71000 57070
rect 70813 56966 70824 57012
rect 70870 56966 70928 57012
rect 70974 56966 71000 57012
rect 70813 56908 71000 56966
rect 70813 56862 70824 56908
rect 70870 56862 70928 56908
rect 70974 56862 71000 56908
rect 70813 56804 71000 56862
rect 70813 56758 70824 56804
rect 70870 56758 70928 56804
rect 70974 56758 71000 56804
rect 70813 56700 71000 56758
rect 70813 56654 70824 56700
rect 70870 56654 70928 56700
rect 70974 56654 71000 56700
rect 70813 56596 71000 56654
rect 70813 56550 70824 56596
rect 70870 56550 70928 56596
rect 70974 56550 71000 56596
rect 70813 56492 71000 56550
rect 70813 56446 70824 56492
rect 70870 56446 70928 56492
rect 70974 56446 71000 56492
rect 70813 56388 71000 56446
rect 70813 56342 70824 56388
rect 70870 56342 70928 56388
rect 70974 56342 71000 56388
rect 70813 56284 71000 56342
rect 70813 56238 70824 56284
rect 70870 56238 70928 56284
rect 70974 56238 71000 56284
rect 70813 56180 71000 56238
rect 70813 56134 70824 56180
rect 70870 56134 70928 56180
rect 70974 56134 71000 56180
rect 70813 56076 71000 56134
rect 70813 56030 70824 56076
rect 70870 56030 70928 56076
rect 70974 56030 71000 56076
rect 70813 55972 71000 56030
rect 70813 55926 70824 55972
rect 70870 55926 70928 55972
rect 70974 55926 71000 55972
rect 70813 55868 71000 55926
rect 70813 55822 70824 55868
rect 70870 55822 70928 55868
rect 70974 55822 71000 55868
rect 70813 55764 71000 55822
rect 70813 55718 70824 55764
rect 70870 55718 70928 55764
rect 70974 55718 71000 55764
rect 70813 55660 71000 55718
rect 70813 55614 70824 55660
rect 70870 55614 70928 55660
rect 70974 55614 71000 55660
rect 70813 55556 71000 55614
rect 70813 55510 70824 55556
rect 70870 55510 70928 55556
rect 70974 55510 71000 55556
rect 70813 55452 71000 55510
rect 70813 55406 70824 55452
rect 70870 55406 70928 55452
rect 70974 55406 71000 55452
rect 70813 55348 71000 55406
rect 70813 55302 70824 55348
rect 70870 55302 70928 55348
rect 70974 55302 71000 55348
rect 70813 55244 71000 55302
rect 70813 55198 70824 55244
rect 70870 55198 70928 55244
rect 70974 55198 71000 55244
rect 70813 55140 71000 55198
rect 70813 55094 70824 55140
rect 70870 55094 70928 55140
rect 70974 55094 71000 55140
rect 70813 55036 71000 55094
rect 70813 54990 70824 55036
rect 70870 54990 70928 55036
rect 70974 54990 71000 55036
rect 70813 54932 71000 54990
rect 70813 54886 70824 54932
rect 70870 54886 70928 54932
rect 70974 54886 71000 54932
rect 70813 54828 71000 54886
rect 70813 54782 70824 54828
rect 70870 54782 70928 54828
rect 70974 54782 71000 54828
rect 70813 54724 71000 54782
rect 70813 54678 70824 54724
rect 70870 54678 70928 54724
rect 70974 54678 71000 54724
rect 70813 54620 71000 54678
rect 70813 54574 70824 54620
rect 70870 54574 70928 54620
rect 70974 54574 71000 54620
rect 70813 54516 71000 54574
rect 70813 54470 70824 54516
rect 70870 54470 70928 54516
rect 70974 54470 71000 54516
rect 70813 54412 71000 54470
rect 70813 54366 70824 54412
rect 70870 54366 70928 54412
rect 70974 54366 71000 54412
rect 70813 54308 71000 54366
rect 70813 54262 70824 54308
rect 70870 54262 70928 54308
rect 70974 54262 71000 54308
rect 70813 54204 71000 54262
rect 70813 54158 70824 54204
rect 70870 54158 70928 54204
rect 70974 54158 71000 54204
rect 70813 54100 71000 54158
rect 70813 54054 70824 54100
rect 70870 54054 70928 54100
rect 70974 54054 71000 54100
rect 70813 53996 71000 54054
rect 70813 53950 70824 53996
rect 70870 53950 70928 53996
rect 70974 53950 71000 53996
rect 70813 53892 71000 53950
rect 70813 53846 70824 53892
rect 70870 53846 70928 53892
rect 70974 53846 71000 53892
rect 70813 53788 71000 53846
rect 70813 53742 70824 53788
rect 70870 53742 70928 53788
rect 70974 53742 71000 53788
rect 70813 53684 71000 53742
rect 70813 53638 70824 53684
rect 70870 53638 70928 53684
rect 70974 53638 71000 53684
rect 70813 53580 71000 53638
rect 70813 53534 70824 53580
rect 70870 53534 70928 53580
rect 70974 53534 71000 53580
rect 70813 53476 71000 53534
rect 70813 53430 70824 53476
rect 70870 53430 70928 53476
rect 70974 53430 71000 53476
rect 70813 53372 71000 53430
rect 70813 53326 70824 53372
rect 70870 53326 70928 53372
rect 70974 53326 71000 53372
rect 70813 53268 71000 53326
rect 70813 53222 70824 53268
rect 70870 53222 70928 53268
rect 70974 53222 71000 53268
rect 70813 53164 71000 53222
rect 70813 53118 70824 53164
rect 70870 53118 70928 53164
rect 70974 53118 71000 53164
rect 70813 53060 71000 53118
rect 70813 53014 70824 53060
rect 70870 53014 70928 53060
rect 70974 53014 71000 53060
rect 70813 52956 71000 53014
rect 70813 52910 70824 52956
rect 70870 52910 70928 52956
rect 70974 52910 71000 52956
rect 70813 52852 71000 52910
rect 70813 52806 70824 52852
rect 70870 52806 70928 52852
rect 70974 52806 71000 52852
rect 70813 52748 71000 52806
rect 70813 52702 70824 52748
rect 70870 52702 70928 52748
rect 70974 52702 71000 52748
rect 70813 52644 71000 52702
rect 70813 52598 70824 52644
rect 70870 52598 70928 52644
rect 70974 52598 71000 52644
rect 70813 52540 71000 52598
rect 70813 52494 70824 52540
rect 70870 52494 70928 52540
rect 70974 52494 71000 52540
rect 70813 52436 71000 52494
rect 70813 52390 70824 52436
rect 70870 52390 70928 52436
rect 70974 52390 71000 52436
rect 70813 52332 71000 52390
rect 70813 52286 70824 52332
rect 70870 52286 70928 52332
rect 70974 52286 71000 52332
rect 70813 52228 71000 52286
rect 70813 52182 70824 52228
rect 70870 52182 70928 52228
rect 70974 52182 71000 52228
rect 70813 52124 71000 52182
rect 70813 52078 70824 52124
rect 70870 52078 70928 52124
rect 70974 52078 71000 52124
rect 70813 52020 71000 52078
rect 70813 51974 70824 52020
rect 70870 51974 70928 52020
rect 70974 51974 71000 52020
rect 70813 51916 71000 51974
rect 70813 51870 70824 51916
rect 70870 51870 70928 51916
rect 70974 51870 71000 51916
rect 70813 51812 71000 51870
rect 70813 51766 70824 51812
rect 70870 51766 70928 51812
rect 70974 51766 71000 51812
rect 70813 51708 71000 51766
rect 70813 51662 70824 51708
rect 70870 51662 70928 51708
rect 70974 51662 71000 51708
rect 70813 51604 71000 51662
rect 70813 51558 70824 51604
rect 70870 51558 70928 51604
rect 70974 51558 71000 51604
rect 70813 51500 71000 51558
rect 70813 51454 70824 51500
rect 70870 51454 70928 51500
rect 70974 51454 71000 51500
rect 70813 51396 71000 51454
rect 70813 51350 70824 51396
rect 70870 51350 70928 51396
rect 70974 51350 71000 51396
rect 70813 51292 71000 51350
rect 70813 51246 70824 51292
rect 70870 51246 70928 51292
rect 70974 51246 71000 51292
rect 70813 51188 71000 51246
rect 70813 51142 70824 51188
rect 70870 51142 70928 51188
rect 70974 51142 71000 51188
rect 70813 51084 71000 51142
rect 70813 51038 70824 51084
rect 70870 51038 70928 51084
rect 70974 51038 71000 51084
rect 70813 50980 71000 51038
rect 70813 50934 70824 50980
rect 70870 50934 70928 50980
rect 70974 50934 71000 50980
rect 70813 50876 71000 50934
rect 70813 50830 70824 50876
rect 70870 50830 70928 50876
rect 70974 50830 71000 50876
rect 70813 50772 71000 50830
rect 70813 50726 70824 50772
rect 70870 50726 70928 50772
rect 70974 50726 71000 50772
rect 70813 50668 71000 50726
rect 70813 50622 70824 50668
rect 70870 50622 70928 50668
rect 70974 50622 71000 50668
rect 70813 50564 71000 50622
rect 70813 50518 70824 50564
rect 70870 50518 70928 50564
rect 70974 50518 71000 50564
rect 70813 50460 71000 50518
rect 70813 50414 70824 50460
rect 70870 50414 70928 50460
rect 70974 50414 71000 50460
rect 70813 50356 71000 50414
rect 70813 50310 70824 50356
rect 70870 50310 70928 50356
rect 70974 50310 71000 50356
rect 70813 50252 71000 50310
rect 70813 50206 70824 50252
rect 70870 50206 70928 50252
rect 70974 50206 71000 50252
rect 70813 50148 71000 50206
rect 70813 50102 70824 50148
rect 70870 50102 70928 50148
rect 70974 50102 71000 50148
rect 70813 50044 71000 50102
rect 70813 49998 70824 50044
rect 70870 49998 70928 50044
rect 70974 49998 71000 50044
rect 70813 49940 71000 49998
rect 70813 49894 70824 49940
rect 70870 49894 70928 49940
rect 70974 49894 71000 49940
rect 70813 49836 71000 49894
rect 70813 49790 70824 49836
rect 70870 49790 70928 49836
rect 70974 49790 71000 49836
rect 70813 49732 71000 49790
rect 70813 49686 70824 49732
rect 70870 49686 70928 49732
rect 70974 49686 71000 49732
rect 70813 49628 71000 49686
rect 70813 49582 70824 49628
rect 70870 49582 70928 49628
rect 70974 49582 71000 49628
rect 70813 49524 71000 49582
rect 70813 49478 70824 49524
rect 70870 49478 70928 49524
rect 70974 49478 71000 49524
rect 70813 49420 71000 49478
rect 70813 49374 70824 49420
rect 70870 49374 70928 49420
rect 70974 49374 71000 49420
rect 70813 49316 71000 49374
rect 70813 49270 70824 49316
rect 70870 49270 70928 49316
rect 70974 49270 71000 49316
rect 70813 49212 71000 49270
rect 70813 49166 70824 49212
rect 70870 49166 70928 49212
rect 70974 49166 71000 49212
rect 70813 49108 71000 49166
rect 70813 49062 70824 49108
rect 70870 49062 70928 49108
rect 70974 49062 71000 49108
rect 70813 49004 71000 49062
rect 70813 48958 70824 49004
rect 70870 48958 70928 49004
rect 70974 48958 71000 49004
rect 70813 48900 71000 48958
rect 70813 48854 70824 48900
rect 70870 48854 70928 48900
rect 70974 48854 71000 48900
rect 70813 48796 71000 48854
rect 70813 48750 70824 48796
rect 70870 48750 70928 48796
rect 70974 48750 71000 48796
rect 70813 48692 71000 48750
rect 70813 48646 70824 48692
rect 70870 48646 70928 48692
rect 70974 48646 71000 48692
rect 70813 48588 71000 48646
rect 70813 48542 70824 48588
rect 70870 48542 70928 48588
rect 70974 48542 71000 48588
rect 70813 48484 71000 48542
rect 70813 48438 70824 48484
rect 70870 48438 70928 48484
rect 70974 48438 71000 48484
rect 70813 48380 71000 48438
rect 70813 48334 70824 48380
rect 70870 48334 70928 48380
rect 70974 48334 71000 48380
rect 70813 48276 71000 48334
rect 70813 48230 70824 48276
rect 70870 48230 70928 48276
rect 70974 48230 71000 48276
rect 70813 48172 71000 48230
rect 70813 48126 70824 48172
rect 70870 48126 70928 48172
rect 70974 48126 71000 48172
rect 70813 48068 71000 48126
rect 70813 48022 70824 48068
rect 70870 48022 70928 48068
rect 70974 48022 71000 48068
rect 70813 47964 71000 48022
rect 70813 47918 70824 47964
rect 70870 47918 70928 47964
rect 70974 47918 71000 47964
rect 70813 47860 71000 47918
rect 70813 47814 70824 47860
rect 70870 47814 70928 47860
rect 70974 47814 71000 47860
rect 70813 47756 71000 47814
rect 70813 47710 70824 47756
rect 70870 47710 70928 47756
rect 70974 47710 71000 47756
rect 70813 47652 71000 47710
rect 70813 47606 70824 47652
rect 70870 47606 70928 47652
rect 70974 47606 71000 47652
rect 70813 47548 71000 47606
rect 70813 47502 70824 47548
rect 70870 47502 70928 47548
rect 70974 47502 71000 47548
rect 70813 47444 71000 47502
rect 70813 47398 70824 47444
rect 70870 47398 70928 47444
rect 70974 47398 71000 47444
rect 70813 47340 71000 47398
rect 70813 47294 70824 47340
rect 70870 47294 70928 47340
rect 70974 47294 71000 47340
rect 70813 47236 71000 47294
rect 70813 47190 70824 47236
rect 70870 47190 70928 47236
rect 70974 47190 71000 47236
rect 70813 47132 71000 47190
rect 70813 47086 70824 47132
rect 70870 47086 70928 47132
rect 70974 47086 71000 47132
rect 70813 47028 71000 47086
rect 70813 46982 70824 47028
rect 70870 46982 70928 47028
rect 70974 46982 71000 47028
rect 70813 46924 71000 46982
rect 70813 46878 70824 46924
rect 70870 46878 70928 46924
rect 70974 46878 71000 46924
rect 70813 46820 71000 46878
rect 70813 46774 70824 46820
rect 70870 46774 70928 46820
rect 70974 46774 71000 46820
rect 70813 46716 71000 46774
rect 70813 46670 70824 46716
rect 70870 46670 70928 46716
rect 70974 46670 71000 46716
rect 70813 46612 71000 46670
rect 70813 46566 70824 46612
rect 70870 46566 70928 46612
rect 70974 46566 71000 46612
rect 70813 46508 71000 46566
rect 70813 46462 70824 46508
rect 70870 46462 70928 46508
rect 70974 46462 71000 46508
rect 70813 46404 71000 46462
rect 70813 46358 70824 46404
rect 70870 46358 70928 46404
rect 70974 46358 71000 46404
rect 70813 46300 71000 46358
rect 70813 46254 70824 46300
rect 70870 46254 70928 46300
rect 70974 46254 71000 46300
rect 70813 46196 71000 46254
rect 70813 46150 70824 46196
rect 70870 46150 70928 46196
rect 70974 46150 71000 46196
rect 70813 46092 71000 46150
rect 70813 46046 70824 46092
rect 70870 46046 70928 46092
rect 70974 46046 71000 46092
rect 70813 45988 71000 46046
rect 70813 45942 70824 45988
rect 70870 45942 70928 45988
rect 70974 45942 71000 45988
rect 70813 45884 71000 45942
rect 70813 45838 70824 45884
rect 70870 45838 70928 45884
rect 70974 45838 71000 45884
rect 70813 45780 71000 45838
rect 70813 45734 70824 45780
rect 70870 45734 70928 45780
rect 70974 45734 71000 45780
rect 70813 45676 71000 45734
rect 70813 45630 70824 45676
rect 70870 45630 70928 45676
rect 70974 45630 71000 45676
rect 70813 45572 71000 45630
rect 70813 45526 70824 45572
rect 70870 45526 70928 45572
rect 70974 45526 71000 45572
rect 70813 45468 71000 45526
rect 70813 45422 70824 45468
rect 70870 45422 70928 45468
rect 70974 45422 71000 45468
rect 70813 45364 71000 45422
rect 70813 45318 70824 45364
rect 70870 45318 70928 45364
rect 70974 45318 71000 45364
rect 70813 45260 71000 45318
rect 70813 45214 70824 45260
rect 70870 45214 70928 45260
rect 70974 45214 71000 45260
rect 70813 45156 71000 45214
rect 70813 45110 70824 45156
rect 70870 45110 70928 45156
rect 70974 45110 71000 45156
rect 70813 45052 71000 45110
rect 70813 45006 70824 45052
rect 70870 45006 70928 45052
rect 70974 45006 71000 45052
rect 70813 44948 71000 45006
tri 13108 44740 13216 44848 ne
rect 13216 44828 13280 44848
tri 13280 44828 13372 44920 sw
rect 70813 44902 70824 44948
rect 70870 44902 70928 44948
rect 70974 44902 71000 44948
rect 70813 44844 71000 44902
rect 13216 44824 13372 44828
rect 13216 44778 13254 44824
rect 13300 44778 13372 44824
rect 13216 44740 13372 44778
tri 13216 44584 13372 44740 ne
tri 13372 44692 13508 44828 sw
rect 70813 44798 70824 44844
rect 70870 44798 70928 44844
rect 70974 44798 71000 44844
rect 70813 44740 71000 44798
rect 70813 44694 70824 44740
rect 70870 44694 70928 44740
rect 70974 44694 71000 44740
rect 13372 44646 13386 44692
rect 13432 44646 13508 44692
rect 13372 44584 13508 44646
tri 13508 44584 13616 44692 sw
rect 70813 44636 71000 44694
rect 70813 44590 70824 44636
rect 70870 44590 70928 44636
rect 70974 44590 71000 44636
tri 13372 44486 13470 44584 ne
rect 13470 44560 13616 44584
rect 13470 44514 13518 44560
rect 13564 44514 13616 44560
rect 13470 44486 13616 44514
tri 13470 44340 13616 44486 ne
tri 13616 44428 13772 44584 sw
rect 70813 44532 71000 44590
rect 70813 44486 70824 44532
rect 70870 44486 70928 44532
rect 70974 44486 71000 44532
rect 70813 44428 71000 44486
rect 13616 44382 13650 44428
rect 13696 44382 13772 44428
rect 13616 44340 13772 44382
tri 13616 44220 13736 44340 ne
rect 13736 44324 13772 44340
tri 13772 44324 13876 44428 sw
rect 70813 44382 70824 44428
rect 70870 44382 70928 44428
rect 70974 44382 71000 44428
rect 70813 44324 71000 44382
rect 13736 44296 13876 44324
rect 13736 44250 13782 44296
rect 13828 44250 13876 44296
rect 13736 44220 13876 44250
tri 13736 44096 13860 44220 ne
rect 13860 44164 13876 44220
tri 13876 44164 14036 44324 sw
rect 70813 44278 70824 44324
rect 70870 44278 70928 44324
rect 70974 44278 71000 44324
rect 70813 44220 71000 44278
rect 70813 44174 70824 44220
rect 70870 44174 70928 44220
rect 70974 44174 71000 44220
rect 13860 44118 13914 44164
rect 13960 44118 14036 44164
rect 13860 44096 14036 44118
tri 13860 43966 13990 44096 ne
rect 13990 44070 14036 44096
tri 14036 44070 14130 44164 sw
rect 70813 44116 71000 44174
rect 70813 44070 70824 44116
rect 70870 44070 70928 44116
rect 70974 44070 71000 44116
rect 13990 44032 14130 44070
rect 13990 43986 14046 44032
rect 14092 43986 14130 44032
rect 13990 43966 14130 43986
tri 13990 43852 14104 43966 ne
rect 14104 43900 14130 43966
tri 14130 43900 14300 44070 sw
rect 70813 44012 71000 44070
rect 70813 43966 70824 44012
rect 70870 43966 70928 44012
rect 70974 43966 71000 44012
rect 70813 43908 71000 43966
rect 14104 43854 14178 43900
rect 14224 43854 14300 43900
rect 14104 43852 14300 43854
tri 14104 43700 14256 43852 ne
rect 14256 43768 14300 43852
tri 14300 43768 14432 43900 sw
rect 70813 43862 70824 43908
rect 70870 43862 70928 43908
rect 70974 43862 71000 43908
rect 70813 43804 71000 43862
rect 14256 43722 14310 43768
rect 14356 43722 14432 43768
rect 14256 43700 14432 43722
tri 14256 43550 14406 43700 ne
rect 14406 43636 14432 43700
tri 14432 43636 14564 43768 sw
rect 70813 43758 70824 43804
rect 70870 43758 70928 43804
rect 70974 43758 71000 43804
rect 70813 43700 71000 43758
rect 70813 43654 70824 43700
rect 70870 43654 70928 43700
rect 70974 43654 71000 43700
rect 14406 43590 14442 43636
rect 14488 43590 14564 43636
rect 14406 43550 14564 43590
tri 14406 43446 14510 43550 ne
rect 14510 43504 14564 43550
tri 14564 43504 14696 43636 sw
rect 70813 43596 71000 43654
rect 70813 43550 70824 43596
rect 70870 43550 70928 43596
rect 70974 43550 71000 43596
rect 14510 43458 14574 43504
rect 14620 43458 14696 43504
rect 14510 43446 14696 43458
tri 14510 43284 14672 43446 ne
rect 14672 43372 14696 43446
tri 14696 43372 14828 43504 sw
rect 70813 43492 71000 43550
rect 70813 43446 70824 43492
rect 70870 43446 70928 43492
rect 70974 43446 71000 43492
rect 70813 43388 71000 43446
rect 14672 43326 14706 43372
rect 14752 43326 14828 43372
rect 14672 43284 14828 43326
tri 14672 43134 14822 43284 ne
rect 14822 43240 14828 43284
tri 14828 43240 14960 43372 sw
rect 70813 43342 70824 43388
rect 70870 43342 70928 43388
rect 70974 43342 71000 43388
rect 70813 43284 71000 43342
rect 14822 43194 14838 43240
rect 14884 43194 14960 43240
rect 14822 43134 14960 43194
tri 14822 43030 14926 43134 ne
rect 14926 43120 14960 43134
tri 14960 43120 15080 43240 sw
rect 70813 43238 70824 43284
rect 70870 43238 70928 43284
rect 70974 43238 71000 43284
rect 70813 43180 71000 43238
rect 70813 43134 70824 43180
rect 70870 43134 70928 43180
rect 70974 43134 71000 43180
rect 14926 43108 15080 43120
rect 14926 43062 14970 43108
rect 15016 43062 15080 43108
rect 14926 43030 15080 43062
tri 14926 42876 15080 43030 ne
tri 15080 42976 15224 43120 sw
rect 70813 43076 71000 43134
rect 70813 43030 70824 43076
rect 70870 43030 70928 43076
rect 70974 43030 71000 43076
rect 15080 42930 15102 42976
rect 15148 42930 15224 42976
rect 15080 42876 15224 42930
tri 15080 42764 15192 42876 ne
rect 15192 42868 15224 42876
tri 15224 42868 15332 42976 sw
rect 70813 42972 71000 43030
rect 70813 42926 70824 42972
rect 70870 42926 70928 42972
rect 70974 42926 71000 42972
rect 70813 42868 71000 42926
rect 15192 42844 15332 42868
rect 15192 42798 15234 42844
rect 15280 42798 15332 42844
rect 15192 42764 15332 42798
tri 15192 42632 15324 42764 ne
rect 15324 42712 15332 42764
tri 15332 42712 15488 42868 sw
rect 70813 42822 70824 42868
rect 70870 42822 70928 42868
rect 70974 42822 71000 42868
rect 70813 42764 71000 42822
rect 70813 42718 70824 42764
rect 70870 42718 70928 42764
rect 70974 42718 71000 42764
rect 15324 42666 15366 42712
rect 15412 42666 15488 42712
rect 15324 42632 15488 42666
tri 15324 42510 15446 42632 ne
rect 15446 42614 15488 42632
tri 15488 42614 15586 42712 sw
rect 70813 42660 71000 42718
rect 70813 42614 70824 42660
rect 70870 42614 70928 42660
rect 70974 42614 71000 42660
rect 15446 42580 15586 42614
rect 15446 42534 15498 42580
rect 15544 42534 15586 42580
rect 15446 42510 15586 42534
tri 15446 42388 15568 42510 ne
rect 15568 42448 15586 42510
tri 15586 42448 15752 42614 sw
rect 70813 42556 71000 42614
rect 70813 42510 70824 42556
rect 70870 42510 70928 42556
rect 70974 42510 71000 42556
rect 70813 42452 71000 42510
rect 15568 42402 15630 42448
rect 15676 42402 15752 42448
rect 15568 42388 15752 42402
tri 15568 42244 15712 42388 ne
rect 15712 42348 15752 42388
tri 15752 42348 15852 42448 sw
rect 70813 42406 70824 42452
rect 70870 42406 70928 42452
rect 70974 42406 71000 42452
rect 70813 42348 71000 42406
rect 15712 42316 15852 42348
rect 15712 42270 15762 42316
rect 15808 42270 15852 42316
rect 15712 42244 15852 42270
tri 15712 42138 15818 42244 ne
rect 15818 42184 15852 42244
tri 15852 42184 16016 42348 sw
rect 70813 42302 70824 42348
rect 70870 42302 70928 42348
rect 70974 42302 71000 42348
rect 70813 42244 71000 42302
rect 70813 42198 70824 42244
rect 70870 42198 70928 42244
rect 70974 42198 71000 42244
rect 15818 42138 15894 42184
rect 15940 42138 16016 42184
tri 15818 41990 15966 42138 ne
rect 15966 42052 16016 42138
tri 16016 42052 16148 42184 sw
rect 70813 42140 71000 42198
rect 70813 42094 70824 42140
rect 70870 42094 70928 42140
rect 70974 42094 71000 42140
rect 15966 42006 16026 42052
rect 16072 42006 16148 42052
rect 15966 41990 16148 42006
tri 15966 41828 16128 41990 ne
rect 16128 41920 16148 41990
tri 16148 41920 16280 42052 sw
rect 70813 42036 71000 42094
rect 70813 41990 70824 42036
rect 70870 41990 70928 42036
rect 70974 41990 71000 42036
rect 70813 41932 71000 41990
rect 16128 41874 16158 41920
rect 16204 41874 16280 41920
rect 16128 41828 16280 41874
tri 16128 41678 16278 41828 ne
rect 16278 41788 16280 41828
tri 16280 41788 16412 41920 sw
rect 70813 41886 70824 41932
rect 70870 41886 70928 41932
rect 70974 41886 71000 41932
rect 70813 41828 71000 41886
rect 16278 41742 16290 41788
rect 16336 41742 16412 41788
rect 16278 41678 16412 41742
tri 16278 41574 16382 41678 ne
rect 16382 41656 16412 41678
tri 16412 41656 16544 41788 sw
rect 70813 41782 70824 41828
rect 70870 41782 70928 41828
rect 70974 41782 71000 41828
rect 70813 41724 71000 41782
rect 70813 41678 70824 41724
rect 70870 41678 70928 41724
rect 70974 41678 71000 41724
rect 16382 41610 16422 41656
rect 16468 41610 16544 41656
rect 16382 41574 16544 41610
tri 16382 41412 16544 41574 ne
tri 16544 41524 16676 41656 sw
rect 70813 41620 71000 41678
rect 70813 41574 70824 41620
rect 70870 41574 70928 41620
rect 70974 41574 71000 41620
rect 16544 41478 16554 41524
rect 16600 41478 16676 41524
rect 16544 41412 16676 41478
tri 16676 41412 16788 41524 sw
rect 70813 41516 71000 41574
rect 70813 41470 70824 41516
rect 70870 41470 70928 41516
rect 70974 41470 71000 41516
rect 70813 41412 71000 41470
tri 16544 41308 16648 41412 ne
rect 16648 41392 16788 41412
rect 16648 41346 16686 41392
rect 16732 41346 16788 41392
rect 16648 41308 16788 41346
tri 16648 41168 16788 41308 ne
tri 16788 41260 16940 41412 sw
rect 70813 41366 70824 41412
rect 70870 41366 70928 41412
rect 70974 41366 71000 41412
rect 70813 41308 71000 41366
rect 70813 41262 70824 41308
rect 70870 41262 70928 41308
rect 70974 41262 71000 41308
rect 16788 41214 16818 41260
rect 16864 41214 16940 41260
rect 16788 41168 16940 41214
tri 16788 41054 16902 41168 ne
rect 16902 41158 16940 41168
tri 16940 41158 17042 41260 sw
rect 70813 41204 71000 41262
rect 70813 41158 70824 41204
rect 70870 41158 70928 41204
rect 70974 41158 71000 41204
rect 16902 41128 17042 41158
rect 16902 41082 16950 41128
rect 16996 41082 17042 41128
rect 16902 41054 17042 41082
tri 16902 40924 17032 41054 ne
rect 17032 40996 17042 41054
tri 17042 40996 17204 41158 sw
rect 70813 41100 71000 41158
rect 70813 41054 70824 41100
rect 70870 41054 70928 41100
rect 70974 41054 71000 41100
rect 70813 40996 71000 41054
rect 17032 40950 17082 40996
rect 17128 40950 17204 40996
rect 17032 40924 17204 40950
tri 17032 40788 17168 40924 ne
rect 17168 40892 17204 40924
tri 17204 40892 17308 40996 sw
rect 70813 40950 70824 40996
rect 70870 40950 70928 40996
rect 70974 40950 71000 40996
rect 70813 40892 71000 40950
rect 17168 40864 17308 40892
rect 17168 40818 17214 40864
rect 17260 40818 17308 40864
rect 17168 40788 17308 40818
tri 17168 40680 17276 40788 ne
rect 17276 40732 17308 40788
tri 17308 40732 17468 40892 sw
rect 70813 40846 70824 40892
rect 70870 40846 70928 40892
rect 70974 40846 71000 40892
rect 70813 40788 71000 40846
rect 70813 40742 70824 40788
rect 70870 40742 70928 40788
rect 70974 40742 71000 40788
rect 17276 40686 17346 40732
rect 17392 40686 17468 40732
rect 17276 40680 17468 40686
tri 17276 40534 17422 40680 ne
rect 17422 40600 17468 40680
tri 17468 40600 17600 40732 sw
rect 70813 40684 71000 40742
rect 70813 40638 70824 40684
rect 70870 40638 70928 40684
rect 70974 40638 71000 40684
rect 17422 40554 17478 40600
rect 17524 40554 17600 40600
rect 17422 40534 17600 40554
tri 17422 40372 17584 40534 ne
rect 17584 40468 17600 40534
tri 17600 40468 17732 40600 sw
rect 70813 40580 71000 40638
rect 70813 40534 70824 40580
rect 70870 40534 70928 40580
rect 70974 40534 71000 40580
rect 70813 40476 71000 40534
rect 17584 40422 17610 40468
rect 17656 40422 17732 40468
rect 17584 40372 17732 40422
tri 17584 40268 17688 40372 ne
rect 17688 40336 17732 40372
tri 17732 40336 17864 40468 sw
rect 70813 40430 70824 40476
rect 70870 40430 70928 40476
rect 70974 40430 71000 40476
rect 70813 40372 71000 40430
rect 17688 40290 17742 40336
rect 17788 40290 17864 40336
rect 17688 40268 17864 40290
tri 17688 40118 17838 40268 ne
rect 17838 40204 17864 40268
tri 17864 40204 17996 40336 sw
rect 70813 40326 70824 40372
rect 70870 40326 70928 40372
rect 70974 40326 71000 40372
rect 70813 40268 71000 40326
rect 70813 40222 70824 40268
rect 70870 40222 70928 40268
rect 70974 40222 71000 40268
rect 17838 40158 17874 40204
rect 17920 40158 17996 40204
rect 17838 40118 17996 40158
tri 17838 40014 17942 40118 ne
rect 17942 40072 17996 40118
tri 17996 40072 18128 40204 sw
rect 70813 40164 71000 40222
rect 70813 40118 70824 40164
rect 70870 40118 70928 40164
rect 70974 40118 71000 40164
rect 17942 40026 18006 40072
rect 18052 40026 18128 40072
rect 17942 40014 18128 40026
tri 17942 39852 18104 40014 ne
rect 18104 39948 18128 40014
tri 18128 39948 18252 40072 sw
rect 70813 40060 71000 40118
rect 70813 40014 70824 40060
rect 70870 40014 70928 40060
rect 70974 40014 71000 40060
rect 70813 39956 71000 40014
rect 18104 39940 18252 39948
rect 18104 39894 18138 39940
rect 18184 39894 18252 39940
rect 18104 39852 18252 39894
tri 18104 39704 18252 39852 ne
tri 18252 39808 18392 39948 sw
rect 70813 39910 70824 39956
rect 70870 39910 70928 39956
rect 70974 39910 71000 39956
rect 70813 39852 71000 39910
rect 18252 39762 18270 39808
rect 18316 39762 18392 39808
rect 18252 39704 18392 39762
tri 18252 39598 18358 39704 ne
rect 18358 39702 18392 39704
tri 18392 39702 18498 39808 sw
rect 70813 39806 70824 39852
rect 70870 39806 70928 39852
rect 70974 39806 71000 39852
rect 70813 39748 71000 39806
rect 70813 39702 70824 39748
rect 70870 39702 70928 39748
rect 70974 39702 71000 39748
rect 18358 39676 18498 39702
rect 18358 39630 18402 39676
rect 18448 39630 18498 39676
rect 18358 39598 18498 39630
tri 18358 39460 18496 39598 ne
rect 18496 39544 18498 39598
tri 18498 39544 18656 39702 sw
rect 70813 39644 71000 39702
rect 70813 39598 70824 39644
rect 70870 39598 70928 39644
rect 70974 39598 71000 39644
rect 18496 39498 18534 39544
rect 18580 39498 18656 39544
rect 18496 39460 18656 39498
tri 18496 39332 18624 39460 ne
rect 18624 39436 18656 39460
tri 18656 39436 18764 39544 sw
rect 70813 39540 71000 39598
rect 70813 39494 70824 39540
rect 70870 39494 70928 39540
rect 70974 39494 71000 39540
rect 70813 39436 71000 39494
rect 18624 39412 18764 39436
rect 18624 39366 18666 39412
rect 18712 39366 18764 39412
rect 18624 39332 18764 39366
tri 18624 39216 18740 39332 ne
rect 18740 39280 18764 39332
tri 18764 39280 18920 39436 sw
rect 70813 39390 70824 39436
rect 70870 39390 70928 39436
rect 70974 39390 71000 39436
rect 70813 39332 71000 39390
rect 70813 39286 70824 39332
rect 70870 39286 70928 39332
rect 70974 39286 71000 39332
rect 18740 39234 18798 39280
rect 18844 39234 18920 39280
rect 18740 39216 18920 39234
tri 18740 39078 18878 39216 ne
rect 18878 39182 18920 39216
tri 18920 39182 19018 39280 sw
rect 70813 39228 71000 39286
rect 70813 39182 70824 39228
rect 70870 39182 70928 39228
rect 70974 39182 71000 39228
rect 18878 39148 19018 39182
rect 18878 39102 18930 39148
rect 18976 39102 19018 39148
rect 18878 39078 19018 39102
tri 18878 38970 18986 39078 ne
rect 18986 39016 19018 39078
tri 19018 39016 19184 39182 sw
rect 70813 39124 71000 39182
rect 70813 39078 70824 39124
rect 70870 39078 70928 39124
rect 70974 39078 71000 39124
rect 70813 39020 71000 39078
rect 18986 38970 19062 39016
rect 19108 38970 19184 39016
tri 18986 38812 19144 38970 ne
rect 19144 38884 19184 38970
tri 19184 38884 19316 39016 sw
rect 70813 38974 70824 39020
rect 70870 38974 70928 39020
rect 70974 38974 71000 39020
rect 70813 38916 71000 38974
rect 19144 38838 19194 38884
rect 19240 38838 19316 38884
rect 19144 38812 19316 38838
tri 19144 38662 19294 38812 ne
rect 19294 38752 19316 38812
tri 19316 38752 19448 38884 sw
rect 70813 38870 70824 38916
rect 70870 38870 70928 38916
rect 70974 38870 71000 38916
rect 70813 38812 71000 38870
rect 70813 38766 70824 38812
rect 70870 38766 70928 38812
rect 70974 38766 71000 38812
rect 19294 38706 19326 38752
rect 19372 38706 19448 38752
rect 19294 38662 19448 38706
tri 19294 38558 19398 38662 ne
rect 19398 38620 19448 38662
tri 19448 38620 19580 38752 sw
rect 70813 38708 71000 38766
rect 70813 38662 70824 38708
rect 70870 38662 70928 38708
rect 70974 38662 71000 38708
rect 19398 38574 19458 38620
rect 19504 38574 19580 38620
rect 19398 38558 19580 38574
tri 19398 38396 19560 38558 ne
rect 19560 38488 19580 38558
tri 19580 38488 19712 38620 sw
rect 70813 38604 71000 38662
rect 70813 38558 70824 38604
rect 70870 38558 70928 38604
rect 70974 38558 71000 38604
rect 70813 38500 71000 38558
rect 19560 38442 19590 38488
rect 19636 38442 19712 38488
rect 19560 38396 19712 38442
tri 19560 38246 19710 38396 ne
rect 19710 38356 19712 38396
tri 19712 38356 19844 38488 sw
rect 70813 38454 70824 38500
rect 70870 38454 70928 38500
rect 70974 38454 71000 38500
rect 70813 38396 71000 38454
rect 19710 38310 19722 38356
rect 19768 38310 19844 38356
rect 19710 38246 19844 38310
tri 19710 38142 19814 38246 ne
rect 19814 38240 19844 38246
tri 19844 38240 19960 38356 sw
rect 70813 38350 70824 38396
rect 70870 38350 70928 38396
rect 70974 38350 71000 38396
rect 70813 38292 71000 38350
rect 70813 38246 70824 38292
rect 70870 38246 70928 38292
rect 70974 38246 71000 38292
rect 19814 38224 19960 38240
rect 19814 38178 19854 38224
rect 19900 38178 19960 38224
rect 19814 38142 19960 38178
tri 19814 37996 19960 38142 ne
tri 19960 38092 20108 38240 sw
rect 70813 38188 71000 38246
rect 70813 38142 70824 38188
rect 70870 38142 70928 38188
rect 70974 38142 71000 38188
rect 19960 38046 19986 38092
rect 20032 38046 20108 38092
rect 19960 37996 20108 38046
tri 19960 37876 20080 37996 ne
rect 20080 37980 20108 37996
tri 20108 37980 20220 38092 sw
rect 70813 38084 71000 38142
rect 70813 38038 70824 38084
rect 70870 38038 70928 38084
rect 70974 38038 71000 38084
rect 70813 37980 71000 38038
rect 20080 37960 20220 37980
rect 20080 37914 20118 37960
rect 20164 37914 20220 37960
rect 20080 37876 20220 37914
tri 20080 37752 20204 37876 ne
rect 20204 37828 20220 37876
tri 20220 37828 20372 37980 sw
rect 70813 37934 70824 37980
rect 70870 37934 70928 37980
rect 70974 37934 71000 37980
rect 70813 37876 71000 37934
rect 70813 37830 70824 37876
rect 70870 37830 70928 37876
rect 70974 37830 71000 37876
rect 20204 37782 20250 37828
rect 20296 37782 20372 37828
rect 20204 37752 20372 37782
tri 20204 37622 20334 37752 ne
rect 20334 37726 20372 37752
tri 20372 37726 20474 37828 sw
rect 70813 37772 71000 37830
rect 70813 37726 70824 37772
rect 70870 37726 70928 37772
rect 70974 37726 71000 37772
rect 20334 37696 20474 37726
rect 20334 37650 20382 37696
rect 20428 37650 20474 37696
rect 20334 37622 20474 37650
tri 20334 37508 20448 37622 ne
rect 20448 37564 20474 37622
tri 20474 37564 20636 37726 sw
rect 70813 37668 71000 37726
rect 70813 37622 70824 37668
rect 70870 37622 70928 37668
rect 70974 37622 71000 37668
rect 70813 37564 71000 37622
rect 20448 37518 20514 37564
rect 20560 37518 20636 37564
rect 20448 37508 20636 37518
tri 20448 37356 20600 37508 ne
rect 20600 37460 20636 37508
tri 20636 37460 20740 37564 sw
rect 70813 37518 70824 37564
rect 70870 37518 70928 37564
rect 70974 37518 71000 37564
rect 70813 37460 71000 37518
rect 20600 37432 20740 37460
rect 20600 37386 20646 37432
rect 20692 37386 20740 37432
rect 20600 37356 20740 37386
tri 20600 37252 20704 37356 ne
rect 20704 37300 20740 37356
tri 20740 37300 20900 37460 sw
rect 70813 37414 70824 37460
rect 70870 37414 70928 37460
rect 70974 37414 71000 37460
rect 70813 37356 71000 37414
rect 70813 37310 70824 37356
rect 70870 37310 70928 37356
rect 70974 37310 71000 37356
rect 20704 37254 20778 37300
rect 20824 37254 20900 37300
rect 20704 37252 20900 37254
tri 20704 37102 20854 37252 ne
rect 20854 37168 20900 37252
tri 20900 37168 21032 37300 sw
rect 70813 37252 71000 37310
rect 70813 37206 70824 37252
rect 70870 37206 70928 37252
rect 70974 37206 71000 37252
rect 20854 37122 20910 37168
rect 20956 37122 21032 37168
rect 20854 37102 21032 37122
tri 20854 36940 21016 37102 ne
rect 21016 37036 21032 37102
tri 21032 37036 21164 37168 sw
rect 70813 37148 71000 37206
rect 70813 37102 70824 37148
rect 70870 37102 70928 37148
rect 70974 37102 71000 37148
rect 70813 37044 71000 37102
rect 21016 36990 21042 37036
rect 21088 36990 21164 37036
rect 21016 36940 21164 36990
tri 21016 36836 21120 36940 ne
rect 21120 36904 21164 36940
tri 21164 36904 21296 37036 sw
rect 70813 36998 70824 37044
rect 70870 36998 70928 37044
rect 70974 36998 71000 37044
rect 70813 36940 71000 36998
rect 21120 36858 21174 36904
rect 21220 36858 21296 36904
rect 21120 36836 21296 36858
tri 21120 36686 21270 36836 ne
rect 21270 36776 21296 36836
tri 21296 36776 21424 36904 sw
rect 70813 36894 70824 36940
rect 70870 36894 70928 36940
rect 70974 36894 71000 36940
rect 70813 36836 71000 36894
rect 70813 36790 70824 36836
rect 70870 36790 70928 36836
rect 70974 36790 71000 36836
rect 21270 36772 21424 36776
rect 21270 36726 21306 36772
rect 21352 36726 21424 36772
rect 21270 36686 21424 36726
tri 21270 36532 21424 36686 ne
tri 21424 36640 21560 36776 sw
rect 70813 36732 71000 36790
rect 70813 36686 70824 36732
rect 70870 36686 70928 36732
rect 70974 36686 71000 36732
rect 21424 36594 21438 36640
rect 21484 36594 21560 36640
rect 21424 36532 21560 36594
tri 21424 36420 21536 36532 ne
rect 21536 36524 21560 36532
tri 21560 36524 21676 36640 sw
rect 70813 36628 71000 36686
rect 70813 36582 70824 36628
rect 70870 36582 70928 36628
rect 70974 36582 71000 36628
rect 70813 36524 71000 36582
rect 21536 36508 21676 36524
rect 21536 36462 21570 36508
rect 21616 36462 21676 36508
rect 21536 36420 21676 36462
tri 21536 36288 21668 36420 ne
rect 21668 36376 21676 36420
tri 21676 36376 21824 36524 sw
rect 70813 36478 70824 36524
rect 70870 36478 70928 36524
rect 70974 36478 71000 36524
rect 70813 36420 71000 36478
rect 21668 36330 21702 36376
rect 21748 36330 21824 36376
rect 21668 36288 21824 36330
tri 21668 36166 21790 36288 ne
rect 21790 36270 21824 36288
tri 21824 36270 21930 36376 sw
rect 70813 36374 70824 36420
rect 70870 36374 70928 36420
rect 70974 36374 71000 36420
rect 70813 36316 71000 36374
rect 70813 36270 70824 36316
rect 70870 36270 70928 36316
rect 70974 36270 71000 36316
rect 21790 36244 21930 36270
rect 21790 36198 21834 36244
rect 21880 36198 21930 36244
rect 21790 36166 21930 36198
tri 21790 36044 21912 36166 ne
rect 21912 36112 21930 36166
tri 21930 36112 22088 36270 sw
rect 70813 36212 71000 36270
rect 70813 36166 70824 36212
rect 70870 36166 70928 36212
rect 70974 36166 71000 36212
rect 21912 36066 21966 36112
rect 22012 36066 22088 36112
rect 21912 36044 22088 36066
tri 21912 35900 22056 36044 ne
rect 22056 36004 22088 36044
tri 22088 36004 22196 36112 sw
rect 70813 36108 71000 36166
rect 70813 36062 70824 36108
rect 70870 36062 70928 36108
rect 70974 36062 71000 36108
rect 70813 36004 71000 36062
rect 22056 35980 22196 36004
rect 22056 35934 22098 35980
rect 22144 35934 22196 35980
rect 22056 35900 22196 35934
tri 22056 35796 22160 35900 ne
rect 22160 35848 22196 35900
tri 22196 35848 22352 36004 sw
rect 70813 35958 70824 36004
rect 70870 35958 70928 36004
rect 70974 35958 71000 36004
rect 70813 35900 71000 35958
rect 70813 35854 70824 35900
rect 70870 35854 70928 35900
rect 70974 35854 71000 35900
rect 22160 35802 22230 35848
rect 22276 35802 22352 35848
rect 22160 35796 22352 35802
tri 22160 35646 22310 35796 ne
rect 22310 35716 22352 35796
tri 22352 35716 22484 35848 sw
rect 70813 35796 71000 35854
rect 70813 35750 70824 35796
rect 70870 35750 70928 35796
rect 70974 35750 71000 35796
rect 22310 35670 22362 35716
rect 22408 35670 22484 35716
rect 22310 35646 22484 35670
tri 22310 35484 22472 35646 ne
rect 22472 35584 22484 35646
tri 22484 35584 22616 35716 sw
rect 70813 35692 71000 35750
rect 70813 35646 70824 35692
rect 70870 35646 70928 35692
rect 70974 35646 71000 35692
rect 70813 35588 71000 35646
rect 22472 35538 22494 35584
rect 22540 35538 22616 35584
rect 22472 35484 22616 35538
tri 22472 35380 22576 35484 ne
rect 22576 35452 22616 35484
tri 22616 35452 22748 35584 sw
rect 70813 35542 70824 35588
rect 70870 35542 70928 35588
rect 70974 35542 71000 35588
rect 70813 35484 71000 35542
rect 22576 35406 22626 35452
rect 22672 35406 22748 35452
rect 22576 35380 22748 35406
tri 22576 35230 22726 35380 ne
rect 22726 35320 22748 35380
tri 22748 35320 22880 35452 sw
rect 70813 35438 70824 35484
rect 70870 35438 70928 35484
rect 70974 35438 71000 35484
rect 70813 35380 71000 35438
rect 70813 35334 70824 35380
rect 70870 35334 70928 35380
rect 70974 35334 71000 35380
rect 22726 35274 22758 35320
rect 22804 35274 22880 35320
rect 22726 35230 22880 35274
tri 22726 35126 22830 35230 ne
rect 22830 35188 22880 35230
tri 22880 35188 23012 35320 sw
rect 70813 35276 71000 35334
rect 70813 35230 70824 35276
rect 70870 35230 70928 35276
rect 70974 35230 71000 35276
rect 22830 35142 22890 35188
rect 22936 35142 23012 35188
rect 22830 35126 23012 35142
tri 22830 34964 22992 35126 ne
rect 22992 35068 23012 35126
tri 23012 35068 23132 35188 sw
rect 70813 35172 71000 35230
rect 70813 35126 70824 35172
rect 70870 35126 70928 35172
rect 70974 35126 71000 35172
rect 70813 35068 71000 35126
rect 22992 35056 23132 35068
rect 22992 35010 23022 35056
rect 23068 35010 23132 35056
rect 22992 34964 23132 35010
tri 22992 34824 23132 34964 ne
tri 23132 34924 23276 35068 sw
rect 70813 35022 70824 35068
rect 70870 35022 70928 35068
rect 70974 35022 71000 35068
rect 70813 34964 71000 35022
rect 23132 34878 23154 34924
rect 23200 34878 23276 34924
rect 23132 34824 23276 34878
tri 23132 34710 23246 34824 ne
rect 23246 34814 23276 34824
tri 23276 34814 23386 34924 sw
rect 70813 34918 70824 34964
rect 70870 34918 70928 34964
rect 70974 34918 71000 34964
rect 70813 34860 71000 34918
rect 70813 34814 70824 34860
rect 70870 34814 70928 34860
rect 70974 34814 71000 34860
rect 23246 34792 23386 34814
rect 23246 34746 23286 34792
rect 23332 34746 23386 34792
rect 23246 34710 23386 34746
tri 23246 34580 23376 34710 ne
rect 23376 34660 23386 34710
tri 23386 34660 23540 34814 sw
rect 70813 34756 71000 34814
rect 70813 34710 70824 34756
rect 70870 34710 70928 34756
rect 70974 34710 71000 34756
rect 23376 34614 23418 34660
rect 23464 34614 23540 34660
rect 23376 34580 23540 34614
tri 23376 34444 23512 34580 ne
rect 23512 34548 23540 34580
tri 23540 34548 23652 34660 sw
rect 70813 34652 71000 34710
rect 70813 34606 70824 34652
rect 70870 34606 70928 34652
rect 70974 34606 71000 34652
rect 70813 34548 71000 34606
rect 23512 34528 23652 34548
rect 23512 34482 23550 34528
rect 23596 34482 23652 34528
rect 23512 34444 23652 34482
tri 23512 34336 23620 34444 ne
rect 23620 34396 23652 34444
tri 23652 34396 23804 34548 sw
rect 70813 34502 70824 34548
rect 70870 34502 70928 34548
rect 70974 34502 71000 34548
rect 70813 34444 71000 34502
rect 70813 34398 70824 34444
rect 70870 34398 70928 34444
rect 70974 34398 71000 34444
rect 23620 34350 23682 34396
rect 23728 34350 23804 34396
rect 23620 34336 23804 34350
tri 23620 34190 23766 34336 ne
rect 23766 34294 23804 34336
tri 23804 34294 23906 34396 sw
rect 70813 34340 71000 34398
rect 70813 34294 70824 34340
rect 70870 34294 70928 34340
rect 70974 34294 71000 34340
rect 23766 34264 23906 34294
rect 23766 34218 23814 34264
rect 23860 34218 23906 34264
rect 23766 34190 23906 34218
tri 23766 34086 23870 34190 ne
rect 23870 34132 23906 34190
tri 23906 34132 24068 34294 sw
rect 70813 34236 71000 34294
rect 70813 34190 70824 34236
rect 70870 34190 70928 34236
rect 70974 34190 71000 34236
rect 70813 34132 71000 34190
rect 23870 34086 23946 34132
rect 23992 34086 24068 34132
tri 23870 33924 24032 34086 ne
rect 24032 34000 24068 34086
tri 24068 34000 24200 34132 sw
rect 70813 34086 70824 34132
rect 70870 34086 70928 34132
rect 70974 34086 71000 34132
rect 70813 34028 71000 34086
rect 24032 33954 24078 34000
rect 24124 33954 24200 34000
rect 24032 33924 24200 33954
tri 24032 33774 24182 33924 ne
rect 24182 33868 24200 33924
tri 24200 33868 24332 34000 sw
rect 70813 33982 70824 34028
rect 70870 33982 70928 34028
rect 70974 33982 71000 34028
rect 70813 33924 71000 33982
rect 70813 33878 70824 33924
rect 70870 33878 70928 33924
rect 70974 33878 71000 33924
rect 24182 33822 24210 33868
rect 24256 33822 24332 33868
rect 24182 33774 24332 33822
tri 24182 33670 24286 33774 ne
rect 24286 33736 24332 33774
tri 24332 33736 24464 33868 sw
rect 70813 33820 71000 33878
rect 70813 33774 70824 33820
rect 70870 33774 70928 33820
rect 70974 33774 71000 33820
rect 24286 33690 24342 33736
rect 24388 33690 24464 33736
rect 24286 33670 24464 33690
tri 24286 33508 24448 33670 ne
rect 24448 33604 24464 33670
tri 24464 33604 24596 33736 sw
rect 70813 33716 71000 33774
rect 70813 33670 70824 33716
rect 70870 33670 70928 33716
rect 70974 33670 71000 33716
rect 70813 33612 71000 33670
rect 24448 33558 24474 33604
rect 24520 33558 24596 33604
rect 24448 33508 24596 33558
tri 24448 33360 24596 33508 ne
tri 24596 33472 24728 33604 sw
rect 70813 33566 70824 33612
rect 70870 33566 70928 33612
rect 70974 33566 71000 33612
rect 70813 33508 71000 33566
rect 24596 33426 24606 33472
rect 24652 33426 24728 33472
rect 24596 33360 24728 33426
tri 24596 33254 24702 33360 ne
rect 24702 33358 24728 33360
tri 24728 33358 24842 33472 sw
rect 70813 33462 70824 33508
rect 70870 33462 70928 33508
rect 70974 33462 71000 33508
rect 70813 33404 71000 33462
rect 70813 33358 70824 33404
rect 70870 33358 70928 33404
rect 70974 33358 71000 33404
rect 24702 33340 24842 33358
rect 24702 33294 24738 33340
rect 24784 33294 24842 33340
rect 24702 33254 24842 33294
tri 24702 33116 24840 33254 ne
rect 24840 33208 24842 33254
tri 24842 33208 24992 33358 sw
rect 70813 33300 71000 33358
rect 70813 33254 70824 33300
rect 70870 33254 70928 33300
rect 70974 33254 71000 33300
rect 24840 33162 24870 33208
rect 24916 33162 24992 33208
rect 24840 33116 24992 33162
tri 24840 32988 24968 33116 ne
rect 24968 33092 24992 33116
tri 24992 33092 25108 33208 sw
rect 70813 33196 71000 33254
rect 70813 33150 70824 33196
rect 70870 33150 70928 33196
rect 70974 33150 71000 33196
rect 70813 33092 71000 33150
rect 24968 33076 25108 33092
rect 24968 33030 25002 33076
rect 25048 33030 25108 33076
rect 24968 32988 25108 33030
tri 24968 32872 25084 32988 ne
rect 25084 32944 25108 32988
tri 25108 32944 25256 33092 sw
rect 70813 33046 70824 33092
rect 70870 33046 70928 33092
rect 70974 33046 71000 33092
rect 70813 32988 71000 33046
rect 25084 32898 25134 32944
rect 25180 32898 25256 32944
rect 25084 32872 25256 32898
tri 25084 32734 25222 32872 ne
rect 25222 32838 25256 32872
tri 25256 32838 25362 32944 sw
rect 70813 32942 70824 32988
rect 70870 32942 70928 32988
rect 70974 32942 71000 32988
rect 70813 32884 71000 32942
rect 70813 32838 70824 32884
rect 70870 32838 70928 32884
rect 70974 32838 71000 32884
rect 25222 32812 25362 32838
rect 25222 32766 25266 32812
rect 25312 32766 25362 32812
rect 25222 32734 25362 32766
tri 25222 32628 25328 32734 ne
rect 25328 32680 25362 32734
tri 25362 32680 25520 32838 sw
rect 70813 32780 71000 32838
rect 70813 32734 70824 32780
rect 70870 32734 70928 32780
rect 70974 32734 71000 32780
rect 25328 32634 25398 32680
rect 25444 32634 25520 32680
rect 25328 32628 25520 32634
tri 25328 32468 25488 32628 ne
rect 25488 32548 25520 32628
tri 25520 32548 25652 32680 sw
rect 70813 32676 71000 32734
rect 70813 32630 70824 32676
rect 70870 32630 70928 32676
rect 70974 32630 71000 32676
rect 70813 32572 71000 32630
rect 25488 32502 25530 32548
rect 25576 32502 25652 32548
rect 25488 32468 25652 32502
tri 25488 32318 25638 32468 ne
rect 25638 32416 25652 32468
tri 25652 32416 25784 32548 sw
rect 70813 32526 70824 32572
rect 70870 32526 70928 32572
rect 70974 32526 71000 32572
rect 70813 32468 71000 32526
rect 70813 32422 70824 32468
rect 70870 32422 70928 32468
rect 70974 32422 71000 32468
rect 25638 32370 25662 32416
rect 25708 32370 25784 32416
rect 25638 32318 25784 32370
tri 25638 32214 25742 32318 ne
rect 25742 32284 25784 32318
tri 25784 32284 25916 32416 sw
rect 70813 32364 71000 32422
rect 70813 32318 70824 32364
rect 70870 32318 70928 32364
rect 70974 32318 71000 32364
rect 25742 32238 25794 32284
rect 25840 32238 25916 32284
rect 25742 32214 25916 32238
tri 25742 32052 25904 32214 ne
rect 25904 32152 25916 32214
tri 25916 32152 26048 32284 sw
rect 70813 32260 71000 32318
rect 70813 32214 70824 32260
rect 70870 32214 70928 32260
rect 70974 32214 71000 32260
rect 70813 32156 71000 32214
rect 25904 32106 25926 32152
rect 25972 32106 26048 32152
rect 25904 32052 26048 32106
tri 25904 31948 26008 32052 ne
rect 26008 32020 26048 32052
tri 26048 32020 26180 32152 sw
rect 70813 32110 70824 32156
rect 70870 32110 70928 32156
rect 70974 32110 71000 32156
rect 70813 32052 71000 32110
rect 26008 31974 26058 32020
rect 26104 31974 26180 32020
rect 26008 31948 26180 31974
tri 26008 31798 26158 31948 ne
rect 26158 31896 26180 31948
tri 26180 31896 26304 32020 sw
rect 70813 32006 70824 32052
rect 70870 32006 70928 32052
rect 70974 32006 71000 32052
rect 70813 31948 71000 32006
rect 70813 31902 70824 31948
rect 70870 31902 70928 31948
rect 70974 31902 71000 31948
rect 26158 31888 26304 31896
rect 26158 31842 26190 31888
rect 26236 31842 26304 31888
rect 26158 31798 26304 31842
tri 26158 31652 26304 31798 ne
tri 26304 31756 26444 31896 sw
rect 70813 31844 71000 31902
rect 70813 31798 70824 31844
rect 70870 31798 70928 31844
rect 70974 31798 71000 31844
rect 26304 31710 26322 31756
rect 26368 31710 26444 31756
rect 26304 31652 26444 31710
tri 26304 31532 26424 31652 ne
rect 26424 31636 26444 31652
tri 26444 31636 26564 31756 sw
rect 70813 31740 71000 31798
rect 70813 31694 70824 31740
rect 70870 31694 70928 31740
rect 70974 31694 71000 31740
rect 70813 31636 71000 31694
rect 26424 31624 26564 31636
rect 26424 31578 26454 31624
rect 26500 31578 26564 31624
rect 26424 31532 26564 31578
tri 26424 31408 26548 31532 ne
rect 26548 31492 26564 31532
tri 26564 31492 26708 31636 sw
rect 70813 31590 70824 31636
rect 70870 31590 70928 31636
rect 70974 31590 71000 31636
rect 70813 31532 71000 31590
rect 26548 31446 26586 31492
rect 26632 31446 26708 31492
rect 26548 31408 26708 31446
tri 26548 31278 26678 31408 ne
rect 26678 31382 26708 31408
tri 26708 31382 26818 31492 sw
rect 70813 31486 70824 31532
rect 70870 31486 70928 31532
rect 70974 31486 71000 31532
rect 70813 31428 71000 31486
rect 70813 31382 70824 31428
rect 70870 31382 70928 31428
rect 70974 31382 71000 31428
rect 26678 31360 26818 31382
rect 26678 31314 26718 31360
rect 26764 31314 26818 31360
rect 26678 31278 26818 31314
tri 26678 31164 26792 31278 ne
rect 26792 31228 26818 31278
tri 26818 31228 26972 31382 sw
rect 70813 31324 71000 31382
rect 70813 31278 70824 31324
rect 70870 31278 70928 31324
rect 70974 31278 71000 31324
rect 26792 31182 26850 31228
rect 26896 31182 26972 31228
rect 26792 31164 26972 31182
tri 26792 31012 26944 31164 ne
rect 26944 31116 26972 31164
tri 26972 31116 27084 31228 sw
rect 70813 31220 71000 31278
rect 70813 31174 70824 31220
rect 70870 31174 70928 31220
rect 70974 31174 71000 31220
rect 70813 31116 71000 31174
rect 26944 31096 27084 31116
rect 26944 31050 26982 31096
rect 27028 31050 27084 31096
rect 26944 31012 27084 31050
tri 26944 30908 27048 31012 ne
rect 27048 30964 27084 31012
tri 27084 30964 27236 31116 sw
rect 70813 31070 70824 31116
rect 70870 31070 70928 31116
rect 70974 31070 71000 31116
rect 70813 31012 71000 31070
rect 70813 30966 70824 31012
rect 70870 30966 70928 31012
rect 70974 30966 71000 31012
rect 27048 30918 27114 30964
rect 27160 30918 27236 30964
rect 27048 30908 27236 30918
tri 27048 30758 27198 30908 ne
rect 27198 30832 27236 30908
tri 27236 30832 27368 30964 sw
rect 70813 30908 71000 30966
rect 70813 30862 70824 30908
rect 70870 30862 70928 30908
rect 70974 30862 71000 30908
rect 27198 30786 27246 30832
rect 27292 30786 27368 30832
rect 27198 30758 27368 30786
tri 27198 30596 27360 30758 ne
rect 27360 30700 27368 30758
tri 27368 30700 27500 30832 sw
rect 70813 30804 71000 30862
rect 70813 30758 70824 30804
rect 70870 30758 70928 30804
rect 70974 30758 71000 30804
rect 70813 30700 71000 30758
rect 27360 30654 27378 30700
rect 27424 30654 27500 30700
rect 27360 30596 27500 30654
tri 27360 30492 27464 30596 ne
rect 27464 30568 27500 30596
tri 27500 30568 27632 30700 sw
rect 70813 30654 70824 30700
rect 70870 30654 70928 30700
rect 70974 30654 71000 30700
rect 70813 30596 71000 30654
rect 27464 30522 27510 30568
rect 27556 30522 27632 30568
rect 27464 30492 27632 30522
tri 27464 30342 27614 30492 ne
rect 27614 30436 27632 30492
tri 27632 30436 27764 30568 sw
rect 70813 30550 70824 30596
rect 70870 30550 70928 30596
rect 70974 30550 71000 30596
rect 70813 30492 71000 30550
rect 70813 30446 70824 30492
rect 70870 30446 70928 30492
rect 70974 30446 71000 30492
rect 27614 30390 27642 30436
rect 27688 30390 27764 30436
rect 27614 30342 27764 30390
tri 27614 30238 27718 30342 ne
rect 27718 30304 27764 30342
tri 27764 30304 27896 30436 sw
rect 70813 30388 71000 30446
rect 70813 30342 70824 30388
rect 70870 30342 70928 30388
rect 70974 30342 71000 30388
rect 27718 30258 27774 30304
rect 27820 30258 27896 30304
rect 27718 30238 27896 30258
tri 27718 30076 27880 30238 ne
rect 27880 30180 27896 30238
tri 27896 30180 28020 30304 sw
rect 70813 30284 71000 30342
rect 70813 30238 70824 30284
rect 70870 30238 70928 30284
rect 70974 30238 71000 30284
rect 70813 30180 71000 30238
rect 27880 30172 28020 30180
rect 27880 30126 27906 30172
rect 27952 30126 28020 30172
rect 27880 30076 28020 30126
tri 27880 29944 28012 30076 ne
rect 28012 30040 28020 30076
tri 28020 30040 28160 30180 sw
rect 70813 30134 70824 30180
rect 70870 30134 70928 30180
rect 70974 30134 71000 30180
rect 70813 30076 71000 30134
rect 28012 29994 28038 30040
rect 28084 29994 28160 30040
rect 28012 29944 28160 29994
tri 28012 29822 28134 29944 ne
rect 28134 29926 28160 29944
tri 28160 29926 28274 30040 sw
rect 70813 30030 70824 30076
rect 70870 30030 70928 30076
rect 70974 30030 71000 30076
rect 70813 29972 71000 30030
rect 70813 29926 70824 29972
rect 70870 29926 70928 29972
rect 70974 29926 71000 29972
rect 28134 29908 28274 29926
rect 28134 29862 28170 29908
rect 28216 29862 28274 29908
rect 28134 29822 28274 29862
tri 28134 29700 28256 29822 ne
rect 28256 29776 28274 29822
tri 28274 29776 28424 29926 sw
rect 70813 29868 71000 29926
rect 70813 29822 70824 29868
rect 70870 29822 70928 29868
rect 70974 29822 71000 29868
rect 28256 29730 28302 29776
rect 28348 29730 28424 29776
rect 28256 29700 28424 29730
tri 28256 29556 28400 29700 ne
rect 28400 29660 28424 29700
tri 28424 29660 28540 29776 sw
rect 70813 29764 71000 29822
rect 70813 29718 70824 29764
rect 70870 29718 70928 29764
rect 70974 29718 71000 29764
rect 70813 29660 71000 29718
rect 28400 29644 28540 29660
rect 28400 29598 28434 29644
rect 28480 29598 28540 29644
rect 28400 29556 28540 29598
tri 28400 29452 28504 29556 ne
rect 28504 29512 28540 29556
tri 28540 29512 28688 29660 sw
rect 70813 29614 70824 29660
rect 70870 29614 70928 29660
rect 70974 29614 71000 29660
rect 70813 29556 71000 29614
rect 28504 29466 28566 29512
rect 28612 29466 28688 29512
rect 28504 29452 28688 29466
tri 28504 29302 28654 29452 ne
rect 28654 29406 28688 29452
tri 28688 29406 28794 29512 sw
rect 70813 29510 70824 29556
rect 70870 29510 70928 29556
rect 70974 29510 71000 29556
rect 70813 29452 71000 29510
rect 70813 29406 70824 29452
rect 70870 29406 70928 29452
rect 70974 29406 71000 29452
rect 28654 29380 28794 29406
rect 28654 29334 28698 29380
rect 28744 29334 28794 29380
rect 28654 29302 28794 29334
tri 28654 29198 28758 29302 ne
rect 28758 29248 28794 29302
tri 28794 29248 28952 29406 sw
rect 70813 29348 71000 29406
rect 70813 29302 70824 29348
rect 70870 29302 70928 29348
rect 70974 29302 71000 29348
rect 28758 29202 28830 29248
rect 28876 29202 28952 29248
rect 28758 29198 28952 29202
tri 28758 29036 28920 29198 ne
rect 28920 29116 28952 29198
tri 28952 29116 29084 29248 sw
rect 70813 29244 71000 29302
rect 70813 29198 70824 29244
rect 70870 29198 70928 29244
rect 70974 29198 71000 29244
rect 70813 29140 71000 29198
rect 28920 29070 28962 29116
rect 29008 29070 29084 29116
rect 28920 29036 29084 29070
tri 28920 28886 29070 29036 ne
rect 29070 28984 29084 29036
tri 29084 28984 29216 29116 sw
rect 70813 29094 70824 29140
rect 70870 29094 70928 29140
rect 70974 29094 71000 29140
rect 70813 29036 71000 29094
rect 70813 28990 70824 29036
rect 70870 28990 70928 29036
rect 70974 28990 71000 29036
rect 29070 28938 29094 28984
rect 29140 28938 29216 28984
rect 29070 28886 29216 28938
tri 29070 28782 29174 28886 ne
rect 29174 28852 29216 28886
tri 29216 28852 29348 28984 sw
rect 70813 28932 71000 28990
rect 70813 28886 70824 28932
rect 70870 28886 70928 28932
rect 70974 28886 71000 28932
rect 29174 28806 29226 28852
rect 29272 28806 29348 28852
rect 29174 28782 29348 28806
tri 29174 28620 29336 28782 ne
rect 29336 28724 29348 28782
tri 29348 28724 29476 28852 sw
rect 70813 28828 71000 28886
rect 70813 28782 70824 28828
rect 70870 28782 70928 28828
rect 70974 28782 71000 28828
rect 70813 28724 71000 28782
rect 29336 28720 29476 28724
rect 29336 28674 29358 28720
rect 29404 28674 29476 28720
rect 29336 28620 29476 28674
tri 29336 28480 29476 28620 ne
tri 29476 28588 29612 28724 sw
rect 70813 28678 70824 28724
rect 70870 28678 70928 28724
rect 70974 28678 71000 28724
rect 70813 28620 71000 28678
rect 29476 28542 29490 28588
rect 29536 28542 29612 28588
rect 29476 28480 29612 28542
tri 29476 28366 29590 28480 ne
rect 29590 28470 29612 28480
tri 29612 28470 29730 28588 sw
rect 70813 28574 70824 28620
rect 70870 28574 70928 28620
rect 70974 28574 71000 28620
rect 70813 28516 71000 28574
rect 70813 28470 70824 28516
rect 70870 28470 70928 28516
rect 70974 28470 71000 28516
rect 29590 28456 29730 28470
rect 29590 28410 29622 28456
rect 29668 28410 29730 28456
rect 29590 28366 29730 28410
tri 29590 28236 29720 28366 ne
rect 29720 28324 29730 28366
tri 29730 28324 29876 28470 sw
rect 70813 28412 71000 28470
rect 70813 28366 70824 28412
rect 70870 28366 70928 28412
rect 70974 28366 71000 28412
rect 29720 28278 29754 28324
rect 29800 28278 29876 28324
rect 29720 28236 29876 28278
tri 29720 28100 29856 28236 ne
rect 29856 28204 29876 28236
tri 29876 28204 29996 28324 sw
rect 70813 28308 71000 28366
rect 70813 28262 70824 28308
rect 70870 28262 70928 28308
rect 70974 28262 71000 28308
rect 70813 28204 71000 28262
rect 29856 28192 29996 28204
rect 29856 28146 29886 28192
rect 29932 28146 29996 28192
rect 29856 28100 29996 28146
tri 29856 27992 29964 28100 ne
rect 29964 28060 29996 28100
tri 29996 28060 30140 28204 sw
rect 70813 28158 70824 28204
rect 70870 28158 70928 28204
rect 70974 28158 71000 28204
rect 70813 28100 71000 28158
rect 29964 28014 30018 28060
rect 30064 28014 30140 28060
rect 29964 27992 30140 28014
tri 29964 27846 30110 27992 ne
rect 30110 27950 30140 27992
tri 30140 27950 30250 28060 sw
rect 70813 28054 70824 28100
rect 70870 28054 70928 28100
rect 70974 28054 71000 28100
rect 70813 27996 71000 28054
rect 70813 27950 70824 27996
rect 70870 27950 70928 27996
rect 70974 27950 71000 27996
rect 30110 27928 30250 27950
rect 30110 27882 30150 27928
rect 30196 27882 30250 27928
rect 30110 27846 30250 27882
tri 30110 27742 30214 27846 ne
rect 30214 27796 30250 27846
tri 30250 27796 30404 27950 sw
rect 70813 27892 71000 27950
rect 70813 27846 70824 27892
rect 70870 27846 70928 27892
rect 70974 27846 71000 27892
rect 30214 27750 30282 27796
rect 30328 27750 30404 27796
rect 30214 27742 30404 27750
tri 30214 27580 30376 27742 ne
rect 30376 27664 30404 27742
tri 30404 27664 30536 27796 sw
rect 70813 27788 71000 27846
rect 70813 27742 70824 27788
rect 70870 27742 70928 27788
rect 70974 27742 71000 27788
rect 70813 27684 71000 27742
rect 30376 27618 30414 27664
rect 30460 27618 30536 27664
rect 30376 27580 30536 27618
tri 30376 27430 30526 27580 ne
rect 30526 27532 30536 27580
tri 30536 27532 30668 27664 sw
rect 70813 27638 70824 27684
rect 70870 27638 70928 27684
rect 70974 27638 71000 27684
rect 70813 27580 71000 27638
rect 70813 27534 70824 27580
rect 70870 27534 70928 27580
rect 70974 27534 71000 27580
rect 30526 27486 30546 27532
rect 30592 27486 30668 27532
rect 30526 27430 30668 27486
tri 30526 27326 30630 27430 ne
rect 30630 27400 30668 27430
tri 30668 27400 30800 27532 sw
rect 70813 27476 71000 27534
rect 70813 27430 70824 27476
rect 70870 27430 70928 27476
rect 70974 27430 71000 27476
rect 30630 27354 30678 27400
rect 30724 27354 30800 27400
rect 30630 27326 30800 27354
tri 30630 27164 30792 27326 ne
rect 30792 27268 30800 27326
tri 30800 27268 30932 27400 sw
rect 70813 27372 71000 27430
rect 70813 27326 70824 27372
rect 70870 27326 70928 27372
rect 70974 27326 71000 27372
rect 70813 27268 71000 27326
rect 30792 27222 30810 27268
rect 30856 27222 30932 27268
rect 30792 27164 30932 27222
tri 30792 27060 30896 27164 ne
rect 30896 27136 30932 27164
tri 30932 27136 31064 27268 sw
rect 70813 27222 70824 27268
rect 70870 27222 70928 27268
rect 70974 27222 71000 27268
rect 70813 27164 71000 27222
rect 30896 27090 30942 27136
rect 30988 27090 31064 27136
rect 30896 27060 31064 27090
tri 30896 26910 31046 27060 ne
rect 31046 27014 31064 27060
tri 31064 27014 31186 27136 sw
rect 70813 27118 70824 27164
rect 70870 27118 70928 27164
rect 70974 27118 71000 27164
rect 70813 27060 71000 27118
rect 70813 27014 70824 27060
rect 70870 27014 70928 27060
rect 70974 27014 71000 27060
rect 31046 27004 31186 27014
rect 31046 26958 31074 27004
rect 31120 26958 31186 27004
rect 31046 26910 31186 26958
tri 31046 26772 31184 26910 ne
rect 31184 26872 31186 26910
tri 31186 26872 31328 27014 sw
rect 70813 26956 71000 27014
rect 70813 26910 70824 26956
rect 70870 26910 70928 26956
rect 70974 26910 71000 26956
rect 31184 26826 31206 26872
rect 31252 26826 31328 26872
rect 31184 26772 31328 26826
tri 31184 26644 31312 26772 ne
rect 31312 26748 31328 26772
tri 31328 26748 31452 26872 sw
rect 70813 26852 71000 26910
rect 70813 26806 70824 26852
rect 70870 26806 70928 26852
rect 70974 26806 71000 26852
rect 70813 26748 71000 26806
rect 31312 26740 31452 26748
rect 31312 26694 31338 26740
rect 31384 26694 31452 26740
rect 31312 26644 31452 26694
tri 31312 26528 31428 26644 ne
rect 31428 26608 31452 26644
tri 31452 26608 31592 26748 sw
rect 70813 26702 70824 26748
rect 70870 26702 70928 26748
rect 70974 26702 71000 26748
rect 70813 26644 71000 26702
rect 31428 26562 31470 26608
rect 31516 26562 31592 26608
rect 31428 26528 31592 26562
tri 31428 26390 31566 26528 ne
rect 31566 26494 31592 26528
tri 31592 26494 31706 26608 sw
rect 70813 26598 70824 26644
rect 70870 26598 70928 26644
rect 70974 26598 71000 26644
rect 70813 26540 71000 26598
rect 70813 26494 70824 26540
rect 70870 26494 70928 26540
rect 70974 26494 71000 26540
rect 31566 26476 31706 26494
rect 31566 26430 31602 26476
rect 31648 26430 31706 26476
rect 31566 26390 31706 26430
tri 31566 26284 31672 26390 ne
rect 31672 26344 31706 26390
tri 31706 26344 31856 26494 sw
rect 70813 26436 71000 26494
rect 70813 26390 70824 26436
rect 70870 26390 70928 26436
rect 70974 26390 71000 26436
rect 31672 26298 31734 26344
rect 31780 26298 31856 26344
rect 31672 26284 31856 26298
tri 31672 26124 31832 26284 ne
rect 31832 26228 31856 26284
tri 31856 26228 31972 26344 sw
rect 70813 26332 71000 26390
rect 70813 26286 70824 26332
rect 70870 26286 70928 26332
rect 70974 26286 71000 26332
rect 70813 26228 71000 26286
rect 31832 26212 31972 26228
rect 31832 26166 31866 26212
rect 31912 26166 31972 26212
rect 31832 26124 31972 26166
tri 31832 26020 31936 26124 ne
rect 31936 26080 31972 26124
tri 31972 26080 32120 26228 sw
rect 70813 26182 70824 26228
rect 70870 26182 70928 26228
rect 70974 26182 71000 26228
rect 70813 26124 71000 26182
rect 31936 26034 31998 26080
rect 32044 26034 32120 26080
rect 31936 26020 32120 26034
tri 31936 25870 32086 26020 ne
rect 32086 25948 32120 26020
tri 32120 25948 32252 26080 sw
rect 70813 26078 70824 26124
rect 70870 26078 70928 26124
rect 70974 26078 71000 26124
rect 70813 26020 71000 26078
rect 70813 25974 70824 26020
rect 70870 25974 70928 26020
rect 70974 25974 71000 26020
rect 32086 25902 32130 25948
rect 32176 25902 32252 25948
rect 32086 25870 32252 25902
tri 32086 25708 32248 25870 ne
rect 32248 25816 32252 25870
tri 32252 25816 32384 25948 sw
rect 70813 25916 71000 25974
rect 70813 25870 70824 25916
rect 70870 25870 70928 25916
rect 70974 25870 71000 25916
rect 32248 25770 32262 25816
rect 32308 25770 32384 25816
rect 32248 25708 32384 25770
tri 32248 25604 32352 25708 ne
rect 32352 25684 32384 25708
tri 32384 25684 32516 25816 sw
rect 70813 25812 71000 25870
rect 70813 25766 70824 25812
rect 70870 25766 70928 25812
rect 70974 25766 71000 25812
rect 70813 25708 71000 25766
rect 32352 25638 32394 25684
rect 32440 25638 32516 25684
rect 32352 25604 32516 25638
tri 32352 25454 32502 25604 ne
rect 32502 25552 32516 25604
tri 32516 25552 32648 25684 sw
rect 70813 25662 70824 25708
rect 70870 25662 70928 25708
rect 70974 25662 71000 25708
rect 70813 25604 71000 25662
rect 70813 25558 70824 25604
rect 70870 25558 70928 25604
rect 70974 25558 71000 25604
rect 32502 25506 32526 25552
rect 32572 25506 32648 25552
rect 32502 25454 32648 25506
tri 32502 25308 32648 25454 ne
tri 32648 25420 32780 25552 sw
rect 70813 25500 71000 25558
rect 70813 25454 70824 25500
rect 70870 25454 70928 25500
rect 70974 25454 71000 25500
rect 32648 25374 32658 25420
rect 32704 25374 32780 25420
rect 32648 25308 32780 25374
tri 32648 25188 32768 25308 ne
rect 32768 25292 32780 25308
tri 32780 25292 32908 25420 sw
rect 70813 25396 71000 25454
rect 70813 25350 70824 25396
rect 70870 25350 70928 25396
rect 70974 25350 71000 25396
rect 70813 25292 71000 25350
rect 32768 25288 32908 25292
rect 32768 25242 32790 25288
rect 32836 25242 32908 25288
rect 32768 25188 32908 25242
tri 32768 25064 32892 25188 ne
rect 32892 25156 32908 25188
tri 32908 25156 33044 25292 sw
rect 70813 25246 70824 25292
rect 70870 25246 70928 25292
rect 70974 25246 71000 25292
rect 70813 25188 71000 25246
rect 32892 25110 32922 25156
rect 32968 25110 33044 25156
rect 32892 25064 33044 25110
tri 32892 24934 33022 25064 ne
rect 33022 25038 33044 25064
tri 33044 25038 33162 25156 sw
rect 70813 25142 70824 25188
rect 70870 25142 70928 25188
rect 70974 25142 71000 25188
rect 70813 25084 71000 25142
rect 70813 25038 70824 25084
rect 70870 25038 70928 25084
rect 70974 25038 71000 25084
rect 33022 25024 33162 25038
rect 33022 24978 33054 25024
rect 33100 24978 33162 25024
rect 33022 24934 33162 24978
tri 33022 24820 33136 24934 ne
rect 33136 24892 33162 24934
tri 33162 24892 33308 25038 sw
rect 70813 24980 71000 25038
rect 70813 24934 70824 24980
rect 70870 24934 70928 24980
rect 70974 24934 71000 24980
rect 33136 24846 33186 24892
rect 33232 24846 33308 24892
rect 33136 24820 33308 24846
tri 33136 24668 33288 24820 ne
rect 33288 24772 33308 24820
tri 33308 24772 33428 24892 sw
rect 70813 24876 71000 24934
rect 70813 24830 70824 24876
rect 70870 24830 70928 24876
rect 70974 24830 71000 24876
rect 70813 24772 71000 24830
rect 33288 24760 33428 24772
rect 33288 24714 33318 24760
rect 33364 24714 33428 24760
rect 33288 24668 33428 24714
tri 33288 24564 33392 24668 ne
rect 33392 24628 33428 24668
tri 33428 24628 33572 24772 sw
rect 70813 24726 70824 24772
rect 70870 24726 70928 24772
rect 70974 24726 71000 24772
rect 70813 24668 71000 24726
rect 33392 24582 33450 24628
rect 33496 24582 33572 24628
rect 33392 24564 33572 24582
tri 33392 24414 33542 24564 ne
rect 33542 24496 33572 24564
tri 33572 24496 33704 24628 sw
rect 70813 24622 70824 24668
rect 70870 24622 70928 24668
rect 70974 24622 71000 24668
rect 70813 24564 71000 24622
rect 70813 24518 70824 24564
rect 70870 24518 70928 24564
rect 70974 24518 71000 24564
rect 33542 24450 33582 24496
rect 33628 24450 33704 24496
rect 33542 24414 33704 24450
tri 33542 24252 33704 24414 ne
tri 33704 24364 33836 24496 sw
rect 70813 24460 71000 24518
rect 70813 24414 70824 24460
rect 70870 24414 70928 24460
rect 70974 24414 71000 24460
rect 33704 24318 33714 24364
rect 33760 24318 33836 24364
rect 33704 24252 33836 24318
tri 33704 24148 33808 24252 ne
rect 33808 24232 33836 24252
tri 33836 24232 33968 24364 sw
rect 70813 24356 71000 24414
rect 70813 24310 70824 24356
rect 70870 24310 70928 24356
rect 70974 24310 71000 24356
rect 70813 24252 71000 24310
rect 33808 24186 33846 24232
rect 33892 24186 33968 24232
rect 33808 24148 33968 24186
tri 33808 23998 33958 24148 ne
rect 33958 24100 33968 24148
tri 33968 24100 34100 24232 sw
rect 70813 24206 70824 24252
rect 70870 24206 70928 24252
rect 70974 24206 71000 24252
rect 70813 24148 71000 24206
rect 70813 24102 70824 24148
rect 70870 24102 70928 24148
rect 70974 24102 71000 24148
rect 33958 24054 33978 24100
rect 34024 24054 34100 24100
rect 33958 23998 34100 24054
tri 33958 23894 34062 23998 ne
rect 34062 23968 34100 23998
tri 34100 23968 34232 24100 sw
rect 70813 24044 71000 24102
rect 70813 23998 70824 24044
rect 70870 23998 70928 24044
rect 70974 23998 71000 24044
rect 34062 23922 34110 23968
rect 34156 23922 34232 23968
rect 34062 23894 34232 23922
tri 34062 23732 34224 23894 ne
rect 34224 23836 34232 23894
tri 34232 23836 34364 23968 sw
rect 70813 23940 71000 23998
rect 70813 23894 70824 23940
rect 70870 23894 70928 23940
rect 70974 23894 71000 23940
rect 70813 23836 71000 23894
rect 34224 23790 34242 23836
rect 34288 23790 34364 23836
rect 34224 23732 34364 23790
tri 34224 23600 34356 23732 ne
rect 34356 23704 34364 23732
tri 34364 23704 34496 23836 sw
rect 70813 23790 70824 23836
rect 70870 23790 70928 23836
rect 70974 23790 71000 23836
rect 70813 23732 71000 23790
rect 34356 23658 34374 23704
rect 34420 23658 34496 23704
rect 34356 23600 34496 23658
tri 34356 23478 34478 23600 ne
rect 34478 23582 34496 23600
tri 34496 23582 34618 23704 sw
rect 70813 23686 70824 23732
rect 70870 23686 70928 23732
rect 70974 23686 71000 23732
rect 70813 23628 71000 23686
rect 70813 23582 70824 23628
rect 70870 23582 70928 23628
rect 70974 23582 71000 23628
rect 34478 23572 34618 23582
rect 34478 23526 34506 23572
rect 34552 23526 34618 23572
rect 34478 23478 34618 23526
tri 34478 23356 34600 23478 ne
rect 34600 23440 34618 23478
tri 34618 23440 34760 23582 sw
rect 70813 23524 71000 23582
rect 70813 23478 70824 23524
rect 70870 23478 70928 23524
rect 70974 23478 71000 23524
rect 34600 23394 34638 23440
rect 34684 23394 34760 23440
rect 34600 23356 34760 23394
tri 34600 23212 34744 23356 ne
rect 34744 23316 34760 23356
tri 34760 23316 34884 23440 sw
rect 70813 23420 71000 23478
rect 70813 23374 70824 23420
rect 70870 23374 70928 23420
rect 70974 23374 71000 23420
rect 70813 23316 71000 23374
rect 34744 23308 34884 23316
rect 34744 23262 34770 23308
rect 34816 23262 34884 23308
rect 34744 23212 34884 23262
tri 34744 23108 34848 23212 ne
rect 34848 23176 34884 23212
tri 34884 23176 35024 23316 sw
rect 70813 23270 70824 23316
rect 70870 23270 70928 23316
rect 70974 23270 71000 23316
rect 70813 23212 71000 23270
rect 34848 23130 34902 23176
rect 34948 23130 35024 23176
rect 34848 23108 35024 23130
tri 34848 22958 34998 23108 ne
rect 34998 23062 35024 23108
tri 35024 23062 35138 23176 sw
rect 70813 23166 70824 23212
rect 70870 23166 70928 23212
rect 70974 23166 71000 23212
rect 70813 23108 71000 23166
rect 70813 23062 70824 23108
rect 70870 23062 70928 23108
rect 70974 23062 71000 23108
rect 34998 23044 35138 23062
rect 34998 22998 35034 23044
rect 35080 22998 35138 23044
rect 34998 22958 35138 22998
tri 34998 22854 35102 22958 ne
rect 35102 22912 35138 22958
tri 35138 22912 35288 23062 sw
rect 70813 23004 71000 23062
rect 70813 22958 70824 23004
rect 70870 22958 70928 23004
rect 70974 22958 71000 23004
rect 35102 22866 35166 22912
rect 35212 22866 35288 22912
rect 35102 22854 35288 22866
tri 35102 22692 35264 22854 ne
rect 35264 22780 35288 22854
tri 35288 22780 35420 22912 sw
rect 70813 22900 71000 22958
rect 70813 22854 70824 22900
rect 70870 22854 70928 22900
rect 70974 22854 71000 22900
rect 70813 22796 71000 22854
rect 35264 22734 35298 22780
rect 35344 22734 35420 22780
rect 35264 22692 35420 22734
tri 35264 22542 35414 22692 ne
rect 35414 22648 35420 22692
tri 35420 22648 35552 22780 sw
rect 70813 22750 70824 22796
rect 70870 22750 70928 22796
rect 70974 22750 71000 22796
rect 70813 22692 71000 22750
rect 35414 22602 35430 22648
rect 35476 22602 35552 22648
rect 35414 22542 35552 22602
tri 35414 22438 35518 22542 ne
rect 35518 22516 35552 22542
tri 35552 22516 35684 22648 sw
rect 70813 22646 70824 22692
rect 70870 22646 70928 22692
rect 70974 22646 71000 22692
rect 70813 22588 71000 22646
rect 70813 22542 70824 22588
rect 70870 22542 70928 22588
rect 70974 22542 71000 22588
rect 35518 22470 35562 22516
rect 35608 22470 35684 22516
rect 35518 22438 35684 22470
tri 35518 22276 35680 22438 ne
rect 35680 22384 35684 22438
tri 35684 22384 35816 22516 sw
rect 70813 22484 71000 22542
rect 70813 22438 70824 22484
rect 70870 22438 70928 22484
rect 70974 22438 71000 22484
rect 35680 22338 35694 22384
rect 35740 22338 35816 22384
rect 35680 22276 35816 22338
tri 35680 22172 35784 22276 ne
rect 35784 22252 35816 22276
tri 35816 22252 35948 22384 sw
rect 70813 22380 71000 22438
rect 70813 22334 70824 22380
rect 70870 22334 70928 22380
rect 70974 22334 71000 22380
rect 70813 22276 71000 22334
rect 35784 22206 35826 22252
rect 35872 22206 35948 22252
rect 35784 22172 35948 22206
tri 35784 22022 35934 22172 ne
rect 35934 22126 35948 22172
tri 35948 22126 36074 22252 sw
rect 70813 22230 70824 22276
rect 70870 22230 70928 22276
rect 70974 22230 71000 22276
rect 70813 22172 71000 22230
rect 70813 22126 70824 22172
rect 70870 22126 70928 22172
rect 70974 22126 71000 22172
rect 35934 22120 36074 22126
rect 35934 22074 35958 22120
rect 36004 22074 36074 22120
rect 35934 22022 36074 22074
tri 35934 21892 36064 22022 ne
rect 36064 21988 36074 22022
tri 36074 21988 36212 22126 sw
rect 70813 22068 71000 22126
rect 70813 22022 70824 22068
rect 70870 22022 70928 22068
rect 70974 22022 71000 22068
rect 36064 21942 36090 21988
rect 36136 21942 36212 21988
rect 36064 21892 36212 21942
tri 36064 21756 36200 21892 ne
rect 36200 21860 36212 21892
tri 36212 21860 36340 21988 sw
rect 70813 21964 71000 22022
rect 70813 21918 70824 21964
rect 70870 21918 70928 21964
rect 70974 21918 71000 21964
rect 70813 21860 71000 21918
rect 36200 21856 36340 21860
rect 36200 21810 36222 21856
rect 36268 21810 36340 21856
rect 36200 21756 36340 21810
tri 36200 21648 36308 21756 ne
rect 36308 21724 36340 21756
tri 36340 21724 36476 21860 sw
rect 70813 21814 70824 21860
rect 70870 21814 70928 21860
rect 70974 21814 71000 21860
rect 70813 21756 71000 21814
rect 36308 21678 36354 21724
rect 36400 21678 36476 21724
rect 36308 21648 36476 21678
tri 36308 21502 36454 21648 ne
rect 36454 21606 36476 21648
tri 36476 21606 36594 21724 sw
rect 70813 21710 70824 21756
rect 70870 21710 70928 21756
rect 70974 21710 71000 21756
rect 70813 21652 71000 21710
rect 70813 21606 70824 21652
rect 70870 21606 70928 21652
rect 70974 21606 71000 21652
rect 36454 21592 36594 21606
rect 36454 21546 36486 21592
rect 36532 21546 36594 21592
rect 36454 21502 36594 21546
tri 36454 21398 36558 21502 ne
rect 36558 21460 36594 21502
tri 36594 21460 36740 21606 sw
rect 70813 21548 71000 21606
rect 70813 21502 70824 21548
rect 70870 21502 70928 21548
rect 70974 21502 71000 21548
rect 36558 21414 36618 21460
rect 36664 21414 36740 21460
rect 36558 21398 36740 21414
tri 36558 21236 36720 21398 ne
rect 36720 21340 36740 21398
tri 36740 21340 36860 21460 sw
rect 70813 21444 71000 21502
rect 70813 21398 70824 21444
rect 70870 21398 70928 21444
rect 70974 21398 71000 21444
rect 70813 21340 71000 21398
rect 36720 21328 36860 21340
rect 36720 21282 36750 21328
rect 36796 21282 36860 21328
rect 36720 21236 36860 21282
tri 36720 21132 36824 21236 ne
rect 36824 21196 36860 21236
tri 36860 21196 37004 21340 sw
rect 70813 21294 70824 21340
rect 70870 21294 70928 21340
rect 70974 21294 71000 21340
rect 70813 21236 71000 21294
rect 36824 21150 36882 21196
rect 36928 21150 37004 21196
rect 36824 21132 37004 21150
tri 36824 20982 36974 21132 ne
rect 36974 21064 37004 21132
tri 37004 21064 37136 21196 sw
rect 70813 21190 70824 21236
rect 70870 21190 70928 21236
rect 70974 21190 71000 21236
rect 70813 21132 71000 21190
rect 70813 21086 70824 21132
rect 70870 21086 70928 21132
rect 70974 21086 71000 21132
rect 36974 21018 37014 21064
rect 37060 21018 37136 21064
rect 36974 20982 37136 21018
tri 36974 20820 37136 20982 ne
tri 37136 20932 37268 21064 sw
rect 70813 21028 71000 21086
rect 70813 20982 70824 21028
rect 70870 20982 70928 21028
rect 70974 20982 71000 21028
rect 37136 20886 37146 20932
rect 37192 20886 37268 20932
rect 37136 20820 37268 20886
tri 37136 20716 37240 20820 ne
rect 37240 20800 37268 20820
tri 37268 20800 37400 20932 sw
rect 70813 20924 71000 20982
rect 70813 20878 70824 20924
rect 70870 20878 70928 20924
rect 70974 20878 71000 20924
rect 70813 20820 71000 20878
rect 37240 20754 37278 20800
rect 37324 20754 37400 20800
rect 37240 20716 37400 20754
tri 37240 20566 37390 20716 ne
rect 37390 20670 37400 20716
tri 37400 20670 37530 20800 sw
rect 70813 20774 70824 20820
rect 70870 20774 70928 20820
rect 70974 20774 71000 20820
rect 70813 20716 71000 20774
rect 70813 20670 70824 20716
rect 70870 20670 70928 20716
rect 70974 20670 71000 20716
rect 37390 20668 37530 20670
rect 37390 20622 37410 20668
rect 37456 20622 37530 20668
rect 37390 20566 37530 20622
tri 37390 20428 37528 20566 ne
rect 37528 20536 37530 20566
tri 37530 20536 37664 20670 sw
rect 70813 20612 71000 20670
rect 70813 20566 70824 20612
rect 70870 20566 70928 20612
rect 70974 20566 71000 20612
rect 37528 20490 37542 20536
rect 37588 20490 37664 20536
rect 37528 20428 37664 20490
tri 37528 20300 37656 20428 ne
rect 37656 20404 37664 20428
tri 37664 20404 37796 20536 sw
rect 70813 20508 71000 20566
rect 70813 20462 70824 20508
rect 70870 20462 70928 20508
rect 70974 20462 71000 20508
rect 70813 20404 71000 20462
rect 37656 20358 37674 20404
rect 37720 20358 37796 20404
rect 37656 20300 37796 20358
tri 37656 20184 37772 20300 ne
rect 37772 20272 37796 20300
tri 37796 20272 37928 20404 sw
rect 70813 20358 70824 20404
rect 70870 20358 70928 20404
rect 70974 20358 71000 20404
rect 70813 20300 71000 20358
rect 37772 20226 37806 20272
rect 37852 20226 37928 20272
rect 37772 20184 37928 20226
tri 37772 20046 37910 20184 ne
rect 37910 20150 37928 20184
tri 37928 20150 38050 20272 sw
rect 70813 20254 70824 20300
rect 70870 20254 70928 20300
rect 70974 20254 71000 20300
rect 70813 20196 71000 20254
rect 70813 20150 70824 20196
rect 70870 20150 70928 20196
rect 70974 20150 71000 20196
rect 37910 20140 38050 20150
rect 37910 20094 37938 20140
rect 37984 20094 38050 20140
rect 37910 20046 38050 20094
tri 37910 19940 38016 20046 ne
rect 38016 20008 38050 20046
tri 38050 20008 38192 20150 sw
rect 70813 20092 71000 20150
rect 70813 20046 70824 20092
rect 70870 20046 70928 20092
rect 70974 20046 71000 20092
rect 38016 19962 38070 20008
rect 38116 19962 38192 20008
rect 38016 19940 38192 19962
tri 38016 19780 38176 19940 ne
rect 38176 19884 38192 19940
tri 38192 19884 38316 20008 sw
rect 70813 19988 71000 20046
rect 70813 19942 70824 19988
rect 70870 19942 70928 19988
rect 70974 19942 71000 19988
rect 70813 19884 71000 19942
rect 38176 19876 38316 19884
rect 38176 19830 38202 19876
rect 38248 19830 38316 19876
rect 38176 19780 38316 19830
tri 38176 19676 38280 19780 ne
rect 38280 19744 38316 19780
tri 38316 19744 38456 19884 sw
rect 70813 19838 70824 19884
rect 70870 19838 70928 19884
rect 70974 19838 71000 19884
rect 70813 19780 71000 19838
rect 38280 19698 38334 19744
rect 38380 19698 38456 19744
rect 38280 19676 38456 19698
tri 38280 19526 38430 19676 ne
rect 38430 19612 38456 19676
tri 38456 19612 38588 19744 sw
rect 70813 19734 70824 19780
rect 70870 19734 70928 19780
rect 70974 19734 71000 19780
rect 70813 19676 71000 19734
rect 70813 19630 70824 19676
rect 70870 19630 70928 19676
rect 70974 19630 71000 19676
rect 38430 19566 38466 19612
rect 38512 19566 38588 19612
rect 38430 19526 38588 19566
tri 38430 19422 38534 19526 ne
rect 38534 19480 38588 19526
tri 38588 19480 38720 19612 sw
rect 70813 19572 71000 19630
rect 70813 19526 70824 19572
rect 70870 19526 70928 19572
rect 70974 19526 71000 19572
rect 38534 19434 38598 19480
rect 38644 19434 38720 19480
rect 38534 19422 38720 19434
tri 38534 19260 38696 19422 ne
rect 38696 19348 38720 19422
tri 38720 19348 38852 19480 sw
rect 70813 19468 71000 19526
rect 70813 19422 70824 19468
rect 70870 19422 70928 19468
rect 70974 19422 71000 19468
rect 70813 19364 71000 19422
rect 38696 19302 38730 19348
rect 38776 19302 38852 19348
rect 38696 19260 38852 19302
tri 38696 19110 38846 19260 ne
rect 38846 19216 38852 19260
tri 38852 19216 38984 19348 sw
rect 70813 19318 70824 19364
rect 70870 19318 70928 19364
rect 70974 19318 71000 19364
rect 70813 19260 71000 19318
rect 38846 19170 38862 19216
rect 38908 19170 38984 19216
rect 38846 19110 38984 19170
tri 38846 19006 38950 19110 ne
rect 38950 19084 38984 19110
tri 38984 19084 39116 19216 sw
rect 70813 19214 70824 19260
rect 70870 19214 70928 19260
rect 70974 19214 71000 19260
rect 70813 19156 71000 19214
rect 70813 19110 70824 19156
rect 70870 19110 70928 19156
rect 70974 19110 71000 19156
rect 38950 19038 38994 19084
rect 39040 19038 39116 19084
rect 38950 19006 39116 19038
tri 38950 18844 39112 19006 ne
rect 39112 18964 39116 19006
tri 39116 18964 39236 19084 sw
rect 70813 19052 71000 19110
rect 70813 19006 70824 19052
rect 70870 19006 70928 19052
rect 70974 19006 71000 19052
rect 39112 18952 39236 18964
rect 39112 18906 39126 18952
rect 39172 18906 39236 18952
rect 39112 18844 39236 18906
tri 39112 18720 39236 18844 ne
tri 39236 18820 39380 18964 sw
rect 70813 18948 71000 19006
rect 70813 18902 70824 18948
rect 70870 18902 70928 18948
rect 70974 18902 71000 18948
rect 70813 18844 71000 18902
rect 39236 18774 39258 18820
rect 39304 18774 39380 18820
rect 39236 18720 39380 18774
tri 39236 18590 39366 18720 ne
rect 39366 18694 39380 18720
tri 39380 18694 39506 18820 sw
rect 70813 18798 70824 18844
rect 70870 18798 70928 18844
rect 70974 18798 71000 18844
rect 70813 18740 71000 18798
rect 70813 18694 70824 18740
rect 70870 18694 70928 18740
rect 70974 18694 71000 18740
rect 39366 18688 39506 18694
rect 39366 18642 39390 18688
rect 39436 18642 39506 18688
rect 39366 18590 39506 18642
tri 39366 18476 39480 18590 ne
rect 39480 18556 39506 18590
tri 39506 18556 39644 18694 sw
rect 70813 18636 71000 18694
rect 70813 18590 70824 18636
rect 70870 18590 70928 18636
rect 70974 18590 71000 18636
rect 39480 18510 39522 18556
rect 39568 18510 39644 18556
rect 39480 18476 39644 18510
tri 39480 18324 39632 18476 ne
rect 39632 18428 39644 18476
tri 39644 18428 39772 18556 sw
rect 70813 18532 71000 18590
rect 70813 18486 70824 18532
rect 70870 18486 70928 18532
rect 70974 18486 71000 18532
rect 70813 18428 71000 18486
rect 39632 18424 39772 18428
rect 39632 18378 39654 18424
rect 39700 18378 39772 18424
rect 39632 18324 39772 18378
tri 39632 18220 39736 18324 ne
rect 39736 18292 39772 18324
tri 39772 18292 39908 18428 sw
rect 70813 18382 70824 18428
rect 70870 18382 70928 18428
rect 70974 18382 71000 18428
rect 70813 18324 71000 18382
rect 39736 18246 39786 18292
rect 39832 18246 39908 18292
rect 39736 18220 39908 18246
tri 39736 18070 39886 18220 ne
rect 39886 18174 39908 18220
tri 39908 18174 40026 18292 sw
rect 70813 18278 70824 18324
rect 70870 18278 70928 18324
rect 70974 18278 71000 18324
rect 70813 18220 71000 18278
rect 70813 18174 70824 18220
rect 70870 18174 70928 18220
rect 70974 18174 71000 18220
rect 39886 18160 40026 18174
rect 39886 18114 39918 18160
rect 39964 18114 40026 18160
rect 39886 18070 40026 18114
tri 39886 17966 39990 18070 ne
rect 39990 18028 40026 18070
tri 40026 18028 40172 18174 sw
rect 70813 18116 71000 18174
rect 70813 18070 70824 18116
rect 70870 18070 70928 18116
rect 70974 18070 71000 18116
rect 39990 17982 40050 18028
rect 40096 17982 40172 18028
rect 39990 17966 40172 17982
tri 39990 17804 40152 17966 ne
rect 40152 17896 40172 17966
tri 40172 17896 40304 18028 sw
rect 70813 18012 71000 18070
rect 70813 17966 70824 18012
rect 70870 17966 70928 18012
rect 70974 17966 71000 18012
rect 70813 17908 71000 17966
rect 40152 17850 40182 17896
rect 40228 17850 40304 17896
rect 40152 17804 40304 17850
tri 40152 17654 40302 17804 ne
rect 40302 17764 40304 17804
tri 40304 17764 40436 17896 sw
rect 70813 17862 70824 17908
rect 70870 17862 70928 17908
rect 70974 17862 71000 17908
rect 70813 17804 71000 17862
rect 40302 17718 40314 17764
rect 40360 17718 40436 17764
rect 40302 17654 40436 17718
tri 40302 17550 40406 17654 ne
rect 40406 17632 40436 17654
tri 40436 17632 40568 17764 sw
rect 70813 17758 70824 17804
rect 70870 17758 70928 17804
rect 70974 17758 71000 17804
rect 70813 17700 71000 17758
rect 70813 17654 70824 17700
rect 70870 17654 70928 17700
rect 70974 17654 71000 17700
rect 40406 17586 40446 17632
rect 40492 17586 40568 17632
rect 40406 17550 40568 17586
tri 40406 17388 40568 17550 ne
tri 40568 17500 40700 17632 sw
rect 70813 17596 71000 17654
rect 70813 17550 70824 17596
rect 70870 17550 70928 17596
rect 70974 17550 71000 17596
rect 40568 17454 40578 17500
rect 40624 17454 40700 17500
rect 40568 17388 40700 17454
tri 40568 17256 40700 17388 ne
tri 40700 17368 40832 17500 sw
rect 70813 17492 71000 17550
rect 70813 17446 70824 17492
rect 70870 17446 70928 17492
rect 70974 17446 71000 17492
rect 70813 17388 71000 17446
rect 40700 17322 40710 17368
rect 40756 17322 40832 17368
rect 40700 17256 40832 17322
tri 40700 17134 40822 17256 ne
rect 40822 17238 40832 17256
tri 40832 17238 40962 17368 sw
rect 70813 17342 70824 17388
rect 70870 17342 70928 17388
rect 70974 17342 71000 17388
rect 70813 17284 71000 17342
rect 70813 17238 70824 17284
rect 70870 17238 70928 17284
rect 70974 17238 71000 17284
rect 40822 17236 40962 17238
rect 40822 17190 40842 17236
rect 40888 17190 40962 17236
rect 40822 17134 40962 17190
tri 40822 17012 40944 17134 ne
rect 40944 17104 40962 17134
tri 40962 17104 41096 17238 sw
rect 70813 17180 71000 17238
rect 70813 17134 70824 17180
rect 70870 17134 70928 17180
rect 70974 17134 71000 17180
rect 40944 17058 40974 17104
rect 41020 17058 41096 17104
rect 40944 17012 41096 17058
tri 40944 16868 41088 17012 ne
rect 41088 16972 41096 17012
tri 41096 16972 41228 17104 sw
rect 70813 17076 71000 17134
rect 70813 17030 70824 17076
rect 70870 17030 70928 17076
rect 70974 17030 71000 17076
rect 70813 16972 71000 17030
rect 41088 16926 41106 16972
rect 41152 16926 41228 16972
rect 41088 16868 41228 16926
tri 41088 16764 41192 16868 ne
rect 41192 16840 41228 16868
tri 41228 16840 41360 16972 sw
rect 70813 16926 70824 16972
rect 70870 16926 70928 16972
rect 70974 16926 71000 16972
rect 70813 16868 71000 16926
rect 41192 16794 41238 16840
rect 41284 16794 41360 16840
rect 41192 16764 41360 16794
tri 41192 16614 41342 16764 ne
rect 41342 16718 41360 16764
tri 41360 16718 41482 16840 sw
rect 70813 16822 70824 16868
rect 70870 16822 70928 16868
rect 70974 16822 71000 16868
rect 70813 16764 71000 16822
rect 70813 16718 70824 16764
rect 70870 16718 70928 16764
rect 70974 16718 71000 16764
rect 41342 16708 41482 16718
rect 41342 16662 41370 16708
rect 41416 16662 41482 16708
rect 41342 16614 41482 16662
tri 41342 16510 41446 16614 ne
rect 41446 16576 41482 16614
tri 41482 16576 41624 16718 sw
rect 70813 16660 71000 16718
rect 70813 16614 70824 16660
rect 70870 16614 70928 16660
rect 70974 16614 71000 16660
rect 41446 16530 41502 16576
rect 41548 16530 41624 16576
rect 41446 16510 41624 16530
tri 41446 16348 41608 16510 ne
rect 41608 16444 41624 16510
tri 41624 16444 41756 16576 sw
rect 70813 16556 71000 16614
rect 70813 16510 70824 16556
rect 70870 16510 70928 16556
rect 70974 16510 71000 16556
rect 70813 16452 71000 16510
rect 41608 16398 41634 16444
rect 41680 16398 41756 16444
rect 41608 16348 41756 16398
tri 41608 16244 41712 16348 ne
rect 41712 16312 41756 16348
tri 41756 16312 41888 16444 sw
rect 70813 16406 70824 16452
rect 70870 16406 70928 16452
rect 70974 16406 71000 16452
rect 70813 16348 71000 16406
rect 41712 16266 41766 16312
rect 41812 16266 41888 16312
rect 41712 16244 41888 16266
tri 41712 16094 41862 16244 ne
rect 41862 16180 41888 16244
tri 41888 16180 42020 16312 sw
rect 70813 16302 70824 16348
rect 70870 16302 70928 16348
rect 70974 16302 71000 16348
rect 70813 16244 71000 16302
rect 70813 16198 70824 16244
rect 70870 16198 70928 16244
rect 70974 16198 71000 16244
rect 41862 16134 41898 16180
rect 41944 16134 42020 16180
rect 41862 16094 42020 16134
tri 41862 15990 41966 16094 ne
rect 41966 16048 42020 16094
tri 42020 16048 42152 16180 sw
rect 70813 16140 71000 16198
rect 70813 16094 70824 16140
rect 70870 16094 70928 16140
rect 70974 16094 71000 16140
rect 41966 16002 42030 16048
rect 42076 16002 42152 16048
rect 41966 15990 42152 16002
tri 41966 15828 42128 15990 ne
rect 42128 15916 42152 15990
tri 42152 15916 42284 16048 sw
rect 70813 16036 71000 16094
rect 70813 15990 70824 16036
rect 70870 15990 70928 16036
rect 70974 15990 71000 16036
rect 70813 15932 71000 15990
rect 42128 15870 42162 15916
rect 42208 15870 42284 15916
rect 42128 15828 42284 15870
tri 42128 15678 42278 15828 ne
rect 42278 15792 42284 15828
tri 42284 15792 42408 15916 sw
rect 70813 15886 70824 15932
rect 70870 15886 70928 15932
rect 70974 15886 71000 15932
rect 70813 15828 71000 15886
rect 42278 15784 42408 15792
rect 42278 15738 42294 15784
rect 42340 15738 42408 15784
rect 42278 15678 42408 15738
tri 42278 15548 42408 15678 ne
tri 42408 15652 42548 15792 sw
rect 70813 15782 70824 15828
rect 70870 15782 70928 15828
rect 70974 15782 71000 15828
rect 70813 15724 71000 15782
rect 70813 15678 70824 15724
rect 70870 15678 70928 15724
rect 70974 15678 71000 15724
rect 42408 15606 42426 15652
rect 42472 15606 42548 15652
rect 42408 15548 42548 15606
tri 42548 15548 42652 15652 sw
rect 70813 15620 71000 15678
rect 70813 15574 70824 15620
rect 70870 15574 70928 15620
rect 70974 15574 71000 15620
tri 42408 15412 42544 15548 ne
rect 42544 15520 42652 15548
rect 42544 15474 42558 15520
rect 42604 15474 42652 15520
rect 42544 15412 42652 15474
tri 42544 15304 42652 15412 ne
tri 42652 15388 42812 15548 sw
rect 70813 15516 71000 15574
rect 70813 15470 70824 15516
rect 70870 15470 70928 15516
rect 70974 15470 71000 15516
rect 70813 15412 71000 15470
rect 42652 15342 42690 15388
rect 42736 15342 42812 15388
rect 42652 15304 42812 15342
tri 42652 15158 42798 15304 ne
rect 42798 15262 42812 15304
tri 42812 15262 42938 15388 sw
rect 70813 15366 70824 15412
rect 70870 15366 70928 15412
rect 70974 15366 71000 15412
rect 70813 15308 71000 15366
rect 70813 15262 70824 15308
rect 70870 15262 70928 15308
rect 70974 15262 71000 15308
rect 42798 15256 42938 15262
rect 42798 15210 42822 15256
rect 42868 15210 42938 15256
rect 42798 15158 42938 15210
tri 42798 15054 42902 15158 ne
rect 42902 15124 42938 15158
tri 42938 15124 43076 15262 sw
rect 70813 15204 71000 15262
rect 70813 15158 70824 15204
rect 70870 15158 70928 15204
rect 70974 15158 71000 15204
rect 42902 15078 42954 15124
rect 43000 15078 43076 15124
rect 42902 15054 43076 15078
tri 42902 14892 43064 15054 ne
rect 43064 14996 43076 15054
tri 43076 14996 43204 15124 sw
rect 70813 15100 71000 15158
rect 70813 15054 70824 15100
rect 70870 15054 70928 15100
rect 70974 15054 71000 15100
rect 70813 14996 71000 15054
rect 43064 14992 43204 14996
rect 43064 14946 43086 14992
rect 43132 14946 43204 14992
rect 43064 14892 43204 14946
tri 43064 14788 43168 14892 ne
rect 43168 14860 43204 14892
tri 43204 14860 43340 14996 sw
rect 70813 14950 70824 14996
rect 70870 14950 70928 14996
rect 70974 14950 71000 14996
rect 70813 14892 71000 14950
rect 43168 14814 43218 14860
rect 43264 14814 43340 14860
rect 43168 14788 43340 14814
tri 43168 14638 43318 14788 ne
rect 43318 14728 43340 14788
tri 43340 14728 43472 14860 sw
rect 70813 14846 70824 14892
rect 70870 14846 70928 14892
rect 70974 14846 71000 14892
rect 70813 14788 71000 14846
rect 70813 14742 70824 14788
rect 70870 14742 70928 14788
rect 70974 14742 71000 14788
rect 43318 14682 43350 14728
rect 43396 14682 43472 14728
rect 43318 14638 43472 14682
tri 43318 14534 43422 14638 ne
rect 43422 14596 43472 14638
tri 43472 14596 43604 14728 sw
rect 70813 14684 71000 14742
rect 70813 14638 70824 14684
rect 70870 14638 70928 14684
rect 70974 14638 71000 14684
rect 43422 14550 43482 14596
rect 43528 14550 43604 14596
rect 43422 14534 43604 14550
tri 43422 14372 43584 14534 ne
rect 43584 14464 43604 14534
tri 43604 14464 43736 14596 sw
rect 70813 14580 71000 14638
rect 70813 14534 70824 14580
rect 70870 14534 70928 14580
rect 70974 14534 71000 14580
rect 70813 14476 71000 14534
rect 43584 14418 43614 14464
rect 43660 14418 43736 14464
rect 43584 14372 43736 14418
tri 43584 14222 43734 14372 ne
rect 43734 14332 43736 14372
tri 43736 14332 43868 14464 sw
rect 70813 14430 70824 14476
rect 70870 14430 70928 14476
rect 70974 14430 71000 14476
rect 70813 14372 71000 14430
rect 43734 14286 43746 14332
rect 43792 14286 43868 14332
rect 43734 14222 43868 14286
tri 43734 14118 43838 14222 ne
rect 43838 14200 43868 14222
tri 43868 14200 44000 14332 sw
rect 70813 14326 70824 14372
rect 70870 14326 70928 14372
rect 70974 14326 71000 14372
rect 70813 14268 71000 14326
rect 70813 14222 70824 14268
rect 70870 14222 70928 14268
rect 70974 14222 71000 14268
rect 43838 14154 43878 14200
rect 43924 14154 44000 14200
rect 43838 14118 44000 14154
tri 43838 13956 44000 14118 ne
tri 44000 14084 44116 14200 sw
rect 70813 14164 71000 14222
rect 70813 14118 70824 14164
rect 70870 14118 70928 14164
rect 70974 14118 71000 14164
rect 44000 14068 44116 14084
rect 44000 14022 44010 14068
rect 44056 14022 44116 14068
rect 44000 13956 44116 14022
tri 44000 13840 44116 13956 ne
tri 44116 13936 44264 14084 sw
rect 70813 14060 71000 14118
rect 70813 14014 70824 14060
rect 70870 14014 70928 14060
rect 70974 14014 71000 14060
rect 70813 13956 71000 14014
rect 44116 13890 44142 13936
rect 44188 13890 44264 13936
rect 44116 13840 44264 13890
tri 44116 13702 44254 13840 ne
rect 44254 13806 44264 13840
tri 44264 13806 44394 13936 sw
rect 70813 13910 70824 13956
rect 70870 13910 70928 13956
rect 70974 13910 71000 13956
rect 70813 13852 71000 13910
rect 70813 13806 70824 13852
rect 70870 13806 70928 13852
rect 70974 13806 71000 13852
rect 44254 13804 44394 13806
rect 44254 13758 44274 13804
rect 44320 13758 44394 13804
rect 44254 13702 44394 13758
tri 44254 13596 44360 13702 ne
rect 44360 13672 44394 13702
tri 44394 13672 44528 13806 sw
rect 70813 13748 71000 13806
rect 70813 13702 70824 13748
rect 70870 13702 70928 13748
rect 70974 13702 71000 13748
rect 44360 13626 44406 13672
rect 44452 13626 44528 13672
rect 44360 13596 44528 13626
tri 44360 13436 44520 13596 ne
rect 44520 13540 44528 13596
tri 44528 13540 44660 13672 sw
rect 70813 13644 71000 13702
rect 70813 13598 70824 13644
rect 70870 13598 70928 13644
rect 70974 13598 71000 13644
rect 70813 13540 71000 13598
rect 44520 13494 44538 13540
rect 44584 13494 44660 13540
rect 44520 13436 44660 13494
tri 44520 13352 44604 13436 ne
rect 44604 13408 44660 13436
tri 44660 13408 44792 13540 sw
rect 70813 13494 70824 13540
rect 70870 13494 70928 13540
rect 70974 13494 71000 13540
rect 70813 13436 71000 13494
rect 44604 13362 44670 13408
rect 44716 13362 44792 13408
rect 44604 13352 44792 13362
tri 44604 13165 44791 13352 ne
rect 44791 13280 44792 13352
tri 44792 13280 44920 13408 sw
rect 70813 13390 70824 13436
rect 70870 13390 70928 13436
rect 70974 13390 71000 13436
rect 70813 13280 71000 13390
rect 44791 13269 71000 13280
rect 44791 13256 45088 13269
rect 44791 13210 44850 13256
rect 44896 13223 45088 13256
rect 45134 13223 45192 13269
rect 45238 13223 45296 13269
rect 45342 13223 45400 13269
rect 45446 13223 45504 13269
rect 45550 13223 45608 13269
rect 45654 13223 45712 13269
rect 45758 13223 45816 13269
rect 45862 13223 45920 13269
rect 45966 13223 46024 13269
rect 46070 13223 46128 13269
rect 46174 13223 46232 13269
rect 46278 13223 46336 13269
rect 46382 13223 46440 13269
rect 46486 13223 46544 13269
rect 46590 13223 46648 13269
rect 46694 13223 46752 13269
rect 46798 13223 46856 13269
rect 46902 13223 46960 13269
rect 47006 13223 47064 13269
rect 47110 13223 47168 13269
rect 47214 13223 47272 13269
rect 47318 13223 47376 13269
rect 47422 13223 47480 13269
rect 47526 13223 47584 13269
rect 47630 13223 47688 13269
rect 47734 13223 47792 13269
rect 47838 13223 47896 13269
rect 47942 13223 48000 13269
rect 48046 13223 48104 13269
rect 48150 13223 48208 13269
rect 48254 13223 48312 13269
rect 48358 13223 48416 13269
rect 48462 13223 48520 13269
rect 48566 13223 48624 13269
rect 48670 13223 48728 13269
rect 48774 13223 48832 13269
rect 48878 13223 48936 13269
rect 48982 13223 49040 13269
rect 49086 13223 49144 13269
rect 49190 13223 49248 13269
rect 49294 13223 49352 13269
rect 49398 13223 49456 13269
rect 49502 13223 49560 13269
rect 49606 13223 49664 13269
rect 49710 13223 49768 13269
rect 49814 13223 49872 13269
rect 49918 13223 49976 13269
rect 50022 13223 50080 13269
rect 50126 13223 50184 13269
rect 50230 13223 50288 13269
rect 50334 13223 50392 13269
rect 50438 13223 50496 13269
rect 50542 13223 50600 13269
rect 50646 13223 50704 13269
rect 50750 13223 50808 13269
rect 50854 13223 50912 13269
rect 50958 13223 51016 13269
rect 51062 13223 51120 13269
rect 51166 13223 51224 13269
rect 51270 13223 51328 13269
rect 51374 13223 51432 13269
rect 51478 13223 51536 13269
rect 51582 13223 51640 13269
rect 51686 13223 51744 13269
rect 51790 13223 51848 13269
rect 51894 13223 51952 13269
rect 51998 13223 52056 13269
rect 52102 13223 52160 13269
rect 52206 13223 52264 13269
rect 52310 13223 52368 13269
rect 52414 13223 52472 13269
rect 52518 13223 52576 13269
rect 52622 13223 52680 13269
rect 52726 13223 52784 13269
rect 52830 13223 52888 13269
rect 52934 13223 52992 13269
rect 53038 13223 53096 13269
rect 53142 13223 53200 13269
rect 53246 13223 53304 13269
rect 53350 13223 53408 13269
rect 53454 13223 53512 13269
rect 53558 13223 53616 13269
rect 53662 13223 53720 13269
rect 53766 13223 53824 13269
rect 53870 13223 53928 13269
rect 53974 13223 54032 13269
rect 54078 13223 54136 13269
rect 54182 13223 54240 13269
rect 54286 13223 54344 13269
rect 54390 13223 54448 13269
rect 54494 13223 54552 13269
rect 54598 13223 54656 13269
rect 54702 13223 54760 13269
rect 54806 13223 54864 13269
rect 54910 13223 54968 13269
rect 55014 13223 55072 13269
rect 55118 13223 55176 13269
rect 55222 13223 55280 13269
rect 55326 13223 55384 13269
rect 55430 13223 55488 13269
rect 55534 13223 55592 13269
rect 55638 13223 55696 13269
rect 55742 13223 55800 13269
rect 55846 13223 55904 13269
rect 55950 13223 56008 13269
rect 56054 13223 56112 13269
rect 56158 13223 56216 13269
rect 56262 13223 56320 13269
rect 56366 13223 56424 13269
rect 56470 13223 56528 13269
rect 56574 13223 56632 13269
rect 56678 13223 56736 13269
rect 56782 13223 56840 13269
rect 56886 13223 56944 13269
rect 56990 13223 57048 13269
rect 57094 13223 57152 13269
rect 57198 13223 57256 13269
rect 57302 13223 57360 13269
rect 57406 13223 57464 13269
rect 57510 13223 57568 13269
rect 57614 13223 57672 13269
rect 57718 13223 57776 13269
rect 57822 13223 57880 13269
rect 57926 13223 57984 13269
rect 58030 13223 58088 13269
rect 58134 13223 58192 13269
rect 58238 13223 58296 13269
rect 58342 13223 58400 13269
rect 58446 13223 58504 13269
rect 58550 13223 58608 13269
rect 58654 13223 58712 13269
rect 58758 13223 58816 13269
rect 58862 13223 58920 13269
rect 58966 13223 59024 13269
rect 59070 13223 59128 13269
rect 59174 13223 59232 13269
rect 59278 13223 59336 13269
rect 59382 13223 59440 13269
rect 59486 13223 59544 13269
rect 59590 13223 59648 13269
rect 59694 13223 59752 13269
rect 59798 13223 59856 13269
rect 59902 13223 59960 13269
rect 60006 13223 60064 13269
rect 60110 13223 60168 13269
rect 60214 13223 60272 13269
rect 60318 13223 60376 13269
rect 60422 13223 60480 13269
rect 60526 13223 60584 13269
rect 60630 13223 60688 13269
rect 60734 13223 60792 13269
rect 60838 13223 60896 13269
rect 60942 13223 61000 13269
rect 61046 13223 61104 13269
rect 61150 13223 61208 13269
rect 61254 13223 61312 13269
rect 61358 13223 61416 13269
rect 61462 13223 61520 13269
rect 61566 13223 61624 13269
rect 61670 13223 61728 13269
rect 61774 13223 61832 13269
rect 61878 13223 61936 13269
rect 61982 13223 62040 13269
rect 62086 13223 62144 13269
rect 62190 13223 62248 13269
rect 62294 13223 62352 13269
rect 62398 13223 62456 13269
rect 62502 13223 62560 13269
rect 62606 13223 62664 13269
rect 62710 13223 62768 13269
rect 62814 13223 62872 13269
rect 62918 13223 62976 13269
rect 63022 13223 63080 13269
rect 63126 13223 63184 13269
rect 63230 13223 63288 13269
rect 63334 13223 63392 13269
rect 63438 13223 63496 13269
rect 63542 13223 63600 13269
rect 63646 13223 63704 13269
rect 63750 13223 63808 13269
rect 63854 13223 63912 13269
rect 63958 13223 64016 13269
rect 64062 13223 64120 13269
rect 64166 13223 64224 13269
rect 64270 13223 64328 13269
rect 64374 13223 64432 13269
rect 64478 13223 64536 13269
rect 64582 13223 64640 13269
rect 64686 13223 64744 13269
rect 64790 13223 64848 13269
rect 64894 13223 64952 13269
rect 64998 13223 65056 13269
rect 65102 13223 65160 13269
rect 65206 13223 65264 13269
rect 65310 13223 65368 13269
rect 65414 13223 65472 13269
rect 65518 13223 65576 13269
rect 65622 13223 65680 13269
rect 65726 13223 65784 13269
rect 65830 13223 65888 13269
rect 65934 13223 65992 13269
rect 66038 13223 66096 13269
rect 66142 13223 66200 13269
rect 66246 13223 66304 13269
rect 66350 13223 66408 13269
rect 66454 13223 66512 13269
rect 66558 13223 66616 13269
rect 66662 13223 66720 13269
rect 66766 13223 66824 13269
rect 66870 13223 66928 13269
rect 66974 13223 67032 13269
rect 67078 13223 67136 13269
rect 67182 13223 67240 13269
rect 67286 13223 67344 13269
rect 67390 13223 67448 13269
rect 67494 13223 67552 13269
rect 67598 13223 67656 13269
rect 67702 13223 67760 13269
rect 67806 13223 67864 13269
rect 67910 13223 67968 13269
rect 68014 13223 68072 13269
rect 68118 13223 68176 13269
rect 68222 13223 68280 13269
rect 68326 13223 68384 13269
rect 68430 13223 68488 13269
rect 68534 13223 68592 13269
rect 68638 13223 68696 13269
rect 68742 13223 68800 13269
rect 68846 13223 68904 13269
rect 68950 13223 69008 13269
rect 69054 13223 69112 13269
rect 69158 13223 69216 13269
rect 69262 13223 69320 13269
rect 69366 13223 69424 13269
rect 69470 13223 69528 13269
rect 69574 13223 69632 13269
rect 69678 13223 69736 13269
rect 69782 13223 69840 13269
rect 69886 13223 69944 13269
rect 69990 13223 70048 13269
rect 70094 13223 70152 13269
rect 70198 13223 70256 13269
rect 70302 13223 70360 13269
rect 70406 13223 70464 13269
rect 70510 13223 70568 13269
rect 70614 13223 70672 13269
rect 70718 13223 70776 13269
rect 70822 13223 70880 13269
rect 70926 13223 71000 13269
rect 44896 13210 71000 13223
rect 44791 13165 71000 13210
tri 44791 13108 44848 13165 ne
rect 44848 13119 45088 13165
rect 45134 13119 45192 13165
rect 45238 13119 45296 13165
rect 45342 13119 45400 13165
rect 45446 13119 45504 13165
rect 45550 13119 45608 13165
rect 45654 13119 45712 13165
rect 45758 13119 45816 13165
rect 45862 13119 45920 13165
rect 45966 13119 46024 13165
rect 46070 13119 46128 13165
rect 46174 13119 46232 13165
rect 46278 13119 46336 13165
rect 46382 13119 46440 13165
rect 46486 13119 46544 13165
rect 46590 13119 46648 13165
rect 46694 13119 46752 13165
rect 46798 13119 46856 13165
rect 46902 13119 46960 13165
rect 47006 13119 47064 13165
rect 47110 13119 47168 13165
rect 47214 13119 47272 13165
rect 47318 13119 47376 13165
rect 47422 13119 47480 13165
rect 47526 13119 47584 13165
rect 47630 13119 47688 13165
rect 47734 13119 47792 13165
rect 47838 13119 47896 13165
rect 47942 13119 48000 13165
rect 48046 13119 48104 13165
rect 48150 13119 48208 13165
rect 48254 13119 48312 13165
rect 48358 13119 48416 13165
rect 48462 13119 48520 13165
rect 48566 13119 48624 13165
rect 48670 13119 48728 13165
rect 48774 13119 48832 13165
rect 48878 13119 48936 13165
rect 48982 13119 49040 13165
rect 49086 13119 49144 13165
rect 49190 13119 49248 13165
rect 49294 13119 49352 13165
rect 49398 13119 49456 13165
rect 49502 13119 49560 13165
rect 49606 13119 49664 13165
rect 49710 13119 49768 13165
rect 49814 13119 49872 13165
rect 49918 13119 49976 13165
rect 50022 13119 50080 13165
rect 50126 13119 50184 13165
rect 50230 13119 50288 13165
rect 50334 13119 50392 13165
rect 50438 13119 50496 13165
rect 50542 13119 50600 13165
rect 50646 13119 50704 13165
rect 50750 13119 50808 13165
rect 50854 13119 50912 13165
rect 50958 13119 51016 13165
rect 51062 13119 51120 13165
rect 51166 13119 51224 13165
rect 51270 13119 51328 13165
rect 51374 13119 51432 13165
rect 51478 13119 51536 13165
rect 51582 13119 51640 13165
rect 51686 13119 51744 13165
rect 51790 13119 51848 13165
rect 51894 13119 51952 13165
rect 51998 13119 52056 13165
rect 52102 13119 52160 13165
rect 52206 13119 52264 13165
rect 52310 13119 52368 13165
rect 52414 13119 52472 13165
rect 52518 13119 52576 13165
rect 52622 13119 52680 13165
rect 52726 13119 52784 13165
rect 52830 13119 52888 13165
rect 52934 13119 52992 13165
rect 53038 13119 53096 13165
rect 53142 13119 53200 13165
rect 53246 13119 53304 13165
rect 53350 13119 53408 13165
rect 53454 13119 53512 13165
rect 53558 13119 53616 13165
rect 53662 13119 53720 13165
rect 53766 13119 53824 13165
rect 53870 13119 53928 13165
rect 53974 13119 54032 13165
rect 54078 13119 54136 13165
rect 54182 13119 54240 13165
rect 54286 13119 54344 13165
rect 54390 13119 54448 13165
rect 54494 13119 54552 13165
rect 54598 13119 54656 13165
rect 54702 13119 54760 13165
rect 54806 13119 54864 13165
rect 54910 13119 54968 13165
rect 55014 13119 55072 13165
rect 55118 13119 55176 13165
rect 55222 13119 55280 13165
rect 55326 13119 55384 13165
rect 55430 13119 55488 13165
rect 55534 13119 55592 13165
rect 55638 13119 55696 13165
rect 55742 13119 55800 13165
rect 55846 13119 55904 13165
rect 55950 13119 56008 13165
rect 56054 13119 56112 13165
rect 56158 13119 56216 13165
rect 56262 13119 56320 13165
rect 56366 13119 56424 13165
rect 56470 13119 56528 13165
rect 56574 13119 56632 13165
rect 56678 13119 56736 13165
rect 56782 13119 56840 13165
rect 56886 13119 56944 13165
rect 56990 13119 57048 13165
rect 57094 13119 57152 13165
rect 57198 13119 57256 13165
rect 57302 13119 57360 13165
rect 57406 13119 57464 13165
rect 57510 13119 57568 13165
rect 57614 13119 57672 13165
rect 57718 13119 57776 13165
rect 57822 13119 57880 13165
rect 57926 13119 57984 13165
rect 58030 13119 58088 13165
rect 58134 13119 58192 13165
rect 58238 13119 58296 13165
rect 58342 13119 58400 13165
rect 58446 13119 58504 13165
rect 58550 13119 58608 13165
rect 58654 13119 58712 13165
rect 58758 13119 58816 13165
rect 58862 13119 58920 13165
rect 58966 13119 59024 13165
rect 59070 13119 59128 13165
rect 59174 13119 59232 13165
rect 59278 13119 59336 13165
rect 59382 13119 59440 13165
rect 59486 13119 59544 13165
rect 59590 13119 59648 13165
rect 59694 13119 59752 13165
rect 59798 13119 59856 13165
rect 59902 13119 59960 13165
rect 60006 13119 60064 13165
rect 60110 13119 60168 13165
rect 60214 13119 60272 13165
rect 60318 13119 60376 13165
rect 60422 13119 60480 13165
rect 60526 13119 60584 13165
rect 60630 13119 60688 13165
rect 60734 13119 60792 13165
rect 60838 13119 60896 13165
rect 60942 13119 61000 13165
rect 61046 13119 61104 13165
rect 61150 13119 61208 13165
rect 61254 13119 61312 13165
rect 61358 13119 61416 13165
rect 61462 13119 61520 13165
rect 61566 13119 61624 13165
rect 61670 13119 61728 13165
rect 61774 13119 61832 13165
rect 61878 13119 61936 13165
rect 61982 13119 62040 13165
rect 62086 13119 62144 13165
rect 62190 13119 62248 13165
rect 62294 13119 62352 13165
rect 62398 13119 62456 13165
rect 62502 13119 62560 13165
rect 62606 13119 62664 13165
rect 62710 13119 62768 13165
rect 62814 13119 62872 13165
rect 62918 13119 62976 13165
rect 63022 13119 63080 13165
rect 63126 13119 63184 13165
rect 63230 13119 63288 13165
rect 63334 13119 63392 13165
rect 63438 13119 63496 13165
rect 63542 13119 63600 13165
rect 63646 13119 63704 13165
rect 63750 13119 63808 13165
rect 63854 13119 63912 13165
rect 63958 13119 64016 13165
rect 64062 13119 64120 13165
rect 64166 13119 64224 13165
rect 64270 13119 64328 13165
rect 64374 13119 64432 13165
rect 64478 13119 64536 13165
rect 64582 13119 64640 13165
rect 64686 13119 64744 13165
rect 64790 13119 64848 13165
rect 64894 13119 64952 13165
rect 64998 13119 65056 13165
rect 65102 13119 65160 13165
rect 65206 13119 65264 13165
rect 65310 13119 65368 13165
rect 65414 13119 65472 13165
rect 65518 13119 65576 13165
rect 65622 13119 65680 13165
rect 65726 13119 65784 13165
rect 65830 13119 65888 13165
rect 65934 13119 65992 13165
rect 66038 13119 66096 13165
rect 66142 13119 66200 13165
rect 66246 13119 66304 13165
rect 66350 13119 66408 13165
rect 66454 13119 66512 13165
rect 66558 13119 66616 13165
rect 66662 13119 66720 13165
rect 66766 13119 66824 13165
rect 66870 13119 66928 13165
rect 66974 13119 67032 13165
rect 67078 13119 67136 13165
rect 67182 13119 67240 13165
rect 67286 13119 67344 13165
rect 67390 13119 67448 13165
rect 67494 13119 67552 13165
rect 67598 13119 67656 13165
rect 67702 13119 67760 13165
rect 67806 13119 67864 13165
rect 67910 13119 67968 13165
rect 68014 13119 68072 13165
rect 68118 13119 68176 13165
rect 68222 13119 68280 13165
rect 68326 13119 68384 13165
rect 68430 13119 68488 13165
rect 68534 13119 68592 13165
rect 68638 13119 68696 13165
rect 68742 13119 68800 13165
rect 68846 13119 68904 13165
rect 68950 13119 69008 13165
rect 69054 13119 69112 13165
rect 69158 13119 69216 13165
rect 69262 13119 69320 13165
rect 69366 13119 69424 13165
rect 69470 13119 69528 13165
rect 69574 13119 69632 13165
rect 69678 13119 69736 13165
rect 69782 13119 69840 13165
rect 69886 13119 69944 13165
rect 69990 13119 70048 13165
rect 70094 13119 70152 13165
rect 70198 13119 70256 13165
rect 70302 13119 70360 13165
rect 70406 13119 70464 13165
rect 70510 13119 70568 13165
rect 70614 13119 70672 13165
rect 70718 13119 70776 13165
rect 70822 13119 70880 13165
rect 70926 13119 71000 13165
rect 44848 13108 71000 13119
<< metal2 >>
rect 70584 68116 70702 68200
rect 70584 66916 70613 68116
rect 70669 66916 70702 68116
rect 70584 60120 70702 66916
rect 70584 58920 70613 60120
rect 70669 58920 70702 60120
rect 70584 56910 70702 58920
rect 70584 55710 70613 56910
rect 70669 55710 70702 56910
rect 70584 55302 70702 55710
rect 70584 54102 70613 55302
rect 70669 54102 70702 55302
rect 70584 53722 70702 54102
rect 70584 52522 70613 53722
rect 70669 52522 70702 53722
rect 70584 45739 70702 52522
rect 70584 42875 70613 45739
rect 70669 42875 70702 45739
rect 70584 42497 70702 42875
rect 70584 41297 70613 42497
rect 70669 41297 70702 42497
rect 70584 39332 70702 41297
rect 70584 36468 70613 39332
rect 70669 36468 70702 39332
rect 70584 36132 70702 36468
rect 70584 33268 70613 36132
rect 70669 33268 70702 36132
rect 70584 32920 70702 33268
rect 70584 30056 70613 32920
rect 70669 30056 70702 32920
rect 70584 29752 70702 30056
rect 70584 26888 70613 29752
rect 70669 26888 70702 29752
rect 70584 24906 70702 26888
rect 70584 23706 70613 24906
rect 70669 23706 70702 24906
rect 70584 23599 70702 23706
<< via2 >>
rect 70613 66916 70669 68116
rect 70613 58920 70669 60120
rect 70613 55710 70669 56910
rect 70613 54102 70669 55302
rect 70613 52522 70669 53722
rect 70613 42875 70669 45739
rect 70613 41297 70669 42497
rect 70613 36468 70669 39332
rect 70613 33268 70669 36132
rect 70613 30056 70669 32920
rect 70613 26888 70669 29752
rect 70613 23706 70669 24906
<< metal3 >>
rect 14000 47112 17000 71000
rect 17200 48448 20200 71000
rect 20400 49774 23400 71000
rect 23600 50451 25000 71000
rect 25200 51220 26600 71000
rect 26800 52454 29800 71000
rect 30000 53792 33000 71000
rect 33200 55124 36200 71000
rect 36400 56465 39400 71000
rect 39600 57138 41000 71000
rect 41200 57723 42600 71000
rect 42800 59150 45800 71000
rect 46000 60510 49000 71000
rect 49200 61175 50600 71000
rect 50800 61839 52200 71000
rect 52400 62507 53800 71000
rect 54000 63173 55400 71000
rect 55600 63836 57000 71000
rect 57200 64499 58600 71000
rect 58800 65166 60200 71000
rect 60400 65831 61800 71000
rect 62000 66494 63400 71000
rect 63600 67166 65000 71000
rect 65200 67829 66600 71000
rect 66800 68476 68200 71000
rect 68400 69678 69678 71000
rect 68400 68769 71000 69678
tri 68400 68693 68476 68769 ne
rect 68476 68693 71000 68769
tri 68200 68476 68417 68693 sw
tri 68476 68476 68693 68693 ne
rect 68693 68476 71000 68693
rect 66800 68200 68417 68476
tri 68417 68200 68693 68476 sw
tri 68693 68400 68769 68476 ne
rect 68769 68400 71000 68476
rect 66800 68116 71000 68200
rect 66800 68113 70613 68116
tri 66600 67829 66800 68029 sw
tri 66800 67829 67084 68113 ne
rect 67084 67829 70613 68113
rect 65200 67545 66800 67829
tri 66800 67545 67084 67829 sw
tri 67084 67545 67368 67829 ne
rect 67368 67545 70613 67829
rect 65200 67449 67084 67545
tri 65000 67166 65200 67366 sw
tri 65200 67166 65483 67449 ne
rect 65483 67368 67084 67449
tri 67084 67368 67261 67545 sw
tri 67368 67368 67545 67545 ne
rect 67545 67368 70613 67545
rect 65483 67166 67261 67368
rect 63600 66883 65200 67166
tri 65200 66883 65483 67166 sw
tri 65483 66883 65766 67166 ne
rect 65766 67084 67261 67166
tri 67261 67084 67545 67368 sw
tri 67545 67084 67829 67368 ne
rect 67829 67084 70613 67368
rect 65766 66883 67545 67084
rect 63600 66786 65483 66883
tri 63400 66494 63600 66694 sw
tri 63600 66494 63892 66786 ne
rect 63892 66600 65483 66786
tri 65483 66600 65766 66883 sw
tri 65766 66600 66049 66883 ne
rect 66049 66800 67545 66883
tri 67545 66800 67829 67084 sw
tri 67829 66800 68113 67084 ne
rect 68113 66916 70613 67084
rect 70669 66916 71000 68116
rect 68113 66800 71000 66916
rect 66049 66600 67829 66800
tri 67829 66600 68029 66800 sw
rect 63892 66494 65766 66600
rect 62000 66202 63600 66494
tri 63600 66202 63892 66494 sw
tri 63892 66202 64184 66494 ne
rect 64184 66332 65766 66494
tri 65766 66332 66034 66600 sw
tri 66049 66332 66317 66600 ne
rect 66317 66332 71000 66600
rect 64184 66202 66034 66332
rect 62000 66114 63892 66202
tri 61800 65831 62000 66031 sw
tri 62000 65831 62283 66114 ne
rect 62283 65964 63892 66114
tri 63892 65964 64130 66202 sw
tri 64184 65964 64422 66202 ne
rect 64422 66049 66034 66202
tri 66034 66049 66317 66332 sw
tri 66317 66049 66600 66332 ne
rect 66600 66049 71000 66332
rect 64422 65964 66317 66049
rect 62283 65831 64130 65964
rect 60400 65663 62000 65831
tri 62000 65663 62168 65831 sw
tri 62283 65663 62451 65831 ne
rect 62451 65672 64130 65831
tri 64130 65672 64422 65964 sw
tri 64422 65672 64714 65964 ne
rect 64714 65766 66317 65964
tri 66317 65766 66600 66049 sw
tri 66600 65766 66883 66049 ne
rect 66883 65766 71000 66049
rect 64714 65672 66600 65766
rect 62451 65663 64422 65672
rect 60400 65451 62168 65663
tri 60200 65166 60400 65366 sw
tri 60400 65166 60685 65451 ne
rect 60685 65380 62168 65451
tri 62168 65380 62451 65663 sw
tri 62451 65380 62734 65663 ne
rect 62734 65380 64422 65663
tri 64422 65380 64714 65672 sw
tri 64714 65380 65006 65672 ne
rect 65006 65483 66600 65672
tri 66600 65483 66883 65766 sw
tri 66883 65483 67166 65766 ne
rect 67166 65483 71000 65766
rect 65006 65380 66883 65483
rect 60685 65166 62451 65380
rect 58800 64881 60400 65166
tri 60400 64881 60685 65166 sw
tri 60685 64881 60970 65166 ne
rect 60970 65097 62451 65166
tri 62451 65097 62734 65380 sw
tri 62734 65097 63017 65380 ne
rect 63017 65292 64714 65380
tri 64714 65292 64802 65380 sw
tri 65006 65292 65094 65380 ne
rect 65094 65292 66883 65380
rect 63017 65097 64802 65292
rect 60970 64997 62734 65097
tri 62734 64997 62834 65097 sw
tri 63017 64997 63117 65097 ne
rect 63117 65000 64802 65097
tri 64802 65000 65094 65292 sw
tri 65094 65000 65386 65292 ne
rect 65386 65200 66883 65292
tri 66883 65200 67166 65483 sw
tri 67166 65200 67449 65483 ne
rect 67449 65200 71000 65483
rect 65386 65000 67166 65200
tri 67166 65000 67366 65200 sw
rect 63117 64997 65094 65000
rect 60970 64881 62834 64997
rect 58800 64786 60685 64881
tri 58600 64499 58800 64699 sw
tri 58800 64499 59087 64786 ne
rect 59087 64730 60685 64786
tri 60685 64730 60836 64881 sw
tri 60970 64730 61121 64881 ne
rect 61121 64730 62834 64881
rect 59087 64499 60836 64730
rect 57200 64447 58800 64499
tri 58800 64447 58852 64499 sw
tri 59087 64447 59139 64499 ne
rect 59139 64447 60836 64499
rect 57200 64160 58852 64447
tri 58852 64160 59139 64447 sw
tri 59139 64160 59426 64447 ne
rect 59426 64445 60836 64447
tri 60836 64445 61121 64730 sw
tri 61121 64445 61406 64730 ne
rect 61406 64714 62834 64730
tri 62834 64714 63117 64997 sw
tri 63117 64714 63400 64997 ne
rect 63400 64714 65094 64997
rect 61406 64445 63117 64714
rect 59426 64160 61121 64445
tri 61121 64160 61406 64445 sw
tri 61406 64160 61691 64445 ne
rect 61691 64431 63117 64445
tri 63117 64431 63400 64714 sw
tri 63400 64431 63683 64714 ne
rect 63683 64708 65094 64714
tri 65094 64708 65386 65000 sw
tri 65386 64708 65678 65000 ne
rect 65678 64708 71000 65000
rect 63683 64431 65386 64708
rect 61691 64160 63400 64431
rect 57200 64119 59139 64160
tri 57000 63836 57200 64036 sw
tri 57200 63836 57483 64119 ne
rect 57483 63873 59139 64119
tri 59139 63873 59426 64160 sw
tri 59426 63873 59713 64160 ne
rect 59713 64065 61406 64160
tri 61406 64065 61501 64160 sw
tri 61691 64065 61786 64160 ne
rect 61786 64148 63400 64160
tri 63400 64148 63683 64431 sw
tri 63683 64148 63966 64431 ne
rect 63966 64416 65386 64431
tri 65386 64416 65678 64708 sw
tri 65678 64416 65970 64708 ne
rect 65970 64416 71000 64708
rect 63966 64184 65678 64416
tri 65678 64184 65910 64416 sw
tri 65970 64184 66202 64416 ne
rect 66202 64184 71000 64416
rect 63966 64148 65910 64184
rect 61786 64065 63683 64148
rect 59713 63873 61501 64065
rect 57483 63836 59426 63873
rect 55600 63553 57200 63836
tri 57200 63553 57483 63836 sw
tri 57483 63553 57766 63836 ne
rect 57766 63673 59426 63836
tri 59426 63673 59626 63873 sw
tri 59713 63673 59913 63873 ne
rect 59913 63780 61501 63873
tri 61501 63780 61786 64065 sw
tri 61786 63780 62071 64065 ne
rect 62071 63966 63683 64065
tri 63683 63966 63865 64148 sw
tri 63966 63966 64148 64148 ne
rect 64148 63966 65910 64148
rect 62071 63780 63865 63966
rect 59913 63673 61786 63780
rect 57766 63553 59626 63673
rect 55600 63506 57483 63553
tri 57483 63506 57530 63553 sw
tri 57766 63506 57813 63553 ne
rect 57813 63506 59626 63553
rect 55600 63456 57530 63506
tri 55400 63173 55600 63373 sw
tri 55600 63173 55883 63456 ne
rect 55883 63223 57530 63456
tri 57530 63223 57813 63506 sw
tri 57813 63223 58096 63506 ne
rect 58096 63386 59626 63506
tri 59626 63386 59913 63673 sw
tri 59913 63386 60200 63673 ne
rect 60200 63495 61786 63673
tri 61786 63495 62071 63780 sw
tri 62071 63495 62356 63780 ne
rect 62356 63683 63865 63780
tri 63865 63683 64148 63966 sw
tri 64148 63683 64431 63966 ne
rect 64431 63892 65910 63966
tri 65910 63892 66202 64184 sw
tri 66202 63892 66494 64184 ne
rect 66494 63892 71000 64184
rect 64431 63683 66202 63892
rect 62356 63495 64148 63683
rect 60200 63386 62071 63495
rect 58096 63223 59913 63386
rect 55883 63173 57813 63223
rect 54000 62940 55600 63173
tri 55600 62940 55833 63173 sw
tri 55883 62940 56116 63173 ne
rect 56116 62940 57813 63173
tri 57813 62940 58096 63223 sw
tri 58096 62940 58379 63223 ne
rect 58379 63099 59913 63223
tri 59913 63099 60200 63386 sw
tri 60200 63099 60487 63386 ne
rect 60487 63210 62071 63386
tri 62071 63210 62356 63495 sw
tri 62356 63210 62641 63495 ne
rect 62641 63400 64148 63495
tri 64148 63400 64431 63683 sw
tri 64431 63400 64714 63683 ne
rect 64714 63600 66202 63683
tri 66202 63600 66494 63892 sw
tri 66494 63600 66786 63892 ne
rect 66786 63600 71000 63892
rect 64714 63400 66494 63600
tri 66494 63400 66694 63600 sw
rect 62641 63210 64431 63400
rect 60487 63099 62356 63210
rect 58379 62940 60200 63099
rect 54000 62793 55833 62940
tri 53800 62507 54000 62707 sw
tri 54000 62507 54286 62793 ne
rect 54286 62657 55833 62793
tri 55833 62657 56116 62940 sw
tri 56116 62657 56399 62940 ne
rect 56399 62843 58096 62940
tri 58096 62843 58193 62940 sw
tri 58379 62843 58476 62940 ne
rect 58476 62843 60200 62940
rect 56399 62657 58193 62843
rect 54286 62622 56116 62657
tri 56116 62622 56151 62657 sw
tri 56399 62622 56434 62657 ne
rect 56434 62622 58193 62657
rect 54286 62507 56151 62622
rect 52400 62221 54000 62507
tri 54000 62221 54286 62507 sw
tri 54286 62221 54572 62507 ne
rect 54572 62339 56151 62507
tri 56151 62339 56434 62622 sw
tri 56434 62339 56717 62622 ne
rect 56717 62560 58193 62622
tri 58193 62560 58476 62843 sw
tri 58476 62560 58759 62843 ne
rect 58759 62812 60200 62843
tri 60200 62812 60487 63099 sw
tri 60487 62812 60774 63099 ne
rect 60774 62925 62356 63099
tri 62356 62925 62641 63210 sw
tri 62641 62925 62926 63210 ne
rect 62926 63117 64431 63210
tri 64431 63117 64714 63400 sw
tri 64714 63117 64997 63400 ne
rect 64997 63117 71000 63400
rect 62926 62925 64714 63117
rect 60774 62812 62641 62925
rect 58759 62754 60487 62812
tri 60487 62754 60545 62812 sw
tri 60774 62754 60832 62812 ne
rect 60832 62754 62641 62812
rect 58759 62560 60545 62754
rect 56717 62339 58476 62560
rect 54572 62221 56434 62339
rect 52400 62127 54286 62221
tri 52200 61839 52400 62039 sw
tri 52400 61839 52688 62127 ne
rect 52688 62006 54286 62127
tri 54286 62006 54501 62221 sw
tri 54572 62006 54787 62221 ne
rect 54787 62056 56434 62221
tri 56434 62056 56717 62339 sw
tri 56717 62056 57000 62339 ne
rect 57000 62277 58476 62339
tri 58476 62277 58759 62560 sw
tri 58759 62277 59042 62560 ne
rect 59042 62467 60545 62560
tri 60545 62467 60832 62754 sw
tri 60832 62467 61119 62754 ne
rect 61119 62750 62641 62754
tri 62641 62750 62816 62925 sw
tri 62926 62750 63101 62925 ne
rect 63101 62834 64714 62925
tri 64714 62834 64997 63117 sw
tri 64997 62834 65280 63117 ne
rect 65280 62834 71000 63117
rect 63101 62750 64997 62834
rect 61119 62467 62816 62750
rect 59042 62277 60832 62467
rect 57000 62056 58759 62277
rect 54787 62006 56717 62056
rect 52688 61839 54501 62006
rect 50800 61720 52400 61839
tri 52400 61720 52519 61839 sw
tri 52688 61720 52807 61839 ne
rect 52807 61720 54501 61839
tri 54501 61720 54787 62006 sw
tri 54787 61720 55073 62006 ne
rect 55073 61773 56717 62006
tri 56717 61773 57000 62056 sw
tri 57000 61773 57283 62056 ne
rect 57283 61994 58759 62056
tri 58759 61994 59042 62277 sw
tri 59042 61994 59325 62277 ne
rect 59325 62180 60832 62277
tri 60832 62180 61119 62467 sw
tri 61119 62180 61406 62467 ne
rect 61406 62465 62816 62467
tri 62816 62465 63101 62750 sw
tri 63101 62465 63386 62750 ne
rect 63386 62566 64997 62750
tri 64997 62566 65265 62834 sw
tri 65280 62566 65548 62834 ne
rect 65548 62566 71000 62834
rect 63386 62465 65265 62566
rect 61406 62180 63101 62465
tri 63101 62180 63386 62465 sw
tri 63386 62180 63671 62465 ne
rect 63671 62283 65265 62465
tri 65265 62283 65548 62566 sw
tri 65548 62283 65831 62566 ne
rect 65831 62283 71000 62566
rect 63671 62180 65548 62283
rect 59325 61994 61119 62180
rect 57283 61773 59042 61994
rect 55073 61720 57000 61773
rect 50800 61459 52519 61720
tri 50600 61175 50800 61375 sw
tri 50800 61175 51084 61459 ne
rect 51084 61432 52519 61459
tri 52519 61432 52807 61720 sw
tri 52807 61432 53095 61720 ne
rect 53095 61626 54787 61720
tri 54787 61626 54881 61720 sw
tri 55073 61626 55167 61720 ne
rect 55167 61626 57000 61720
rect 53095 61432 54881 61626
rect 51084 61303 52807 61432
tri 52807 61303 52936 61432 sw
tri 53095 61303 53224 61432 ne
rect 53224 61340 54881 61432
tri 54881 61340 55167 61626 sw
tri 55167 61340 55453 61626 ne
rect 55453 61490 57000 61626
tri 57000 61490 57283 61773 sw
tri 57283 61490 57566 61773 ne
rect 57566 61711 59042 61773
tri 59042 61711 59325 61994 sw
tri 59325 61711 59608 61994 ne
rect 59608 61893 61119 61994
tri 61119 61893 61406 62180 sw
tri 61406 61893 61693 62180 ne
rect 61693 62085 63386 62180
tri 63386 62085 63481 62180 sw
tri 63671 62085 63766 62180 ne
rect 63766 62085 65548 62180
rect 61693 61893 63481 62085
rect 59608 61711 61406 61893
rect 57566 61526 59325 61711
tri 59325 61526 59510 61711 sw
tri 59608 61526 59793 61711 ne
rect 59793 61606 61406 61711
tri 61406 61606 61693 61893 sw
tri 61693 61606 61980 61893 ne
rect 61980 61800 63481 61893
tri 63481 61800 63766 62085 sw
tri 63766 61800 64051 62085 ne
rect 64051 62000 65548 62085
tri 65548 62000 65831 62283 sw
tri 65831 62000 66114 62283 ne
rect 66114 62000 71000 62283
rect 64051 61800 65831 62000
tri 65831 61800 66031 62000 sw
rect 61980 61606 63766 61800
rect 59793 61526 61693 61606
rect 57566 61490 59510 61526
rect 55453 61340 57283 61490
rect 53224 61303 55167 61340
rect 51084 61175 52936 61303
rect 49200 60891 50800 61175
tri 50800 60891 51084 61175 sw
tri 51084 60891 51368 61175 ne
rect 51368 61015 52936 61175
tri 52936 61015 53224 61303 sw
tri 53224 61015 53512 61303 ne
rect 53512 61054 55167 61303
tri 55167 61054 55453 61340 sw
tri 55453 61054 55739 61340 ne
rect 55739 61243 57283 61340
tri 57283 61243 57530 61490 sw
tri 57566 61243 57813 61490 ne
rect 57813 61243 59510 61490
tri 59510 61243 59793 61526 sw
tri 59793 61243 60076 61526 ne
rect 60076 61319 61693 61526
tri 61693 61319 61980 61606 sw
tri 61980 61319 62267 61606 ne
rect 62267 61515 63766 61606
tri 63766 61515 64051 61800 sw
tri 64051 61515 64336 61800 ne
rect 64336 61515 71000 61800
rect 62267 61319 64051 61515
rect 60076 61243 61980 61319
rect 55739 61054 57530 61243
rect 53512 61015 55453 61054
rect 51368 60891 53224 61015
rect 49200 60795 51084 60891
tri 49000 60510 49200 60710 sw
tri 49200 60510 49485 60795 ne
rect 49485 60784 51084 60795
tri 51084 60784 51191 60891 sw
tri 51368 60784 51475 60891 ne
rect 51475 60784 53224 60891
rect 49485 60510 51191 60784
rect 46000 60500 49200 60510
tri 49200 60500 49210 60510 sw
tri 49485 60500 49495 60510 ne
rect 49495 60500 51191 60510
tri 51191 60500 51475 60784 sw
tri 51475 60500 51759 60784 ne
rect 51759 60727 53224 60784
tri 53224 60727 53512 61015 sw
tri 53512 60727 53800 61015 ne
rect 53800 60768 55453 61015
tri 55453 60768 55739 61054 sw
tri 55739 60768 56025 61054 ne
rect 56025 60960 57530 61054
tri 57530 60960 57813 61243 sw
tri 57813 60960 58096 61243 ne
rect 58096 60960 59793 61243
tri 59793 60960 60076 61243 sw
tri 60076 60960 60359 61243 ne
rect 60359 61154 61980 61243
tri 61980 61154 62145 61319 sw
tri 62267 61154 62432 61319 ne
rect 62432 61230 64051 61319
tri 64051 61230 64336 61515 sw
tri 64336 61230 64621 61515 ne
rect 64621 61230 71000 61515
rect 62432 61154 64336 61230
rect 60359 60960 62145 61154
rect 56025 60768 57813 60960
rect 53800 60727 55739 60768
rect 51759 60500 53512 60727
rect 46000 60215 49210 60500
tri 49210 60215 49495 60500 sw
tri 49495 60215 49780 60500 ne
rect 49780 60404 51475 60500
tri 51475 60404 51571 60500 sw
tri 51759 60404 51855 60500 ne
rect 51855 60439 53512 60500
tri 53512 60439 53800 60727 sw
tri 53800 60439 54088 60727 ne
rect 54088 60482 55739 60727
tri 55739 60482 56025 60768 sw
tri 56025 60482 56311 60768 ne
rect 56311 60677 57813 60768
tri 57813 60677 58096 60960 sw
tri 58096 60677 58379 60960 ne
rect 58379 60863 60076 60960
tri 60076 60863 60173 60960 sw
tri 60359 60863 60456 60960 ne
rect 60456 60867 62145 60960
tri 62145 60867 62432 61154 sw
tri 62432 60867 62719 61154 ne
rect 62719 60970 64336 61154
tri 64336 60970 64596 61230 sw
tri 64621 60970 64881 61230 ne
rect 64881 60970 71000 61230
rect 62719 60867 64596 60970
rect 60456 60863 62432 60867
rect 58379 60677 60173 60863
rect 56311 60482 58096 60677
rect 54088 60439 56025 60482
rect 51855 60404 53800 60439
rect 49780 60215 51571 60404
rect 46000 59965 49495 60215
tri 49495 59965 49745 60215 sw
tri 49780 59965 50030 60215 ne
rect 50030 60120 51571 60215
tri 51571 60120 51855 60404 sw
tri 51855 60120 52139 60404 ne
rect 52139 60151 53800 60404
tri 53800 60151 54088 60439 sw
tri 54088 60151 54376 60439 ne
rect 54376 60312 56025 60439
tri 56025 60312 56195 60482 sw
tri 56311 60312 56481 60482 ne
rect 56481 60394 58096 60482
tri 58096 60394 58379 60677 sw
tri 58379 60394 58662 60677 ne
rect 58662 60580 60173 60677
tri 60173 60580 60456 60863 sw
tri 60456 60580 60739 60863 ne
rect 60739 60580 62432 60863
tri 62432 60580 62719 60867 sw
tri 62719 60580 63006 60867 ne
rect 63006 60685 64596 60867
tri 64596 60685 64881 60970 sw
tri 64881 60685 65166 60970 ne
rect 65166 60685 71000 60970
rect 63006 60580 64881 60685
rect 58662 60394 60456 60580
rect 56481 60312 58379 60394
rect 54376 60151 56195 60312
rect 52139 60120 54088 60151
rect 50030 60059 51855 60120
tri 51855 60059 51916 60120 sw
tri 52139 60059 52200 60120 ne
rect 52200 60059 54088 60120
rect 50030 59965 51916 60059
rect 46000 59680 49745 59965
tri 49745 59680 50030 59965 sw
tri 50030 59680 50315 59965 ne
rect 50315 59775 51916 59965
tri 51916 59775 52200 60059 sw
tri 52200 59775 52484 60059 ne
rect 52484 60028 54088 60059
tri 54088 60028 54211 60151 sw
tri 54376 60028 54499 60151 ne
rect 54499 60028 56195 60151
rect 52484 59775 54211 60028
rect 50315 59680 52200 59775
rect 46000 59461 50030 59680
tri 45800 59150 46000 59350 sw
tri 46000 59150 46311 59461 ne
rect 46311 59395 50030 59461
tri 50030 59395 50315 59680 sw
tri 50315 59395 50600 59680 ne
rect 50600 59491 52200 59680
tri 52200 59491 52484 59775 sw
tri 52484 59491 52768 59775 ne
rect 52768 59740 54211 59775
tri 54211 59740 54499 60028 sw
tri 54499 59740 54787 60028 ne
rect 54787 60026 56195 60028
tri 56195 60026 56481 60312 sw
tri 56481 60026 56767 60312 ne
rect 56767 60111 58379 60312
tri 58379 60111 58662 60394 sw
tri 58662 60111 58945 60394 ne
rect 58945 60297 60456 60394
tri 60456 60297 60739 60580 sw
tri 60739 60297 61022 60580 ne
rect 61022 60487 62719 60580
tri 62719 60487 62812 60580 sw
tri 63006 60487 63099 60580 ne
rect 63099 60487 64881 60580
rect 61022 60297 62812 60487
rect 58945 60111 60739 60297
rect 56767 60026 58662 60111
rect 54787 59740 56481 60026
tri 56481 59740 56767 60026 sw
tri 56767 59740 57053 60026 ne
rect 57053 59926 58662 60026
tri 58662 59926 58847 60111 sw
tri 58945 59926 59130 60111 ne
rect 59130 60014 60739 60111
tri 60739 60014 61022 60297 sw
tri 61022 60014 61305 60297 ne
rect 61305 60200 62812 60297
tri 62812 60200 63099 60487 sw
tri 63099 60200 63386 60487 ne
rect 63386 60400 64881 60487
tri 64881 60400 65166 60685 sw
tri 65166 60400 65451 60685 ne
rect 65451 60400 71000 60685
rect 63386 60200 65166 60400
tri 65166 60200 65366 60400 sw
rect 61305 60014 63099 60200
rect 59130 59926 61022 60014
rect 57053 59740 58847 59926
rect 52768 59491 54499 59740
rect 50600 59395 52484 59491
rect 46311 59150 50315 59395
rect 42800 58920 46000 59150
tri 46000 58920 46230 59150 sw
tri 46311 58920 46541 59150 ne
rect 46541 59110 50315 59150
tri 50315 59110 50600 59395 sw
tri 50600 59110 50885 59395 ne
rect 50885 59207 52484 59395
tri 52484 59207 52768 59491 sw
tri 52768 59207 53052 59491 ne
rect 53052 59452 54499 59491
tri 54499 59452 54787 59740 sw
tri 54787 59452 55075 59740 ne
rect 55075 59646 56767 59740
tri 56767 59646 56861 59740 sw
tri 57053 59646 57147 59740 ne
rect 57147 59646 58847 59740
rect 55075 59452 56861 59646
rect 53052 59207 54787 59452
rect 50885 59110 52768 59207
rect 46541 58920 50600 59110
rect 42800 58747 46230 58920
tri 46230 58747 46403 58920 sw
tri 46541 58747 46714 58920 ne
rect 46714 58825 50600 58920
tri 50600 58825 50885 59110 sw
tri 50885 58825 51170 59110 ne
rect 51170 59088 52768 59110
tri 52768 59088 52887 59207 sw
tri 53052 59088 53171 59207 ne
rect 53171 59164 54787 59207
tri 54787 59164 55075 59452 sw
tri 55075 59164 55363 59452 ne
rect 55363 59360 56861 59452
tri 56861 59360 57147 59646 sw
tri 57147 59360 57433 59646 ne
rect 57433 59643 58847 59646
tri 58847 59643 59130 59926 sw
tri 59130 59643 59413 59926 ne
rect 59413 59731 61022 59926
tri 61022 59731 61305 60014 sw
tri 61305 59731 61588 60014 ne
rect 61588 59913 63099 60014
tri 63099 59913 63386 60200 sw
tri 63386 59913 63673 60200 ne
rect 63673 60120 71000 60200
rect 63673 59913 70613 60120
rect 61588 59731 63386 59913
rect 59413 59643 61305 59731
rect 57433 59360 59130 59643
tri 59130 59360 59413 59643 sw
tri 59413 59360 59696 59643 ne
rect 59696 59546 61305 59643
tri 61305 59546 61490 59731 sw
tri 61588 59546 61773 59731 ne
rect 61773 59626 63386 59731
tri 63386 59626 63673 59913 sw
tri 63673 59626 63960 59913 ne
rect 63960 59626 70613 59913
rect 61773 59546 63673 59626
rect 59696 59360 61490 59546
rect 55363 59164 57147 59360
rect 53171 59088 55075 59164
rect 51170 58825 52887 59088
rect 46714 58805 50885 58825
tri 50885 58805 50905 58825 sw
tri 51170 58805 51190 58825 ne
rect 51190 58805 52887 58825
rect 46714 58747 50905 58805
rect 42800 58436 46403 58747
tri 46403 58436 46714 58747 sw
tri 46714 58436 47025 58747 ne
rect 47025 58520 50905 58747
tri 50905 58520 51190 58805 sw
tri 51190 58520 51475 58805 ne
rect 51475 58804 52887 58805
tri 52887 58804 53171 59088 sw
tri 53171 58804 53455 59088 ne
rect 53455 58876 55075 59088
tri 55075 58876 55363 59164 sw
tri 55363 58876 55651 59164 ne
rect 55651 59074 57147 59164
tri 57147 59074 57433 59360 sw
tri 57433 59074 57719 59360 ne
rect 57719 59263 59413 59360
tri 59413 59263 59510 59360 sw
tri 59696 59263 59793 59360 ne
rect 59793 59263 61490 59360
tri 61490 59263 61773 59546 sw
tri 61773 59263 62056 59546 ne
rect 62056 59374 63673 59546
tri 63673 59374 63925 59626 sw
tri 63960 59374 64212 59626 ne
rect 64212 59374 70613 59626
rect 62056 59263 63925 59374
rect 57719 59074 59510 59263
rect 55651 58876 57433 59074
rect 53455 58804 55363 58876
rect 51475 58520 53171 58804
tri 53171 58520 53455 58804 sw
tri 53455 58520 53739 58804 ne
rect 53739 58716 55363 58804
tri 55363 58716 55523 58876 sw
tri 55651 58716 55811 58876 ne
rect 55811 58788 57433 58876
tri 57433 58788 57719 59074 sw
tri 57719 58788 58005 59074 ne
rect 58005 58980 59510 59074
tri 59510 58980 59793 59263 sw
tri 59793 58980 60076 59263 ne
rect 60076 58980 61773 59263
tri 61773 58980 62056 59263 sw
tri 62056 58980 62339 59263 ne
rect 62339 59087 63925 59263
tri 63925 59087 64212 59374 sw
tri 64212 59087 64499 59374 ne
rect 64499 59087 70613 59374
rect 62339 58980 64212 59087
rect 58005 58788 59793 58980
rect 55811 58716 57719 58788
rect 53739 58520 55523 58716
rect 47025 58436 51190 58520
rect 42800 58125 46714 58436
tri 46714 58125 47025 58436 sw
tri 47025 58125 47336 58436 ne
rect 47336 58235 51190 58436
tri 51190 58235 51475 58520 sw
tri 51475 58235 51760 58520 ne
rect 51760 58424 53455 58520
tri 53455 58424 53551 58520 sw
tri 53739 58424 53835 58520 ne
rect 53835 58428 55523 58520
tri 55523 58428 55811 58716 sw
tri 55811 58428 56099 58716 ne
rect 56099 58502 57719 58716
tri 57719 58502 58005 58788 sw
tri 58005 58502 58291 58788 ne
rect 58291 58697 59793 58788
tri 59793 58697 60076 58980 sw
tri 60076 58697 60359 58980 ne
rect 60359 58883 62056 58980
tri 62056 58883 62153 58980 sw
tri 62339 58883 62436 58980 ne
rect 62436 58883 64212 58980
rect 60359 58697 62153 58883
rect 58291 58502 60076 58697
rect 56099 58428 58005 58502
rect 53835 58424 55811 58428
rect 51760 58235 53551 58424
rect 47336 58125 51475 58235
rect 42800 58097 47025 58125
tri 42800 58010 42887 58097 ne
rect 42887 58010 47025 58097
tri 42600 57723 42887 58010 sw
tri 42887 57723 43174 58010 ne
rect 43174 57814 47025 58010
tri 47025 57814 47336 58125 sw
tri 47336 57814 47647 58125 ne
rect 47647 57950 51475 58125
tri 51475 57950 51760 58235 sw
tri 51760 57950 52045 58235 ne
rect 52045 58140 53551 58235
tri 53551 58140 53835 58424 sw
tri 53835 58140 54119 58424 ne
rect 54119 58140 55811 58424
tri 55811 58140 56099 58428 sw
tri 56099 58140 56387 58428 ne
rect 56387 58332 58005 58428
tri 58005 58332 58175 58502 sw
tri 58291 58332 58461 58502 ne
rect 58461 58414 60076 58502
tri 60076 58414 60359 58697 sw
tri 60359 58414 60642 58697 ne
rect 60642 58600 62153 58697
tri 62153 58600 62436 58883 sw
tri 62436 58600 62719 58883 ne
rect 62719 58800 64212 58883
tri 64212 58800 64499 59087 sw
tri 64499 58800 64786 59087 ne
rect 64786 58920 70613 59087
rect 70669 58920 71000 60120
rect 64786 58800 71000 58920
rect 62719 58600 64499 58800
tri 64499 58600 64699 58800 sw
rect 60642 58414 62436 58600
rect 58461 58332 60359 58414
rect 56387 58140 58175 58332
rect 52045 57950 53835 58140
rect 47647 57814 51760 57950
rect 43174 57723 47336 57814
rect 41200 57436 42887 57723
tri 42887 57436 43174 57723 sw
tri 43174 57436 43461 57723 ne
rect 43461 57503 47336 57723
tri 47336 57503 47647 57814 sw
tri 47647 57503 47958 57814 ne
rect 47958 57665 51760 57814
tri 51760 57665 52045 57950 sw
tri 52045 57665 52330 57950 ne
rect 52330 57856 53835 57950
tri 53835 57856 54119 58140 sw
tri 54119 57856 54403 58140 ne
rect 54403 58048 56099 58140
tri 56099 58048 56191 58140 sw
tri 56387 58048 56479 58140 ne
rect 56479 58048 58175 58140
rect 54403 57856 56191 58048
rect 52330 57665 54119 57856
rect 47958 57503 52045 57665
rect 43461 57436 47647 57503
rect 41200 57430 43174 57436
tri 41000 57138 41200 57338 sw
tri 41200 57138 41492 57430 ne
rect 41492 57321 43174 57430
tri 43174 57321 43289 57436 sw
tri 43461 57321 43576 57436 ne
rect 43576 57321 47647 57436
rect 41492 57138 43289 57321
rect 39600 56910 41200 57138
tri 41200 56910 41428 57138 sw
tri 41492 56910 41720 57138 ne
rect 41720 57034 43289 57138
tri 43289 57034 43576 57321 sw
tri 43576 57034 43863 57321 ne
rect 43863 57192 47647 57321
tri 47647 57192 47958 57503 sw
tri 47958 57192 48269 57503 ne
rect 48269 57395 52045 57503
tri 52045 57395 52315 57665 sw
tri 52330 57395 52600 57665 ne
rect 52600 57572 54119 57665
tri 54119 57572 54403 57856 sw
tri 54403 57572 54687 57856 ne
rect 54687 57760 56191 57856
tri 56191 57760 56479 58048 sw
tri 56479 57760 56767 58048 ne
rect 56767 58046 58175 58048
tri 58175 58046 58461 58332 sw
tri 58461 58046 58747 58332 ne
rect 58747 58131 60359 58332
tri 60359 58131 60642 58414 sw
tri 60642 58131 60925 58414 ne
rect 60925 58317 62436 58414
tri 62436 58317 62719 58600 sw
tri 62719 58317 63002 58600 ne
rect 63002 58317 71000 58600
rect 60925 58131 62719 58317
rect 58747 58046 60642 58131
rect 56767 57760 58461 58046
tri 58461 57760 58747 58046 sw
tri 58747 57760 59033 58046 ne
rect 59033 57946 60642 58046
tri 60642 57946 60827 58131 sw
tri 60925 57946 61110 58131 ne
rect 61110 58034 62719 58131
tri 62719 58034 63002 58317 sw
tri 63002 58034 63285 58317 ne
rect 63285 58034 71000 58317
rect 61110 57946 63002 58034
rect 59033 57760 60827 57946
rect 54687 57572 56479 57760
rect 52600 57395 54403 57572
rect 48269 57192 52315 57395
rect 43863 57034 47958 57192
rect 41720 56910 43576 57034
rect 39600 56758 41428 56910
tri 39400 56465 39600 56665 sw
tri 39600 56465 39893 56758 ne
rect 39893 56752 41428 56758
tri 41428 56752 41586 56910 sw
tri 41720 56752 41878 56910 ne
rect 41878 56752 43576 56910
rect 39893 56465 41586 56752
rect 36400 56172 39600 56465
tri 39600 56172 39893 56465 sw
tri 39893 56172 40186 56465 ne
rect 40186 56460 41586 56465
tri 41586 56460 41878 56752 sw
tri 41878 56460 42170 56752 ne
rect 42170 56747 43576 56752
tri 43576 56747 43863 57034 sw
tri 43863 56747 44150 57034 ne
rect 44150 56910 47958 57034
tri 47958 56910 48240 57192 sw
tri 48269 56910 48551 57192 ne
rect 48551 57110 52315 57192
tri 52315 57110 52600 57395 sw
tri 52600 57110 52885 57395 ne
rect 52885 57288 54403 57395
tri 54403 57288 54687 57572 sw
tri 54687 57288 54971 57572 ne
rect 54971 57472 56479 57572
tri 56479 57472 56767 57760 sw
tri 56767 57472 57055 57760 ne
rect 57055 57666 58747 57760
tri 58747 57666 58841 57760 sw
tri 59033 57666 59127 57760 ne
rect 59127 57666 60827 57760
rect 57055 57472 58841 57666
rect 54971 57288 56767 57472
rect 52885 57110 54687 57288
rect 48551 56910 52600 57110
rect 44150 56803 48240 56910
tri 48240 56803 48347 56910 sw
tri 48551 56803 48658 56910 ne
rect 48658 56825 52600 56910
tri 52600 56825 52885 57110 sw
tri 52885 56825 53170 57110 ne
rect 53170 57108 54687 57110
tri 54687 57108 54867 57288 sw
tri 54971 57108 55151 57288 ne
rect 55151 57184 56767 57288
tri 56767 57184 57055 57472 sw
tri 57055 57184 57343 57472 ne
rect 57343 57380 58841 57472
tri 58841 57380 59127 57666 sw
tri 59127 57380 59413 57666 ne
rect 59413 57663 60827 57666
tri 60827 57663 61110 57946 sw
tri 61110 57663 61393 57946 ne
rect 61393 57766 63002 57946
tri 63002 57766 63270 58034 sw
tri 63285 57766 63553 58034 ne
rect 63553 57766 71000 58034
rect 61393 57663 63270 57766
rect 59413 57380 61110 57663
tri 61110 57380 61393 57663 sw
tri 61393 57380 61676 57663 ne
rect 61676 57483 63270 57663
tri 63270 57483 63553 57766 sw
tri 63553 57483 63836 57766 ne
rect 63836 57483 71000 57766
rect 61676 57380 63553 57483
rect 57343 57184 59127 57380
rect 55151 57108 57055 57184
rect 53170 56825 54867 57108
rect 48658 56803 52885 56825
rect 44150 56747 48347 56803
rect 42170 56460 43863 56747
tri 43863 56460 44150 56747 sw
tri 44150 56460 44437 56747 ne
rect 44437 56492 48347 56747
tri 48347 56492 48658 56803 sw
tri 48658 56492 48969 56803 ne
rect 48969 56540 52885 56803
tri 52885 56540 53170 56825 sw
tri 53170 56540 53455 56825 ne
rect 53455 56824 54867 56825
tri 54867 56824 55151 57108 sw
tri 55151 56824 55435 57108 ne
rect 55435 56896 57055 57108
tri 57055 56896 57343 57184 sw
tri 57343 56896 57631 57184 ne
rect 57631 57094 59127 57184
tri 59127 57094 59413 57380 sw
tri 59413 57094 59699 57380 ne
rect 59699 57283 61393 57380
tri 61393 57283 61490 57380 sw
tri 61676 57283 61773 57380 ne
rect 61773 57283 63553 57380
rect 59699 57094 61490 57283
rect 57631 56896 59413 57094
rect 55435 56824 57343 56896
rect 53455 56540 55151 56824
tri 55151 56540 55435 56824 sw
tri 55435 56540 55719 56824 ne
rect 55719 56736 57343 56824
tri 57343 56736 57503 56896 sw
tri 57631 56736 57791 56896 ne
rect 57791 56808 59413 56896
tri 59413 56808 59699 57094 sw
tri 59699 56808 59985 57094 ne
rect 59985 57000 61490 57094
tri 61490 57000 61773 57283 sw
tri 61773 57000 62056 57283 ne
rect 62056 57200 63553 57283
tri 63553 57200 63836 57483 sw
tri 63836 57200 64119 57483 ne
rect 64119 57200 71000 57483
rect 62056 57000 63836 57200
tri 63836 57000 64036 57200 sw
rect 59985 56808 61773 57000
rect 57791 56736 59699 56808
rect 55719 56540 57503 56736
rect 48969 56492 53170 56540
rect 44437 56460 48658 56492
rect 40186 56322 41878 56460
tri 41878 56322 42016 56460 sw
tri 42170 56322 42308 56460 ne
rect 42308 56322 44150 56460
rect 40186 56172 42016 56322
rect 36400 56145 39893 56172
tri 39893 56145 39920 56172 sw
tri 40186 56145 40213 56172 ne
rect 40213 56145 42016 56172
rect 36400 55852 39920 56145
tri 39920 55852 40213 56145 sw
tri 40213 55852 40506 56145 ne
rect 40506 56030 42016 56145
tri 42016 56030 42308 56322 sw
tri 42308 56030 42600 56322 ne
rect 42600 56173 44150 56322
tri 44150 56173 44437 56460 sw
tri 44437 56173 44724 56460 ne
rect 44724 56181 48658 56460
tri 48658 56181 48969 56492 sw
tri 48969 56181 49280 56492 ne
rect 49280 56255 53170 56492
tri 53170 56255 53455 56540 sw
tri 53455 56255 53740 56540 ne
rect 53740 56444 55435 56540
tri 55435 56444 55531 56540 sw
tri 55719 56444 55815 56540 ne
rect 55815 56448 57503 56540
tri 57503 56448 57791 56736 sw
tri 57791 56448 58079 56736 ne
rect 58079 56522 59699 56736
tri 59699 56522 59985 56808 sw
tri 59985 56522 60271 56808 ne
rect 60271 56717 61773 56808
tri 61773 56717 62056 57000 sw
tri 62056 56717 62339 57000 ne
rect 62339 56910 71000 57000
rect 62339 56717 70613 56910
rect 60271 56522 62056 56717
rect 58079 56448 59985 56522
rect 55815 56444 57791 56448
rect 53740 56255 55531 56444
rect 49280 56181 53455 56255
rect 44724 56173 48969 56181
rect 42600 56030 44437 56173
rect 40506 55852 42308 56030
rect 36400 55559 40213 55852
tri 40213 55559 40506 55852 sw
tri 40506 55559 40799 55852 ne
rect 40799 55738 42308 55852
tri 42308 55738 42600 56030 sw
tri 42600 55738 42892 56030 ne
rect 42892 55886 44437 56030
tri 44437 55886 44724 56173 sw
tri 44724 55886 45011 56173 ne
rect 45011 55886 48969 56173
rect 42892 55738 44724 55886
rect 40799 55559 42600 55738
rect 36400 55421 40506 55559
tri 36200 55124 36400 55324 sw
tri 36400 55124 36697 55421 ne
rect 36697 55266 40506 55421
tri 40506 55266 40799 55559 sw
tri 40799 55266 41092 55559 ne
rect 41092 55446 42600 55559
tri 42600 55446 42892 55738 sw
tri 42892 55446 43184 55738 ne
rect 43184 55710 44724 55738
tri 44724 55710 44900 55886 sw
tri 45011 55710 45187 55886 ne
rect 45187 55870 48969 55886
tri 48969 55870 49280 56181 sw
tri 49280 55870 49591 56181 ne
rect 49591 55970 53455 56181
tri 53455 55970 53740 56255 sw
tri 53740 55970 54025 56255 ne
rect 54025 56160 55531 56255
tri 55531 56160 55815 56444 sw
tri 55815 56160 56099 56444 ne
rect 56099 56160 57791 56444
tri 57791 56160 58079 56448 sw
tri 58079 56160 58367 56448 ne
rect 58367 56352 59985 56448
tri 59985 56352 60155 56522 sw
tri 60271 56352 60441 56522 ne
rect 60441 56434 62056 56522
tri 62056 56434 62339 56717 sw
tri 62339 56434 62622 56717 ne
rect 62622 56434 70613 56717
rect 60441 56352 62339 56434
rect 58367 56160 60155 56352
rect 54025 55970 55815 56160
rect 49591 55870 53740 55970
rect 45187 55710 49280 55870
rect 43184 55559 44900 55710
tri 44900 55559 45051 55710 sw
tri 45187 55559 45338 55710 ne
rect 45338 55559 49280 55710
tri 49280 55559 49591 55870 sw
tri 49591 55559 49902 55870 ne
rect 49902 55685 53740 55870
tri 53740 55685 54025 55970 sw
tri 54025 55685 54310 55970 ne
rect 54310 55876 55815 55970
tri 55815 55876 56099 56160 sw
tri 56099 55876 56383 56160 ne
rect 56383 56068 58079 56160
tri 58079 56068 58171 56160 sw
tri 58367 56068 58459 56160 ne
rect 58459 56068 60155 56160
rect 56383 55876 58171 56068
rect 54310 55685 56099 55876
rect 49902 55559 54025 55685
rect 43184 55446 45051 55559
rect 41092 55266 42892 55446
rect 36697 55153 40799 55266
tri 40799 55153 40912 55266 sw
tri 41092 55153 41205 55266 ne
rect 41205 55154 42892 55266
tri 42892 55154 43184 55446 sw
tri 43184 55154 43476 55446 ne
rect 43476 55272 45051 55446
tri 45051 55272 45338 55559 sw
tri 45338 55272 45625 55559 ne
rect 45625 55272 49591 55559
rect 43476 55154 45338 55272
rect 41205 55153 43184 55154
rect 36697 55124 40912 55153
rect 33200 54827 36400 55124
tri 36400 54827 36697 55124 sw
tri 36697 54827 36994 55124 ne
rect 36994 54860 40912 55124
tri 40912 54860 41205 55153 sw
tri 41205 54860 41498 55153 ne
rect 41498 55064 43184 55153
tri 43184 55064 43274 55154 sw
tri 43476 55064 43566 55154 ne
rect 43566 55064 45338 55154
rect 41498 54860 43274 55064
rect 36994 54827 41205 54860
rect 33200 54674 36697 54827
tri 36697 54674 36850 54827 sw
tri 36994 54674 37147 54827 ne
rect 37147 54674 41205 54827
rect 33200 54377 36850 54674
tri 36850 54377 37147 54674 sw
tri 37147 54377 37444 54674 ne
rect 37444 54567 41205 54674
tri 41205 54567 41498 54860 sw
tri 41498 54567 41791 54860 ne
rect 41791 54772 43274 54860
tri 43274 54772 43566 55064 sw
tri 43566 54772 43858 55064 ne
rect 43858 55054 45338 55064
tri 45338 55054 45556 55272 sw
tri 45625 55054 45843 55272 ne
rect 45843 55248 49591 55272
tri 49591 55248 49902 55559 sw
tri 49902 55248 50213 55559 ne
rect 50213 55415 54025 55559
tri 54025 55415 54295 55685 sw
tri 54310 55415 54580 55685 ne
rect 54580 55592 56099 55685
tri 56099 55592 56383 55876 sw
tri 56383 55592 56667 55876 ne
rect 56667 55780 58171 55876
tri 58171 55780 58459 56068 sw
tri 58459 55780 58747 56068 ne
rect 58747 56066 60155 56068
tri 60155 56066 60441 56352 sw
tri 60441 56066 60727 56352 ne
rect 60727 56166 62339 56352
tri 62339 56166 62607 56434 sw
tri 62622 56166 62890 56434 ne
rect 62890 56166 70613 56434
rect 60727 56066 62607 56166
rect 58747 55780 60441 56066
tri 60441 55780 60727 56066 sw
tri 60727 55780 61013 56066 ne
rect 61013 55883 62607 56066
tri 62607 55883 62890 56166 sw
tri 62890 55883 63173 56166 ne
rect 63173 55883 70613 56166
rect 61013 55780 62890 55883
rect 56667 55592 58459 55780
rect 54580 55415 56383 55592
rect 50213 55248 54295 55415
rect 45843 55120 49902 55248
tri 49902 55120 50030 55248 sw
tri 50213 55120 50341 55248 ne
rect 50341 55130 54295 55248
tri 54295 55130 54580 55415 sw
tri 54580 55130 54865 55415 ne
rect 54865 55308 56383 55415
tri 56383 55308 56667 55592 sw
tri 56667 55308 56951 55592 ne
rect 56951 55492 58459 55592
tri 58459 55492 58747 55780 sw
tri 58747 55492 59035 55780 ne
rect 59035 55686 60727 55780
tri 60727 55686 60821 55780 sw
tri 61013 55686 61107 55780 ne
rect 61107 55686 62890 55780
rect 59035 55492 60821 55686
rect 56951 55308 58747 55492
rect 54865 55130 56667 55308
rect 50341 55120 54580 55130
rect 45843 55054 50030 55120
rect 43858 54772 45556 55054
rect 41791 54567 43566 54772
rect 37444 54377 41498 54567
rect 33200 54080 37147 54377
tri 37147 54080 37444 54377 sw
tri 37444 54080 37741 54377 ne
rect 37741 54274 41498 54377
tri 41498 54274 41791 54567 sw
tri 41791 54274 42084 54567 ne
rect 42084 54480 43566 54567
tri 43566 54480 43858 54772 sw
tri 43858 54480 44150 54772 ne
rect 44150 54767 45556 54772
tri 45556 54767 45843 55054 sw
tri 45843 54767 46130 55054 ne
rect 46130 54809 50030 55054
tri 50030 54809 50341 55120 sw
tri 50341 54809 50652 55120 ne
rect 50652 54845 54580 55120
tri 54580 54845 54865 55130 sw
tri 54865 54845 55150 55130 ne
rect 55150 55128 56667 55130
tri 56667 55128 56847 55308 sw
tri 56951 55128 57131 55308 ne
rect 57131 55204 58747 55308
tri 58747 55204 59035 55492 sw
tri 59035 55204 59323 55492 ne
rect 59323 55400 60821 55492
tri 60821 55400 61107 55686 sw
tri 61107 55400 61393 55686 ne
rect 61393 55600 62890 55686
tri 62890 55600 63173 55883 sw
tri 63173 55600 63456 55883 ne
rect 63456 55710 70613 55883
rect 70669 55710 71000 56910
rect 63456 55600 71000 55710
rect 61393 55400 63173 55600
tri 63173 55400 63373 55600 sw
rect 59323 55204 61107 55400
rect 57131 55128 59035 55204
rect 55150 54845 56847 55128
rect 50652 54809 54865 54845
rect 46130 54767 50341 54809
rect 44150 54480 45843 54767
tri 45843 54480 46130 54767 sw
tri 46130 54480 46417 54767 ne
rect 46417 54498 50341 54767
tri 50341 54498 50652 54809 sw
tri 50652 54498 50963 54809 ne
rect 50963 54560 54865 54809
tri 54865 54560 55150 54845 sw
tri 55150 54560 55435 54845 ne
rect 55435 54844 56847 54845
tri 56847 54844 57131 55128 sw
tri 57131 54844 57415 55128 ne
rect 57415 54916 59035 55128
tri 59035 54916 59323 55204 sw
tri 59323 54916 59611 55204 ne
rect 59611 55114 61107 55204
tri 61107 55114 61393 55400 sw
tri 61393 55114 61679 55400 ne
rect 61679 55302 71000 55400
rect 61679 55114 70613 55302
rect 59611 54916 61393 55114
rect 57415 54844 59323 54916
rect 55435 54560 57131 54844
tri 57131 54560 57415 54844 sw
tri 57415 54560 57699 54844 ne
rect 57699 54756 59323 54844
tri 59323 54756 59483 54916 sw
tri 59611 54756 59771 54916 ne
rect 59771 54828 61393 54916
tri 61393 54828 61679 55114 sw
tri 61679 54828 61965 55114 ne
rect 61965 54828 70613 55114
rect 59771 54756 61679 54828
rect 57699 54560 59483 54756
rect 50963 54498 55150 54560
rect 46417 54480 50652 54498
rect 42084 54274 43858 54480
rect 37741 54080 41791 54274
tri 33000 53792 33200 53992 sw
tri 33200 53792 33488 54080 ne
rect 33488 53792 37444 54080
rect 30000 53504 33200 53792
tri 33200 53504 33488 53792 sw
tri 33488 53504 33776 53792 ne
rect 33776 53783 37444 53792
tri 37444 53783 37741 54080 sw
tri 37741 53783 38038 54080 ne
rect 38038 53981 41791 54080
tri 41791 53981 42084 54274 sw
tri 42084 53981 42377 54274 ne
rect 42377 54188 43858 54274
tri 43858 54188 44150 54480 sw
tri 44150 54188 44442 54480 ne
rect 44442 54193 46130 54480
tri 46130 54193 46417 54480 sw
tri 46417 54193 46704 54480 ne
rect 46704 54193 50652 54480
rect 44442 54188 46417 54193
rect 42377 53981 44150 54188
rect 38038 53783 42084 53981
rect 33776 53673 37741 53783
tri 37741 53673 37851 53783 sw
tri 38038 53673 38148 53783 ne
rect 38148 53722 42084 53783
tri 42084 53722 42343 53981 sw
tri 42377 53722 42636 53981 ne
rect 42636 53896 44150 53981
tri 44150 53896 44442 54188 sw
tri 44442 53896 44734 54188 ne
rect 44734 53906 46417 54188
tri 46417 53906 46704 54193 sw
tri 46704 53906 46991 54193 ne
rect 46991 54187 50652 54193
tri 50652 54187 50963 54498 sw
tri 50963 54187 51274 54498 ne
rect 51274 54275 55150 54498
tri 55150 54275 55435 54560 sw
tri 55435 54275 55720 54560 ne
rect 55720 54464 57415 54560
tri 57415 54464 57511 54560 sw
tri 57699 54464 57795 54560 ne
rect 57795 54468 59483 54560
tri 59483 54468 59771 54756 sw
tri 59771 54468 60059 54756 ne
rect 60059 54572 61679 54756
tri 61679 54572 61935 54828 sw
tri 61965 54572 62221 54828 ne
rect 62221 54572 70613 54828
rect 60059 54468 61935 54572
rect 57795 54464 59771 54468
rect 55720 54275 57511 54464
rect 51274 54187 55435 54275
rect 46991 53906 50963 54187
rect 44734 53896 46704 53906
rect 42636 53722 44442 53896
rect 38148 53673 42343 53722
rect 33776 53504 37851 53673
rect 30000 53216 33488 53504
tri 33488 53216 33776 53504 sw
tri 33776 53216 34064 53504 ne
rect 34064 53376 37851 53504
tri 37851 53376 38148 53673 sw
tri 38148 53376 38445 53673 ne
rect 38445 53466 42343 53673
tri 42343 53466 42599 53722 sw
tri 42636 53466 42892 53722 ne
rect 42892 53604 44442 53722
tri 44442 53604 44734 53896 sw
tri 44734 53604 45026 53896 ne
rect 45026 53619 46704 53896
tri 46704 53619 46991 53906 sw
tri 46991 53619 47278 53906 ne
rect 47278 53876 50963 53906
tri 50963 53876 51274 54187 sw
tri 51274 53876 51585 54187 ne
rect 51585 53990 55435 54187
tri 55435 53990 55720 54275 sw
tri 55720 53990 56005 54275 ne
rect 56005 54180 57511 54275
tri 57511 54180 57795 54464 sw
tri 57795 54180 58079 54464 ne
rect 58079 54180 59771 54464
tri 59771 54180 60059 54468 sw
tri 60059 54180 60347 54468 ne
rect 60347 54286 61935 54468
tri 61935 54286 62221 54572 sw
tri 62221 54286 62507 54572 ne
rect 62507 54286 70613 54572
rect 60347 54180 62221 54286
rect 56005 53990 57795 54180
rect 51585 53876 55720 53990
rect 47278 53619 51274 53876
rect 45026 53604 46991 53619
rect 42892 53466 44734 53604
rect 38445 53376 42599 53466
rect 34064 53216 38148 53376
rect 30000 52928 33776 53216
tri 33776 52928 34064 53216 sw
tri 34064 52928 34352 53216 ne
rect 34352 53079 38148 53216
tri 38148 53079 38445 53376 sw
tri 38445 53079 38742 53376 ne
rect 38742 53173 42599 53376
tri 42599 53173 42892 53466 sw
tri 42892 53173 43185 53466 ne
rect 43185 53464 44734 53466
tri 44734 53464 44874 53604 sw
tri 45026 53464 45166 53604 ne
rect 45166 53464 46991 53604
rect 43185 53173 44874 53464
rect 38742 53079 42892 53173
rect 34352 52928 38445 53079
rect 30000 52748 34064 52928
tri 29800 52454 30000 52654 sw
tri 30000 52454 30294 52748 ne
rect 30294 52640 34064 52748
tri 34064 52640 34352 52928 sw
tri 34352 52640 34640 52928 ne
rect 34640 52782 38445 52928
tri 38445 52782 38742 53079 sw
tri 38742 52782 39039 53079 ne
rect 39039 52880 42892 53079
tri 42892 52880 43185 53173 sw
tri 43185 52880 43478 53173 ne
rect 43478 53172 44874 53173
tri 44874 53172 45166 53464 sw
tri 45166 53172 45458 53464 ne
rect 45458 53361 46991 53464
tri 46991 53361 47249 53619 sw
tri 47278 53361 47536 53619 ne
rect 47536 53565 51274 53619
tri 51274 53565 51585 53876 sw
tri 51585 53565 51896 53876 ne
rect 51896 53705 55720 53876
tri 55720 53705 56005 53990 sw
tri 56005 53705 56290 53990 ne
rect 56290 53896 57795 53990
tri 57795 53896 58079 54180 sw
tri 58079 53896 58363 54180 ne
rect 58363 54088 60059 54180
tri 60059 54088 60151 54180 sw
tri 60347 54088 60439 54180 ne
rect 60439 54088 62221 54180
rect 58363 53896 60151 54088
rect 56290 53705 58079 53896
rect 51896 53565 56005 53705
rect 47536 53361 51585 53565
rect 45458 53172 47249 53361
rect 43478 52880 45166 53172
tri 45166 52880 45458 53172 sw
tri 45458 52880 45750 53172 ne
rect 45750 53074 47249 53172
tri 47249 53074 47536 53361 sw
tri 47536 53074 47823 53361 ne
rect 47823 53254 51585 53361
tri 51585 53254 51896 53565 sw
tri 51896 53254 52207 53565 ne
rect 52207 53435 56005 53565
tri 56005 53435 56275 53705 sw
tri 56290 53435 56560 53705 ne
rect 56560 53612 58079 53705
tri 58079 53612 58363 53896 sw
tri 58363 53612 58647 53896 ne
rect 58647 53800 60151 53896
tri 60151 53800 60439 54088 sw
tri 60439 53800 60727 54088 ne
rect 60727 54000 62221 54088
tri 62221 54000 62507 54286 sw
tri 62507 54000 62793 54286 ne
rect 62793 54102 70613 54286
rect 70669 54102 71000 55302
rect 62793 54000 71000 54102
rect 60727 53800 62507 54000
tri 62507 53800 62707 54000 sw
rect 58647 53612 60439 53800
rect 56560 53435 58363 53612
rect 52207 53254 56275 53435
rect 47823 53074 51896 53254
rect 45750 52880 47536 53074
rect 39039 52782 43185 52880
rect 34640 52640 38742 52782
rect 30294 52454 34352 52640
rect 26800 52160 30000 52454
tri 30000 52160 30294 52454 sw
tri 30294 52160 30588 52454 ne
rect 30588 52372 34352 52454
tri 34352 52372 34620 52640 sw
tri 34640 52372 34908 52640 ne
rect 34908 52485 38742 52640
tri 38742 52485 39039 52782 sw
tri 39039 52485 39336 52782 ne
rect 39336 52587 43185 52782
tri 43185 52587 43478 52880 sw
tri 43478 52587 43771 52880 ne
rect 43771 52804 45458 52880
tri 45458 52804 45534 52880 sw
tri 45750 52804 45826 52880 ne
rect 45826 52804 47536 52880
rect 43771 52587 45534 52804
rect 39336 52485 43478 52587
rect 34908 52372 39039 52485
rect 30588 52160 34620 52372
rect 26800 51998 30294 52160
tri 30294 51998 30456 52160 sw
tri 30588 51998 30750 52160 ne
rect 30750 52084 34620 52160
tri 34620 52084 34908 52372 sw
tri 34908 52084 35196 52372 ne
rect 35196 52188 39039 52372
tri 39039 52188 39336 52485 sw
tri 39336 52188 39633 52485 ne
rect 39633 52294 43478 52485
tri 43478 52294 43771 52587 sw
tri 43771 52294 44064 52587 ne
rect 44064 52512 45534 52587
tri 45534 52512 45826 52804 sw
tri 45826 52512 46118 52804 ne
rect 46118 52787 47536 52804
tri 47536 52787 47823 53074 sw
tri 47823 52787 48110 53074 ne
rect 48110 52943 51896 53074
tri 51896 52943 52207 53254 sw
tri 52207 52943 52518 53254 ne
rect 52518 53150 56275 53254
tri 56275 53150 56560 53435 sw
tri 56560 53150 56845 53435 ne
rect 56845 53328 58363 53435
tri 58363 53328 58647 53612 sw
tri 58647 53328 58931 53612 ne
rect 58931 53512 60439 53612
tri 60439 53512 60727 53800 sw
tri 60727 53512 61015 53800 ne
rect 61015 53722 71000 53800
rect 61015 53512 70613 53722
rect 58931 53328 60727 53512
rect 56845 53150 58647 53328
rect 52518 52943 56560 53150
rect 48110 52861 52207 52943
tri 52207 52861 52289 52943 sw
tri 52518 52861 52600 52943 ne
rect 52600 52865 56560 52943
tri 56560 52865 56845 53150 sw
tri 56845 52865 57130 53150 ne
rect 57130 53148 58647 53150
tri 58647 53148 58827 53328 sw
tri 58931 53148 59111 53328 ne
rect 59111 53224 60727 53328
tri 60727 53224 61015 53512 sw
tri 61015 53224 61303 53512 ne
rect 61303 53224 70613 53512
rect 59111 53148 61015 53224
rect 57130 52865 58827 53148
rect 52600 52861 56845 52865
rect 48110 52787 52289 52861
rect 46118 52512 47823 52787
rect 44064 52500 45826 52512
tri 45826 52500 45838 52512 sw
tri 46118 52500 46130 52512 ne
rect 46130 52500 47823 52512
tri 47823 52500 48110 52787 sw
tri 48110 52500 48397 52787 ne
rect 48397 52550 52289 52787
tri 52289 52550 52600 52861 sw
tri 52600 52550 52911 52861 ne
rect 52911 52580 56845 52861
tri 56845 52580 57130 52865 sw
tri 57130 52580 57415 52865 ne
rect 57415 52864 58827 52865
tri 58827 52864 59111 53148 sw
tri 59111 52864 59395 53148 ne
rect 59395 52976 61015 53148
tri 61015 52976 61263 53224 sw
tri 61303 52976 61551 53224 ne
rect 61551 52976 70613 53224
rect 59395 52864 61263 52976
rect 57415 52580 59111 52864
tri 59111 52580 59395 52864 sw
tri 59395 52580 59679 52864 ne
rect 59679 52688 61263 52864
tri 61263 52688 61551 52976 sw
tri 61551 52688 61839 52976 ne
rect 61839 52688 70613 52976
rect 59679 52580 61551 52688
rect 52911 52550 57130 52580
rect 48397 52500 52600 52550
rect 44064 52294 45838 52500
rect 39633 52188 43771 52294
rect 35196 52084 39336 52188
rect 30750 51998 34908 52084
rect 26800 51704 30456 51998
tri 30456 51704 30750 51998 sw
tri 30750 51704 31044 51998 ne
rect 31044 51796 34908 51998
tri 34908 51796 35196 52084 sw
tri 35196 51796 35484 52084 ne
rect 35484 51891 39336 52084
tri 39336 51891 39633 52188 sw
tri 39633 51891 39930 52188 ne
rect 39930 52001 43771 52188
tri 43771 52001 44064 52294 sw
tri 44064 52001 44357 52294 ne
rect 44357 52208 45838 52294
tri 45838 52208 46130 52500 sw
tri 46130 52208 46422 52500 ne
rect 46422 52213 48110 52500
tri 48110 52213 48397 52500 sw
tri 48397 52213 48684 52500 ne
rect 48684 52239 52600 52500
tri 52600 52239 52911 52550 sw
tri 52911 52239 53222 52550 ne
rect 53222 52295 57130 52550
tri 57130 52295 57415 52580 sw
tri 57415 52295 57700 52580 ne
rect 57700 52484 59395 52580
tri 59395 52484 59491 52580 sw
tri 59679 52484 59775 52580 ne
rect 59775 52484 61551 52580
rect 57700 52295 59491 52484
rect 53222 52239 57415 52295
rect 48684 52213 52911 52239
rect 46422 52208 48397 52213
rect 44357 52001 46130 52208
rect 39930 51891 44064 52001
rect 35484 51796 39633 51891
rect 31044 51704 35196 51796
rect 26800 51410 30750 51704
tri 30750 51410 31044 51704 sw
tri 31044 51410 31338 51704 ne
rect 31338 51508 35196 51704
tri 35196 51508 35484 51796 sw
tri 35484 51508 35772 51796 ne
rect 35772 51661 39633 51796
tri 39633 51661 39863 51891 sw
tri 39930 51661 40160 51891 ne
rect 40160 51779 44064 51891
tri 44064 51779 44286 52001 sw
tri 44357 51779 44579 52001 ne
rect 44579 51916 46130 52001
tri 46130 51916 46422 52208 sw
tri 46422 51916 46714 52208 ne
rect 46714 51926 48397 52208
tri 48397 51926 48684 52213 sw
tri 48684 51926 48971 52213 ne
rect 48971 51928 52911 52213
tri 52911 51928 53222 52239 sw
tri 53222 51928 53533 52239 ne
rect 53533 52010 57415 52239
tri 57415 52010 57700 52295 sw
tri 57700 52010 57985 52295 ne
rect 57985 52200 59491 52295
tri 59491 52200 59775 52484 sw
tri 59775 52200 60059 52484 ne
rect 60059 52400 61551 52484
tri 61551 52400 61839 52688 sw
tri 61839 52400 62127 52688 ne
rect 62127 52522 70613 52688
rect 70669 52522 71000 53722
rect 62127 52400 71000 52522
rect 60059 52200 61839 52400
tri 61839 52200 62039 52400 sw
rect 57985 52010 59775 52200
rect 53533 51928 57700 52010
rect 48971 51926 53222 51928
rect 46714 51916 48684 51926
rect 44579 51779 46422 51916
rect 40160 51661 44286 51779
rect 35772 51508 39863 51661
rect 31338 51410 35484 51508
tri 26600 51220 26700 51320 sw
tri 26800 51220 26990 51410 ne
rect 26990 51220 31044 51410
tri 31044 51220 31234 51410 sw
tri 31338 51220 31528 51410 ne
rect 31528 51220 35484 51410
tri 35484 51220 35772 51508 sw
tri 35772 51220 36060 51508 ne
rect 36060 51364 39863 51508
tri 39863 51364 40160 51661 sw
tri 40160 51364 40457 51661 ne
rect 40457 51486 44286 51661
tri 44286 51486 44579 51779 sw
tri 44579 51486 44872 51779 ne
rect 44872 51624 46422 51779
tri 46422 51624 46714 51916 sw
tri 46714 51624 47006 51916 ne
rect 47006 51880 48684 51916
tri 48684 51880 48730 51926 sw
tri 48971 51880 49017 51926 ne
rect 49017 51880 53222 51926
rect 47006 51624 48730 51880
rect 44872 51486 46714 51624
rect 40457 51364 44579 51486
rect 36060 51220 40160 51364
rect 25200 50930 26700 51220
tri 26700 50930 26990 51220 sw
tri 26990 50930 27280 51220 ne
rect 27280 50930 31234 51220
rect 25200 50740 26990 50930
tri 25000 50451 25200 50651 sw
tri 25200 50451 25489 50740 ne
rect 25489 50650 26990 50740
tri 26990 50650 27270 50930 sw
tri 27280 50650 27560 50930 ne
rect 27560 50926 31234 50930
tri 31234 50926 31528 51220 sw
tri 31528 50926 31822 51220 ne
rect 31822 50932 35772 51220
tri 35772 50932 36060 51220 sw
tri 36060 50932 36348 51220 ne
rect 36348 51067 40160 51220
tri 40160 51067 40457 51364 sw
tri 40457 51067 40754 51364 ne
rect 40754 51193 44579 51364
tri 44579 51193 44872 51486 sw
tri 44872 51193 45165 51486 ne
rect 45165 51484 46714 51486
tri 46714 51484 46854 51624 sw
tri 47006 51484 47146 51624 ne
rect 47146 51593 48730 51624
tri 48730 51593 49017 51880 sw
tri 49017 51593 49304 51880 ne
rect 49304 51617 53222 51880
tri 53222 51617 53533 51928 sw
tri 53533 51617 53844 51928 ne
rect 53844 51725 57700 51928
tri 57700 51725 57985 52010 sw
tri 57985 51725 58270 52010 ne
rect 58270 51916 59775 52010
tri 59775 51916 60059 52200 sw
tri 60059 51916 60343 52200 ne
rect 60343 51916 71000 52200
rect 58270 51725 60059 51916
rect 53844 51617 57985 51725
rect 49304 51593 53533 51617
rect 47146 51484 49017 51593
rect 45165 51193 46854 51484
rect 40754 51067 44872 51193
rect 36348 50932 40457 51067
rect 31822 50926 36060 50932
rect 27560 50650 31528 50926
rect 25489 50451 27270 50650
rect 23600 50360 25200 50451
tri 25200 50360 25291 50451 sw
tri 25489 50360 25580 50451 ne
rect 25580 50360 27270 50451
tri 27270 50360 27560 50650 sw
tri 27560 50360 27850 50650 ne
rect 27850 50632 31528 50650
tri 31528 50632 31822 50926 sw
tri 31822 50632 32116 50926 ne
rect 32116 50752 36060 50926
tri 36060 50752 36240 50932 sw
tri 36348 50752 36528 50932 ne
rect 36528 50770 40457 50932
tri 40457 50770 40754 51067 sw
tri 40754 50770 41051 51067 ne
rect 41051 50900 44872 51067
tri 44872 50900 45165 51193 sw
tri 45165 50900 45458 51193 ne
rect 45458 51192 46854 51193
tri 46854 51192 47146 51484 sw
tri 47146 51192 47438 51484 ne
rect 47438 51306 49017 51484
tri 49017 51306 49304 51593 sw
tri 49304 51306 49591 51593 ne
rect 49591 51306 53533 51593
tri 53533 51306 53844 51617 sw
tri 53844 51306 54155 51617 ne
rect 54155 51455 57985 51617
tri 57985 51455 58255 51725 sw
tri 58270 51455 58540 51725 ne
rect 58540 51632 60059 51725
tri 60059 51632 60343 51916 sw
tri 60343 51632 60627 51916 ne
rect 60627 51632 71000 51916
rect 58540 51455 60343 51632
rect 54155 51306 58255 51455
rect 47438 51192 49304 51306
rect 45458 50900 47146 51192
tri 47146 50900 47438 51192 sw
tri 47438 50900 47730 51192 ne
rect 47730 51019 49304 51192
tri 49304 51019 49591 51306 sw
tri 49591 51019 49878 51306 ne
rect 49878 51019 53844 51306
rect 47730 50900 49591 51019
rect 41051 50770 45165 50900
rect 36528 50752 40754 50770
rect 32116 50632 36240 50752
rect 27850 50360 31822 50632
rect 23600 50071 25291 50360
tri 25291 50071 25580 50360 sw
tri 25580 50071 25869 50360 ne
rect 25869 50071 27560 50360
tri 23400 49774 23600 49974 sw
tri 23600 49774 23897 50071 ne
rect 23897 49918 25580 50071
tri 25580 49918 25733 50071 sw
tri 25869 49918 26022 50071 ne
rect 26022 50070 27560 50071
tri 27560 50070 27850 50360 sw
tri 27850 50070 28140 50360 ne
rect 28140 50338 31822 50360
tri 31822 50338 32116 50632 sw
tri 32116 50338 32410 50632 ne
rect 32410 50464 36240 50632
tri 36240 50464 36528 50752 sw
tri 36528 50464 36816 50752 ne
rect 36816 50473 40754 50752
tri 40754 50473 41051 50770 sw
tri 41051 50473 41348 50770 ne
rect 41348 50607 45165 50770
tri 45165 50607 45458 50900 sw
tri 45458 50607 45751 50900 ne
rect 45751 50812 47438 50900
tri 47438 50812 47526 50900 sw
tri 47730 50812 47818 50900 ne
rect 47818 50812 49591 50900
rect 45751 50607 47526 50812
rect 41348 50473 45458 50607
rect 36816 50464 41051 50473
rect 32410 50338 36528 50464
rect 28140 50070 32116 50338
rect 26022 49974 27850 50070
tri 27850 49974 27946 50070 sw
tri 28140 49974 28236 50070 ne
rect 28236 50044 32116 50070
tri 32116 50044 32410 50338 sw
tri 32410 50044 32704 50338 ne
rect 32704 50176 36528 50338
tri 36528 50176 36816 50464 sw
tri 36816 50176 37104 50464 ne
rect 37104 50176 41051 50464
tri 41051 50176 41348 50473 sw
tri 41348 50176 41645 50473 ne
rect 41645 50314 45458 50473
tri 45458 50314 45751 50607 sw
tri 45751 50314 46044 50607 ne
rect 46044 50520 47526 50607
tri 47526 50520 47818 50812 sw
tri 47818 50520 48110 50812 ne
rect 48110 50807 49591 50812
tri 49591 50807 49803 51019 sw
tri 49878 50807 50090 51019 ne
rect 50090 50995 53844 51019
tri 53844 50995 54155 51306 sw
tri 54155 50995 54466 51306 ne
rect 54466 51170 58255 51306
tri 58255 51170 58540 51455 sw
tri 58540 51170 58825 51455 ne
rect 58825 51368 60343 51455
tri 60343 51368 60607 51632 sw
tri 60627 51368 60891 51632 ne
rect 60891 51368 71000 51632
rect 58825 51170 60607 51368
rect 54466 50995 58540 51170
rect 50090 50871 54155 50995
tri 54155 50871 54279 50995 sw
tri 54466 50871 54590 50995 ne
rect 54590 50885 58540 50995
tri 58540 50885 58825 51170 sw
tri 58825 50885 59110 51170 ne
rect 59110 51084 60607 51170
tri 60607 51084 60891 51368 sw
tri 60891 51084 61175 51368 ne
rect 61175 51084 71000 51368
rect 59110 50885 60891 51084
rect 54590 50871 58825 50885
rect 50090 50807 54279 50871
rect 48110 50520 49803 50807
tri 49803 50520 50090 50807 sw
tri 50090 50520 50377 50807 ne
rect 50377 50560 54279 50807
tri 54279 50560 54590 50871 sw
tri 54590 50560 54901 50871 ne
rect 54901 50600 58825 50871
tri 58825 50600 59110 50885 sw
tri 59110 50600 59395 50885 ne
rect 59395 50800 60891 50885
tri 60891 50800 61175 51084 sw
tri 61175 50800 61459 51084 ne
rect 61459 50800 71000 51084
rect 59395 50600 61175 50800
tri 61175 50600 61375 50800 sw
rect 54901 50560 59110 50600
rect 50377 50520 54590 50560
rect 46044 50314 47818 50520
rect 41645 50176 45751 50314
rect 32704 50044 36816 50176
rect 28236 49974 32410 50044
rect 26022 49918 27946 49974
rect 23897 49774 25733 49918
rect 20400 49477 23600 49774
tri 23600 49477 23897 49774 sw
tri 23897 49477 24194 49774 ne
rect 24194 49629 25733 49774
tri 25733 49629 26022 49918 sw
tri 26022 49629 26311 49918 ne
rect 26311 49684 27946 49918
tri 27946 49684 28236 49974 sw
tri 28236 49684 28526 49974 ne
rect 28526 49750 32410 49974
tri 32410 49750 32704 50044 sw
tri 32704 49750 32998 50044 ne
rect 32998 49888 36816 50044
tri 36816 49888 37104 50176 sw
tri 37104 49888 37392 50176 ne
rect 37392 49888 41348 50176
rect 32998 49750 37104 49888
rect 28526 49684 32704 49750
rect 26311 49629 28236 49684
rect 24194 49477 26022 49629
rect 20400 49354 23897 49477
tri 23897 49354 24020 49477 sw
tri 24194 49354 24317 49477 ne
rect 24317 49354 26022 49477
rect 20400 49057 24020 49354
tri 24020 49057 24317 49354 sw
tri 24317 49057 24614 49354 ne
rect 24614 49340 26022 49354
tri 26022 49340 26311 49629 sw
tri 26311 49340 26600 49629 ne
rect 26600 49394 28236 49629
tri 28236 49394 28526 49684 sw
tri 28526 49394 28816 49684 ne
rect 28816 49490 32704 49684
tri 32704 49490 32964 49750 sw
tri 32998 49490 33258 49750 ne
rect 33258 49600 37104 49750
tri 37104 49600 37392 49888 sw
tri 37392 49600 37680 49888 ne
rect 37680 49879 41348 49888
tri 41348 49879 41645 50176 sw
tri 41645 49879 41942 50176 ne
rect 41942 50021 45751 50176
tri 45751 50021 46044 50314 sw
tri 46044 50021 46337 50314 ne
rect 46337 50228 47818 50314
tri 47818 50228 48110 50520 sw
tri 48110 50228 48402 50520 ne
rect 48402 50249 50090 50520
tri 50090 50249 50361 50520 sw
tri 50377 50249 50648 50520 ne
rect 50648 50249 54590 50520
tri 54590 50249 54901 50560 sw
tri 54901 50249 55212 50560 ne
rect 55212 50315 59110 50560
tri 59110 50315 59395 50600 sw
tri 59395 50315 59680 50600 ne
rect 59680 50315 71000 50600
rect 55212 50249 59395 50315
rect 48402 50228 50361 50249
rect 46337 50021 48110 50228
rect 41942 49879 46044 50021
rect 37680 49726 41645 49879
tri 41645 49726 41798 49879 sw
tri 41942 49726 42095 49879 ne
rect 42095 49799 46044 49879
tri 46044 49799 46266 50021 sw
tri 46337 49799 46559 50021 ne
rect 46559 49936 48110 50021
tri 48110 49936 48402 50228 sw
tri 48402 49936 48694 50228 ne
rect 48694 49962 50361 50228
tri 50361 49962 50648 50249 sw
tri 50648 49962 50935 50249 ne
rect 50935 49962 54901 50249
rect 48694 49936 50648 49962
rect 46559 49799 48402 49936
rect 42095 49726 46266 49799
rect 37680 49600 41798 49726
rect 33258 49490 37392 49600
rect 28816 49394 32964 49490
rect 26600 49340 28526 49394
rect 24614 49057 26311 49340
rect 20400 48760 24317 49057
tri 24317 48760 24614 49057 sw
tri 24614 48760 24911 49057 ne
rect 24911 49051 26311 49057
tri 26311 49051 26600 49340 sw
tri 26600 49051 26889 49340 ne
rect 26889 49250 28526 49340
tri 28526 49250 28670 49394 sw
tri 28816 49250 28960 49394 ne
rect 28960 49250 32964 49394
rect 26889 49051 28670 49250
rect 24911 48762 26600 49051
tri 26600 48762 26889 49051 sw
tri 26889 48762 27178 49051 ne
rect 27178 48960 28670 49051
tri 28670 48960 28960 49250 sw
tri 28960 48960 29250 49250 ne
rect 29250 49196 32964 49250
tri 32964 49196 33258 49490 sw
tri 33258 49196 33552 49490 ne
rect 33552 49312 37392 49490
tri 37392 49312 37680 49600 sw
tri 37680 49312 37968 49600 ne
rect 37968 49429 41798 49600
tri 41798 49429 42095 49726 sw
tri 42095 49429 42392 49726 ne
rect 42392 49506 46266 49726
tri 46266 49506 46559 49799 sw
tri 46559 49506 46852 49799 ne
rect 46852 49644 48402 49799
tri 48402 49644 48694 49936 sw
tri 48694 49644 48986 49936 ne
rect 48986 49675 50648 49936
tri 50648 49675 50935 49962 sw
tri 50935 49675 51222 49962 ne
rect 51222 49938 54901 49962
tri 54901 49938 55212 50249 sw
tri 55212 49938 55523 50249 ne
rect 55523 50030 59395 50249
tri 59395 50030 59680 50315 sw
tri 59680 50030 59965 50315 ne
rect 59965 50030 71000 50315
rect 55523 49938 59680 50030
rect 51222 49675 55212 49938
rect 48986 49644 50935 49675
rect 46852 49506 48694 49644
rect 42392 49429 46559 49506
rect 37968 49312 42095 49429
rect 33552 49196 37680 49312
rect 29250 48960 33258 49196
rect 27178 48762 28960 48960
rect 24911 48760 26889 48762
rect 20400 48730 24614 48760
tri 20200 48448 20400 48648 sw
tri 20400 48448 20682 48730 ne
rect 20682 48671 24614 48730
tri 24614 48671 24703 48760 sw
tri 24911 48671 25000 48760 ne
rect 25000 48671 26889 48760
rect 20682 48448 24703 48671
rect 17200 48166 20400 48448
tri 20400 48166 20682 48448 sw
tri 20682 48166 20964 48448 ne
rect 20964 48374 24703 48448
tri 24703 48374 25000 48671 sw
tri 25000 48374 25297 48671 ne
rect 25297 48669 26889 48671
tri 26889 48669 26982 48762 sw
tri 27178 48669 27271 48762 ne
rect 27271 48670 28960 48762
tri 28960 48670 29250 48960 sw
tri 29250 48670 29540 48960 ne
rect 29540 48902 33258 48960
tri 33258 48902 33552 49196 sw
tri 33552 48902 33846 49196 ne
rect 33846 49024 37680 49196
tri 37680 49024 37968 49312 sw
tri 37968 49024 38256 49312 ne
rect 38256 49132 42095 49312
tri 42095 49132 42392 49429 sw
tri 42392 49132 42689 49429 ne
rect 42689 49213 46559 49429
tri 46559 49213 46852 49506 sw
tri 46852 49213 47145 49506 ne
rect 47145 49504 48694 49506
tri 48694 49504 48834 49644 sw
tri 48986 49504 49126 49644 ne
rect 49126 49504 50935 49644
rect 47145 49213 48834 49504
rect 42689 49132 46852 49213
rect 38256 49024 42392 49132
rect 33846 48902 37968 49024
rect 29540 48670 33552 48902
rect 27271 48669 29250 48670
rect 25297 48380 26982 48669
tri 26982 48380 27271 48669 sw
tri 27271 48380 27560 48669 ne
rect 27560 48380 29250 48669
tri 29250 48380 29540 48670 sw
tri 29540 48380 29830 48670 ne
rect 29830 48608 33552 48670
tri 33552 48608 33846 48902 sw
tri 33846 48608 34140 48902 ne
rect 34140 48736 37968 48902
tri 37968 48736 38256 49024 sw
tri 38256 48736 38544 49024 ne
rect 38544 48835 42392 49024
tri 42392 48835 42689 49132 sw
tri 42689 48835 42986 49132 ne
rect 42986 48920 46852 49132
tri 46852 48920 47145 49213 sw
tri 47145 48920 47438 49213 ne
rect 47438 49212 48834 49213
tri 48834 49212 49126 49504 sw
tri 49126 49212 49418 49504 ne
rect 49418 49419 50935 49504
tri 50935 49419 51191 49675 sw
tri 51222 49419 51478 49675 ne
rect 51478 49627 55212 49675
tri 55212 49627 55523 49938 sw
tri 55523 49627 55834 49938 ne
rect 55834 49770 59680 49938
tri 59680 49770 59940 50030 sw
tri 59965 49770 60225 50030 ne
rect 60225 49770 71000 50030
rect 55834 49627 59940 49770
rect 51478 49419 55523 49627
rect 49418 49212 51191 49419
rect 47438 48920 49126 49212
tri 49126 48920 49418 49212 sw
tri 49418 48920 49710 49212 ne
rect 49710 49132 51191 49212
tri 51191 49132 51478 49419 sw
tri 51478 49132 51765 49419 ne
rect 51765 49316 55523 49419
tri 55523 49316 55834 49627 sw
tri 55834 49316 56145 49627 ne
rect 56145 49485 59940 49627
tri 59940 49485 60225 49770 sw
tri 60225 49485 60510 49770 ne
rect 60510 49485 71000 49770
rect 56145 49316 60225 49485
rect 51765 49132 55834 49316
rect 49710 48920 51478 49132
rect 42986 48835 47145 48920
rect 38544 48736 42689 48835
rect 34140 48608 38256 48736
rect 29830 48380 33846 48608
rect 25297 48374 27271 48380
rect 20964 48166 25000 48374
rect 17200 47884 20682 48166
tri 20682 47884 20964 48166 sw
tri 20964 47884 21246 48166 ne
rect 21246 48077 25000 48166
tri 25000 48077 25297 48374 sw
tri 25297 48077 25594 48374 ne
rect 25594 48091 27271 48374
tri 27271 48091 27560 48380 sw
tri 27560 48091 27849 48380 ne
rect 27849 48091 29540 48380
rect 25594 48077 27560 48091
rect 21246 47884 25297 48077
rect 17200 47602 20964 47884
tri 20964 47602 21246 47884 sw
tri 21246 47602 21528 47884 ne
rect 21528 47780 25297 47884
tri 25297 47780 25594 48077 sw
tri 25594 47780 25891 48077 ne
rect 25891 47802 27560 48077
tri 27560 47802 27849 48091 sw
tri 27849 47802 28138 48091 ne
rect 28138 48090 29540 48091
tri 29540 48090 29830 48380 sw
tri 29830 48090 30120 48380 ne
rect 30120 48314 33846 48380
tri 33846 48314 34140 48608 sw
tri 34140 48314 34434 48608 ne
rect 34434 48448 38256 48608
tri 38256 48448 38544 48736 sw
tri 38544 48448 38832 48736 ne
rect 38832 48538 42689 48736
tri 42689 48538 42986 48835 sw
tri 42986 48538 43283 48835 ne
rect 43283 48627 47145 48835
tri 47145 48627 47438 48920 sw
tri 47438 48627 47731 48920 ne
rect 47731 48832 49418 48920
tri 49418 48832 49506 48920 sw
tri 49710 48832 49798 48920 ne
rect 49798 48845 51478 48920
tri 51478 48845 51765 49132 sw
tri 51765 48845 52052 49132 ne
rect 52052 49005 55834 49132
tri 55834 49005 56145 49316 sw
tri 56145 49005 56456 49316 ne
rect 56456 49200 60225 49316
tri 60225 49200 60510 49485 sw
tri 60510 49200 60795 49485 ne
rect 60795 49200 71000 49485
rect 56456 49005 60510 49200
rect 52052 48845 56145 49005
rect 49798 48832 51765 48845
rect 47731 48627 49506 48832
rect 43283 48538 47438 48627
rect 38832 48448 42986 48538
rect 34434 48416 38544 48448
tri 38544 48416 38576 48448 sw
tri 38832 48416 38864 48448 ne
rect 38864 48416 42986 48448
rect 34434 48314 38576 48416
rect 30120 48090 34140 48314
rect 28138 48020 29830 48090
tri 29830 48020 29900 48090 sw
tri 30120 48020 30190 48090 ne
rect 30190 48020 34140 48090
tri 34140 48020 34434 48314 sw
tri 34434 48020 34728 48314 ne
rect 34728 48128 38576 48314
tri 38576 48128 38864 48416 sw
tri 38864 48128 39152 48416 ne
rect 39152 48241 42986 48416
tri 42986 48241 43283 48538 sw
tri 43283 48241 43580 48538 ne
rect 43580 48334 47438 48538
tri 47438 48334 47731 48627 sw
tri 47731 48334 48024 48627 ne
rect 48024 48540 49506 48627
tri 49506 48540 49798 48832 sw
tri 49798 48540 50090 48832 ne
rect 50090 48827 51765 48832
tri 51765 48827 51783 48845 sw
tri 52052 48827 52070 48845 ne
rect 52070 48827 56145 48845
rect 50090 48540 51783 48827
tri 51783 48540 52070 48827 sw
tri 52070 48540 52357 48827 ne
rect 52357 48694 56145 48827
tri 56145 48694 56456 49005 sw
tri 56456 48694 56767 49005 ne
rect 56767 49000 60510 49005
tri 60510 49000 60710 49200 sw
rect 56767 48694 71000 49000
rect 52357 48608 56456 48694
tri 56456 48608 56542 48694 sw
tri 56767 48608 56853 48694 ne
rect 56853 48608 71000 48694
rect 52357 48540 56542 48608
rect 48024 48334 49798 48540
rect 43580 48241 47731 48334
rect 39152 48128 43283 48241
rect 34728 48020 38864 48128
rect 28138 47802 29900 48020
rect 25891 47780 27849 47802
rect 21528 47671 25594 47780
tri 25594 47671 25703 47780 sw
tri 25891 47671 26000 47780 ne
rect 26000 47671 27849 47780
rect 21528 47602 25703 47671
rect 17200 47404 21246 47602
tri 17000 47112 17200 47312 sw
tri 17200 47112 17492 47404 ne
rect 17492 47320 21246 47404
tri 21246 47320 21528 47602 sw
tri 21528 47320 21810 47602 ne
rect 21810 47374 25703 47602
tri 25703 47374 26000 47671 sw
tri 26000 47374 26297 47671 ne
rect 26297 47513 27849 47671
tri 27849 47513 28138 47802 sw
tri 28138 47513 28427 47802 ne
rect 28427 47730 29900 47802
tri 29900 47730 30190 48020 sw
tri 30190 47730 30480 48020 ne
rect 30480 47730 34434 48020
rect 28427 47513 30190 47730
rect 26297 47374 28138 47513
rect 21810 47320 26000 47374
rect 17492 47274 21528 47320
tri 21528 47274 21574 47320 sw
tri 21810 47274 21856 47320 ne
rect 21856 47274 26000 47320
rect 17492 47112 21574 47274
rect 14000 46908 17200 47112
tri 17200 46908 17404 47112 sw
tri 17492 46908 17696 47112 ne
rect 17696 46992 21574 47112
tri 21574 46992 21856 47274 sw
tri 21856 46992 22138 47274 ne
rect 22138 47077 26000 47274
tri 26000 47077 26297 47374 sw
tri 26297 47077 26594 47374 ne
rect 26594 47358 28138 47374
tri 28138 47358 28293 47513 sw
tri 28427 47358 28582 47513 ne
rect 28582 47440 30190 47513
tri 30190 47440 30480 47730 sw
tri 30480 47440 30770 47730 ne
rect 30770 47726 34434 47730
tri 34434 47726 34728 48020 sw
tri 34728 47726 35022 48020 ne
rect 35022 47840 38864 48020
tri 38864 47840 39152 48128 sw
tri 39152 47840 39440 48128 ne
rect 39440 47944 43283 48128
tri 43283 47944 43580 48241 sw
tri 43580 47944 43877 48241 ne
rect 43877 48041 47731 48241
tri 47731 48041 48024 48334 sw
tri 48024 48041 48317 48334 ne
rect 48317 48248 49798 48334
tri 49798 48248 50090 48540 sw
tri 50090 48248 50382 48540 ne
rect 50382 48253 52070 48540
tri 52070 48253 52357 48540 sw
tri 52357 48253 52644 48540 ne
rect 52644 48297 56542 48540
tri 56542 48297 56853 48608 sw
tri 56853 48297 57164 48608 ne
rect 57164 48297 71000 48608
rect 52644 48253 56853 48297
rect 50382 48248 52357 48253
rect 48317 48041 50090 48248
rect 43877 47944 48024 48041
rect 39440 47840 43580 47944
rect 35022 47726 39152 47840
rect 30770 47564 34728 47726
tri 34728 47564 34890 47726 sw
tri 35022 47564 35184 47726 ne
rect 35184 47564 39152 47726
rect 30770 47440 34890 47564
rect 28582 47358 30480 47440
rect 26594 47077 28293 47358
rect 22138 46992 26297 47077
rect 17696 46908 21856 46992
rect 14000 46616 17404 46908
tri 17404 46616 17696 46908 sw
tri 17696 46616 17988 46908 ne
rect 17988 46710 21856 46908
tri 21856 46710 22138 46992 sw
tri 22138 46710 22420 46992 ne
rect 22420 46780 26297 46992
tri 26297 46780 26594 47077 sw
tri 26594 46780 26891 47077 ne
rect 26891 47069 28293 47077
tri 28293 47069 28582 47358 sw
tri 28582 47069 28871 47358 ne
rect 28871 47266 30480 47358
tri 30480 47266 30654 47440 sw
tri 30770 47266 30944 47440 ne
rect 30944 47270 34890 47440
tri 34890 47270 35184 47564 sw
tri 35184 47270 35478 47564 ne
rect 35478 47552 39152 47564
tri 39152 47552 39440 47840 sw
tri 39440 47552 39728 47840 ne
rect 39728 47647 43580 47840
tri 43580 47647 43877 47944 sw
tri 43877 47647 44174 47944 ne
rect 44174 47819 48024 47944
tri 48024 47819 48246 48041 sw
tri 48317 47819 48539 48041 ne
rect 48539 47956 50090 48041
tri 50090 47956 50382 48248 sw
tri 50382 47956 50674 48248 ne
rect 50674 47966 52357 48248
tri 52357 47966 52644 48253 sw
tri 52644 47966 52931 48253 ne
rect 52931 47986 56853 48253
tri 56853 47986 57164 48297 sw
tri 57164 47986 57475 48297 ne
rect 57475 47986 71000 48297
rect 52931 47966 57164 47986
rect 50674 47956 52644 47966
rect 48539 47819 50382 47956
rect 44174 47647 48246 47819
rect 39728 47552 43877 47647
rect 35478 47270 39440 47552
rect 30944 47266 35184 47270
rect 28871 47069 30654 47266
rect 26891 46780 28582 47069
tri 28582 46780 28871 47069 sw
tri 28871 46780 29160 47069 ne
rect 29160 46976 30654 47069
tri 30654 46976 30944 47266 sw
tri 30944 46976 31234 47266 ne
rect 31234 46976 35184 47266
tri 35184 46976 35478 47270 sw
tri 35478 46976 35772 47270 ne
rect 35772 47264 39440 47270
tri 39440 47264 39728 47552 sw
tri 39728 47264 40016 47552 ne
rect 40016 47417 43877 47552
tri 43877 47417 44107 47647 sw
tri 44174 47417 44404 47647 ne
rect 44404 47526 48246 47647
tri 48246 47526 48539 47819 sw
tri 48539 47526 48832 47819 ne
rect 48832 47664 50382 47819
tri 50382 47664 50674 47956 sw
tri 50674 47664 50966 47956 ne
rect 50966 47679 52644 47956
tri 52644 47679 52931 47966 sw
tri 52931 47679 53218 47966 ne
rect 53218 47679 57164 47966
rect 50966 47664 52931 47679
rect 48832 47526 50674 47664
rect 44404 47417 48539 47526
rect 40016 47264 44107 47417
rect 35772 46976 39728 47264
tri 39728 46976 40016 47264 sw
tri 40016 46976 40304 47264 ne
rect 40304 47120 44107 47264
tri 44107 47120 44404 47417 sw
tri 44404 47120 44701 47417 ne
rect 44701 47233 48539 47417
tri 48539 47233 48832 47526 sw
tri 48832 47233 49125 47526 ne
rect 49125 47524 50674 47526
tri 50674 47524 50814 47664 sw
tri 50966 47524 51106 47664 ne
rect 51106 47627 52931 47664
tri 52931 47627 52983 47679 sw
tri 53218 47627 53270 47679 ne
rect 53270 47675 57164 47679
tri 57164 47675 57475 47986 sw
tri 57475 47675 57786 47986 ne
rect 57786 47675 71000 47986
rect 53270 47627 57475 47675
rect 51106 47524 52983 47627
rect 49125 47233 50814 47524
rect 44701 47120 48832 47233
rect 40304 46976 44404 47120
rect 29160 46780 30944 46976
rect 22420 46710 26594 46780
rect 17988 46616 22138 46710
rect 14000 46324 17696 46616
tri 17696 46324 17988 46616 sw
tri 17988 46324 18280 46616 ne
rect 18280 46428 22138 46616
tri 22138 46428 22420 46710 sw
tri 22420 46428 22702 46710 ne
rect 22702 46483 26594 46710
tri 26594 46483 26891 46780 sw
tri 26891 46483 27188 46780 ne
rect 27188 46689 28871 46780
tri 28871 46689 28962 46780 sw
tri 29160 46689 29251 46780 ne
rect 29251 46690 30944 46780
tri 30944 46690 31230 46976 sw
tri 31234 46690 31520 46976 ne
rect 31520 46690 35478 46976
rect 29251 46689 31230 46690
rect 27188 46483 28962 46689
rect 22702 46428 26891 46483
rect 18280 46324 22420 46428
rect 14000 46068 17988 46324
tri 14000 42497 17571 46068 ne
rect 17571 46032 17988 46068
tri 17988 46032 18280 46324 sw
tri 18280 46032 18572 46324 ne
rect 18572 46146 22420 46324
tri 22420 46146 22702 46428 sw
tri 22702 46146 22984 46428 ne
rect 22984 46186 26891 46428
tri 26891 46186 27188 46483 sw
tri 27188 46186 27485 46483 ne
rect 27485 46400 28962 46483
tri 28962 46400 29251 46689 sw
tri 29251 46400 29540 46689 ne
rect 29540 46400 31230 46689
tri 31230 46400 31520 46690 sw
tri 31520 46400 31810 46690 ne
rect 31810 46682 35478 46690
tri 35478 46682 35772 46976 sw
tri 35772 46682 36066 46976 ne
rect 36066 46688 40016 46976
tri 40016 46688 40304 46976 sw
tri 40304 46688 40592 46976 ne
rect 40592 46823 44404 46976
tri 44404 46823 44701 47120 sw
tri 44701 46823 44998 47120 ne
rect 44998 46940 48832 47120
tri 48832 46940 49125 47233 sw
tri 49125 46940 49418 47233 ne
rect 49418 47232 50814 47233
tri 50814 47232 51106 47524 sw
tri 51106 47232 51398 47524 ne
rect 51398 47340 52983 47524
tri 52983 47340 53270 47627 sw
tri 53270 47340 53557 47627 ne
rect 53557 47364 57475 47627
tri 57475 47364 57786 47675 sw
tri 57786 47364 58097 47675 ne
rect 58097 47364 71000 47675
rect 53557 47340 57786 47364
rect 51398 47232 53270 47340
rect 49418 46940 51106 47232
tri 51106 46940 51398 47232 sw
tri 51398 46940 51690 47232 ne
rect 51690 47053 53270 47232
tri 53270 47053 53557 47340 sw
tri 53557 47053 53844 47340 ne
rect 53844 47053 57786 47340
tri 57786 47053 58097 47364 sw
tri 58097 47053 58408 47364 ne
rect 58408 47053 71000 47364
rect 51690 46940 53557 47053
rect 44998 46823 49125 46940
rect 40592 46688 44701 46823
rect 36066 46682 40304 46688
rect 31810 46400 35772 46682
rect 27485 46186 29251 46400
rect 22984 46146 27188 46186
rect 18572 46032 22702 46146
rect 17571 45740 18280 46032
tri 18280 45740 18572 46032 sw
tri 18572 45740 18864 46032 ne
rect 18864 45864 22702 46032
tri 22702 45864 22984 46146 sw
tri 22984 45864 23266 46146 ne
rect 23266 45889 27188 46146
tri 27188 45889 27485 46186 sw
tri 27485 45889 27782 46186 ne
rect 27782 46111 29251 46186
tri 29251 46111 29540 46400 sw
tri 29540 46111 29829 46400 ne
rect 29829 46111 31520 46400
rect 27782 45889 29540 46111
rect 23266 45864 27485 45889
rect 18864 45740 22984 45864
rect 17571 45448 18572 45740
tri 18572 45448 18864 45740 sw
tri 18864 45448 19156 45740 ne
rect 19156 45582 22984 45740
tri 22984 45582 23266 45864 sw
tri 23266 45582 23548 45864 ne
rect 23548 45691 27485 45864
tri 27485 45691 27683 45889 sw
tri 27782 45691 27980 45889 ne
rect 27980 45822 29540 45889
tri 29540 45822 29829 46111 sw
tri 29829 45822 30118 46111 ne
rect 30118 46110 31520 46111
tri 31520 46110 31810 46400 sw
tri 31810 46110 32100 46400 ne
rect 32100 46388 35772 46400
tri 35772 46388 36066 46682 sw
tri 36066 46388 36360 46682 ne
rect 36360 46508 40304 46682
tri 40304 46508 40484 46688 sw
tri 40592 46508 40772 46688 ne
rect 40772 46526 44701 46688
tri 44701 46526 44998 46823 sw
tri 44998 46526 45295 46823 ne
rect 45295 46647 49125 46823
tri 49125 46647 49418 46940 sw
tri 49418 46647 49711 46940 ne
rect 49711 46852 51398 46940
tri 51398 46852 51486 46940 sw
tri 51690 46852 51778 46940 ne
rect 51778 46852 53557 46940
rect 49711 46647 51486 46852
rect 45295 46526 49418 46647
rect 40772 46508 44998 46526
rect 36360 46388 40484 46508
rect 32100 46110 36066 46388
rect 30118 45864 31810 46110
tri 31810 45864 32056 46110 sw
tri 32100 45864 32346 46110 ne
rect 32346 46094 36066 46110
tri 36066 46094 36360 46388 sw
tri 36360 46094 36654 46388 ne
rect 36654 46220 40484 46388
tri 40484 46220 40772 46508 sw
tri 40772 46220 41060 46508 ne
rect 41060 46229 44998 46508
tri 44998 46229 45295 46526 sw
tri 45295 46229 45592 46526 ne
rect 45592 46354 49418 46526
tri 49418 46354 49711 46647 sw
tri 49711 46354 50004 46647 ne
rect 50004 46560 51486 46647
tri 51486 46560 51778 46852 sw
tri 51778 46560 52070 46852 ne
rect 52070 46847 53557 46852
tri 53557 46847 53763 47053 sw
tri 53844 46847 54050 47053 ne
rect 54050 46847 58097 47053
rect 52070 46560 53763 46847
tri 53763 46560 54050 46847 sw
tri 54050 46560 54337 46847 ne
rect 54337 46742 58097 46847
tri 58097 46742 58408 47053 sw
tri 58408 46742 58719 47053 ne
rect 58719 46742 71000 47053
rect 54337 46622 58408 46742
tri 58408 46622 58528 46742 sw
tri 58719 46622 58839 46742 ne
rect 58839 46622 71000 46742
rect 54337 46560 58528 46622
rect 50004 46354 51778 46560
rect 45592 46229 49711 46354
rect 41060 46220 45295 46229
rect 36654 46094 40772 46220
rect 32346 45864 36360 46094
rect 30118 45822 32056 45864
rect 27980 45691 29829 45822
rect 23548 45582 27683 45691
rect 19156 45448 23266 45582
rect 17571 45168 18864 45448
tri 18864 45168 19144 45448 sw
tri 19156 45168 19436 45448 ne
rect 19436 45300 23266 45448
tri 23266 45300 23548 45582 sw
tri 23548 45300 23830 45582 ne
rect 23830 45394 27683 45582
tri 27683 45394 27980 45691 sw
tri 27980 45394 28277 45691 ne
rect 28277 45533 29829 45691
tri 29829 45533 30118 45822 sw
tri 30118 45533 30407 45822 ne
rect 30407 45574 32056 45822
tri 32056 45574 32346 45864 sw
tri 32346 45574 32636 45864 ne
rect 32636 45800 36360 45864
tri 36360 45800 36654 46094 sw
tri 36654 45800 36948 46094 ne
rect 36948 45932 40772 46094
tri 40772 45932 41060 46220 sw
tri 41060 45932 41348 46220 ne
rect 41348 45932 45295 46220
tri 45295 45932 45592 46229 sw
tri 45592 45932 45889 46229 ne
rect 45889 46061 49711 46229
tri 49711 46061 50004 46354 sw
tri 50004 46061 50297 46354 ne
rect 50297 46268 51778 46354
tri 51778 46268 52070 46560 sw
tri 52070 46268 52362 46560 ne
rect 52362 46273 54050 46560
tri 54050 46273 54337 46560 sw
tri 54337 46273 54624 46560 ne
rect 54624 46311 58528 46560
tri 58528 46311 58839 46622 sw
tri 58839 46311 59150 46622 ne
rect 59150 46311 71000 46622
rect 54624 46273 58839 46311
rect 52362 46268 54337 46273
rect 50297 46061 52070 46268
rect 45889 45932 50004 46061
rect 36948 45800 41060 45932
rect 32636 45574 36654 45800
rect 30407 45533 32346 45574
rect 28277 45394 30118 45533
rect 23830 45300 27980 45394
rect 19436 45168 23548 45300
rect 17571 44876 19144 45168
tri 19144 44876 19436 45168 sw
tri 19436 44876 19728 45168 ne
rect 19728 45018 23548 45168
tri 23548 45018 23830 45300 sw
tri 23830 45018 24112 45300 ne
rect 24112 45097 27980 45300
tri 27980 45097 28277 45394 sw
tri 28277 45097 28574 45394 ne
rect 28574 45378 30118 45394
tri 30118 45378 30273 45533 sw
tri 30407 45378 30562 45533 ne
rect 30562 45378 32346 45533
rect 28574 45097 30273 45378
rect 24112 45018 28277 45097
rect 19728 44876 23830 45018
rect 17571 44584 19436 44876
tri 19436 44584 19728 44876 sw
tri 19728 44584 20020 44876 ne
rect 20020 44736 23830 44876
tri 23830 44736 24112 45018 sw
tri 24112 44736 24394 45018 ne
rect 24394 44800 28277 45018
tri 28277 44800 28574 45097 sw
tri 28574 44800 28871 45097 ne
rect 28871 45089 30273 45097
tri 30273 45089 30562 45378 sw
tri 30562 45089 30851 45378 ne
rect 30851 45284 32346 45378
tri 32346 45284 32636 45574 sw
tri 32636 45284 32926 45574 ne
rect 32926 45506 36654 45574
tri 36654 45506 36948 45800 sw
tri 36948 45506 37242 45800 ne
rect 37242 45644 41060 45800
tri 41060 45644 41348 45932 sw
tri 41348 45644 41636 45932 ne
rect 41636 45644 45592 45932
rect 37242 45506 41348 45644
rect 32926 45284 36948 45506
rect 30851 45089 32636 45284
rect 28871 44800 30562 45089
tri 30562 44800 30851 45089 sw
tri 30851 44800 31140 45089 ne
rect 31140 45000 32636 45089
tri 32636 45000 32920 45284 sw
tri 32926 45000 33210 45284 ne
rect 33210 45246 36948 45284
tri 36948 45246 37208 45506 sw
tri 37242 45246 37502 45506 ne
rect 37502 45356 41348 45506
tri 41348 45356 41636 45644 sw
tri 41636 45356 41924 45644 ne
rect 41924 45635 45592 45644
tri 45592 45635 45889 45932 sw
tri 45889 45635 46186 45932 ne
rect 46186 45839 50004 45932
tri 50004 45839 50226 46061 sw
tri 50297 45839 50519 46061 ne
rect 50519 45976 52070 46061
tri 52070 45976 52362 46268 sw
tri 52362 45976 52654 46268 ne
rect 52654 46000 54337 46268
tri 54337 46000 54610 46273 sw
tri 54624 46000 54897 46273 ne
rect 54897 46000 58839 46273
tri 58839 46000 59150 46311 sw
tri 59150 46000 59461 46311 ne
rect 59461 46000 71000 46311
rect 52654 45976 54610 46000
rect 50519 45839 52362 45976
rect 46186 45635 50226 45839
rect 41924 45482 45889 45635
tri 45889 45482 46042 45635 sw
tri 46186 45482 46339 45635 ne
rect 46339 45546 50226 45635
tri 50226 45546 50519 45839 sw
tri 50519 45546 50812 45839 ne
rect 50812 45684 52362 45839
tri 52362 45684 52654 45976 sw
tri 52654 45684 52946 45976 ne
rect 52946 45713 54610 45976
tri 54610 45713 54897 46000 sw
tri 54897 45713 55184 46000 ne
rect 55184 45799 59150 46000
tri 59150 45799 59351 46000 sw
rect 55184 45739 71000 45799
rect 55184 45713 70613 45739
rect 52946 45684 54897 45713
rect 50812 45546 52654 45684
rect 46339 45482 50519 45546
rect 41924 45356 46042 45482
rect 37502 45246 41636 45356
rect 33210 45000 37208 45246
rect 31140 44800 32920 45000
rect 24394 44736 28574 44800
rect 20020 44584 24112 44736
rect 17571 44292 19728 44584
tri 19728 44292 20020 44584 sw
tri 20020 44292 20312 44584 ne
rect 20312 44454 24112 44584
tri 24112 44454 24394 44736 sw
tri 24394 44454 24676 44736 ne
rect 24676 44503 28574 44736
tri 28574 44503 28871 44800 sw
tri 28871 44503 29168 44800 ne
rect 29168 44709 30851 44800
tri 30851 44709 30942 44800 sw
tri 31140 44709 31231 44800 ne
rect 31231 44710 32920 44800
tri 32920 44710 33210 45000 sw
tri 33210 44710 33500 45000 ne
rect 33500 44952 37208 45000
tri 37208 44952 37502 45246 sw
tri 37502 44952 37796 45246 ne
rect 37796 45068 41636 45246
tri 41636 45068 41924 45356 sw
tri 41924 45068 42212 45356 ne
rect 42212 45185 46042 45356
tri 46042 45185 46339 45482 sw
tri 46339 45185 46636 45482 ne
rect 46636 45253 50519 45482
tri 50519 45253 50812 45546 sw
tri 50812 45253 51105 45546 ne
rect 51105 45472 52654 45546
tri 52654 45472 52866 45684 sw
tri 52946 45472 53158 45684 ne
rect 53158 45472 54897 45684
rect 51105 45253 52866 45472
rect 46636 45185 50812 45253
rect 42212 45068 46339 45185
rect 37796 44952 41924 45068
rect 33500 44710 37502 44952
rect 31231 44709 33210 44710
rect 29168 44503 30942 44709
rect 24676 44454 28871 44503
rect 20312 44292 24394 44454
rect 17571 44000 20020 44292
tri 20020 44000 20312 44292 sw
tri 20312 44000 20604 44292 ne
rect 20604 44172 24394 44292
tri 24394 44172 24676 44454 sw
tri 24676 44172 24958 44454 ne
rect 24958 44206 28871 44454
tri 28871 44206 29168 44503 sw
tri 29168 44206 29465 44503 ne
rect 29465 44420 30942 44503
tri 30942 44420 31231 44709 sw
tri 31231 44420 31520 44709 ne
rect 31520 44420 33210 44709
tri 33210 44420 33500 44710 sw
tri 33500 44420 33790 44710 ne
rect 33790 44658 37502 44710
tri 37502 44658 37796 44952 sw
tri 37796 44658 38090 44952 ne
rect 38090 44780 41924 44952
tri 41924 44780 42212 45068 sw
tri 42212 44780 42500 45068 ne
rect 42500 44888 46339 45068
tri 46339 44888 46636 45185 sw
tri 46636 44888 46933 45185 ne
rect 46933 44960 50812 45185
tri 50812 44960 51105 45253 sw
tri 51105 44960 51398 45253 ne
rect 51398 45180 52866 45253
tri 52866 45180 53158 45472 sw
tri 53158 45180 53450 45472 ne
rect 53450 45426 54897 45472
tri 54897 45426 55184 45713 sw
tri 55184 45426 55471 45713 ne
rect 55471 45426 70613 45713
rect 53450 45180 55184 45426
rect 51398 44960 53158 45180
rect 46933 44888 51105 44960
rect 42500 44780 46636 44888
rect 38090 44658 42212 44780
rect 33790 44420 37796 44658
rect 29465 44206 31231 44420
rect 24958 44172 29168 44206
rect 20604 44000 24676 44172
rect 17571 43708 20312 44000
tri 20312 43708 20604 44000 sw
tri 20604 43708 20896 44000 ne
rect 20896 43917 24676 44000
tri 24676 43917 24931 44172 sw
tri 24958 43917 25213 44172 ne
rect 25213 43917 29168 44172
rect 20896 43708 24931 43917
rect 17571 43416 20604 43708
tri 20604 43416 20896 43708 sw
tri 20896 43416 21188 43708 ne
rect 21188 43635 24931 43708
tri 24931 43635 25213 43917 sw
tri 25213 43635 25495 43917 ne
rect 25495 43909 29168 43917
tri 29168 43909 29465 44206 sw
tri 29465 43909 29762 44206 ne
rect 29762 44131 31231 44206
tri 31231 44131 31520 44420 sw
tri 31520 44131 31809 44420 ne
rect 31809 44131 33500 44420
rect 29762 43909 31520 44131
rect 25495 43711 29465 43909
tri 29465 43711 29663 43909 sw
tri 29762 43711 29960 43909 ne
rect 29960 43842 31520 43909
tri 31520 43842 31809 44131 sw
tri 31809 43842 32098 44131 ne
rect 32098 44130 33500 44131
tri 33500 44130 33790 44420 sw
tri 33790 44130 34080 44420 ne
rect 34080 44364 37796 44420
tri 37796 44364 38090 44658 sw
tri 38090 44364 38384 44658 ne
rect 38384 44492 42212 44658
tri 42212 44492 42500 44780 sw
tri 42500 44492 42788 44780 ne
rect 42788 44591 46636 44780
tri 46636 44591 46933 44888 sw
tri 46933 44591 47230 44888 ne
rect 47230 44667 51105 44888
tri 51105 44667 51398 44960 sw
tri 51398 44667 51691 44960 ne
rect 51691 44888 53158 44960
tri 53158 44888 53450 45180 sw
tri 53450 44888 53742 45180 ne
rect 53742 45175 55184 45180
tri 55184 45175 55435 45426 sw
tri 55471 45175 55722 45426 ne
rect 55722 45175 70613 45426
rect 53742 44888 55435 45175
tri 55435 44888 55722 45175 sw
tri 55722 44888 56009 45175 ne
rect 56009 44888 70613 45175
rect 51691 44872 53450 44888
tri 53450 44872 53466 44888 sw
tri 53742 44872 53758 44888 ne
rect 53758 44872 55722 44888
rect 51691 44667 53466 44872
rect 47230 44591 51398 44667
rect 42788 44492 46933 44591
rect 38384 44364 42500 44492
rect 34080 44130 38090 44364
rect 32098 44066 33790 44130
tri 33790 44066 33854 44130 sw
tri 34080 44066 34144 44130 ne
rect 34144 44070 38090 44130
tri 38090 44070 38384 44364 sw
tri 38384 44070 38678 44364 ne
rect 38678 44204 42500 44364
tri 42500 44204 42788 44492 sw
tri 42788 44204 43076 44492 ne
rect 43076 44294 46933 44492
tri 46933 44294 47230 44591 sw
tri 47230 44294 47527 44591 ne
rect 47527 44374 51398 44591
tri 51398 44374 51691 44667 sw
tri 51691 44374 51984 44667 ne
rect 51984 44580 53466 44667
tri 53466 44580 53758 44872 sw
tri 53758 44580 54050 44872 ne
rect 54050 44867 55722 44872
tri 55722 44867 55743 44888 sw
tri 56009 44867 56030 44888 ne
rect 56030 44867 70613 44888
rect 54050 44580 55743 44867
tri 55743 44580 56030 44867 sw
tri 56030 44580 56317 44867 ne
rect 56317 44580 70613 44867
rect 51984 44374 53758 44580
rect 47527 44294 51691 44374
rect 43076 44204 47230 44294
rect 38678 44172 42788 44204
tri 42788 44172 42820 44204 sw
tri 43076 44172 43108 44204 ne
rect 43108 44172 47230 44204
rect 38678 44070 42820 44172
rect 34144 44066 38384 44070
rect 32098 43842 33854 44066
rect 29960 43711 31809 43842
rect 25495 43635 29663 43711
rect 21188 43416 25213 43635
rect 17571 43248 20896 43416
tri 20896 43248 21064 43416 sw
tri 21188 43248 21356 43416 ne
rect 21356 43353 25213 43416
tri 25213 43353 25495 43635 sw
tri 25495 43353 25777 43635 ne
rect 25777 43414 29663 43635
tri 29663 43414 29960 43711 sw
tri 29960 43414 30257 43711 ne
rect 30257 43553 31809 43711
tri 31809 43553 32098 43842 sw
tri 32098 43553 32387 43842 ne
rect 32387 43776 33854 43842
tri 33854 43776 34144 44066 sw
tri 34144 43776 34434 44066 ne
rect 34434 43776 38384 44066
tri 38384 43776 38678 44070 sw
tri 38678 43776 38972 44070 ne
rect 38972 43884 42820 44070
tri 42820 43884 43108 44172 sw
tri 43108 43884 43396 44172 ne
rect 43396 43997 47230 44172
tri 47230 43997 47527 44294 sw
tri 47527 43997 47824 44294 ne
rect 47824 44081 51691 44294
tri 51691 44081 51984 44374 sw
tri 51984 44081 52277 44374 ne
rect 52277 44288 53758 44374
tri 53758 44288 54050 44580 sw
tri 54050 44288 54342 44580 ne
rect 54342 44293 56030 44580
tri 56030 44293 56317 44580 sw
tri 56317 44293 56604 44580 ne
rect 56604 44293 70613 44580
rect 54342 44288 56317 44293
rect 52277 44081 54050 44288
rect 47824 43997 51984 44081
rect 43396 43884 47527 43997
rect 38972 43776 43108 43884
rect 32387 43553 34144 43776
rect 30257 43414 32098 43553
rect 25777 43353 29960 43414
rect 21356 43248 25495 43353
rect 17571 42956 21064 43248
tri 21064 42956 21356 43248 sw
tri 21356 42956 21648 43248 ne
rect 21648 43071 25495 43248
tri 25495 43071 25777 43353 sw
tri 25777 43071 26059 43353 ne
rect 26059 43117 29960 43353
tri 29960 43117 30257 43414 sw
tri 30257 43117 30554 43414 ne
rect 30554 43398 32098 43414
tri 32098 43398 32253 43553 sw
tri 32387 43398 32542 43553 ne
rect 32542 43486 34144 43553
tri 34144 43486 34434 43776 sw
tri 34434 43486 34724 43776 ne
rect 34724 43486 38678 43776
rect 32542 43398 34434 43486
rect 30554 43117 32253 43398
rect 26059 43071 30257 43117
rect 21648 42956 25777 43071
rect 17571 42664 21356 42956
tri 21356 42664 21648 42956 sw
tri 21648 42664 21940 42956 ne
rect 21940 42789 25777 42956
tri 25777 42789 26059 43071 sw
tri 26059 42789 26341 43071 ne
rect 26341 42820 30257 43071
tri 30257 42820 30554 43117 sw
tri 30554 42820 30851 43117 ne
rect 30851 43109 32253 43117
tri 32253 43109 32542 43398 sw
tri 32542 43109 32831 43398 ne
rect 32831 43196 34434 43398
tri 34434 43196 34724 43486 sw
tri 34724 43196 35014 43486 ne
rect 35014 43482 38678 43486
tri 38678 43482 38972 43776 sw
tri 38972 43482 39266 43776 ne
rect 39266 43596 43108 43776
tri 43108 43596 43396 43884 sw
tri 43396 43596 43684 43884 ne
rect 43684 43700 47527 43884
tri 47527 43700 47824 43997 sw
tri 47824 43700 48121 43997 ne
rect 48121 43859 51984 43997
tri 51984 43859 52206 44081 sw
tri 52277 43859 52499 44081 ne
rect 52499 43996 54050 44081
tri 54050 43996 54342 44288 sw
tri 54342 43996 54634 44288 ne
rect 54634 44006 56317 44288
tri 56317 44006 56604 44293 sw
tri 56604 44006 56891 44293 ne
rect 56891 44006 70613 44293
rect 54634 43996 56604 44006
rect 52499 43859 54342 43996
rect 48121 43700 52206 43859
rect 43684 43596 47824 43700
rect 39266 43482 43396 43596
rect 35014 43320 38972 43482
tri 38972 43320 39134 43482 sw
tri 39266 43320 39428 43482 ne
rect 39428 43320 43396 43482
rect 35014 43196 39134 43320
rect 32831 43109 34724 43196
rect 30851 42820 32542 43109
tri 32542 42820 32831 43109 sw
tri 32831 42820 33120 43109 ne
rect 33120 43020 34724 43109
tri 34724 43020 34900 43196 sw
tri 35014 43020 35190 43196 ne
rect 35190 43026 39134 43196
tri 39134 43026 39428 43320 sw
tri 39428 43026 39722 43320 ne
rect 39722 43308 43396 43320
tri 43396 43308 43684 43596 sw
tri 43684 43308 43972 43596 ne
rect 43972 43403 47824 43596
tri 47824 43403 48121 43700 sw
tri 48121 43403 48418 43700 ne
rect 48418 43566 52206 43700
tri 52206 43566 52499 43859 sw
tri 52499 43566 52792 43859 ne
rect 52792 43704 54342 43859
tri 54342 43704 54634 43996 sw
tri 54634 43704 54926 43996 ne
rect 54926 43719 56604 43996
tri 56604 43719 56891 44006 sw
tri 56891 43719 57178 44006 ne
rect 57178 43719 70613 44006
rect 54926 43704 56891 43719
rect 52792 43676 54634 43704
tri 54634 43676 54662 43704 sw
tri 54926 43676 54954 43704 ne
rect 54954 43676 56891 43704
rect 52792 43566 54662 43676
rect 48418 43403 52499 43566
rect 43972 43308 48121 43403
rect 39722 43026 43684 43308
rect 35190 43020 39428 43026
rect 33120 42820 34900 43020
rect 26341 42789 30554 42820
rect 21940 42664 26059 42789
rect 17571 42497 21648 42664
tri 17571 38420 21648 42497 ne
tri 21648 42372 21940 42664 sw
tri 21940 42372 22232 42664 ne
rect 22232 42507 26059 42664
tri 26059 42507 26341 42789 sw
tri 26341 42507 26623 42789 ne
rect 26623 42523 30554 42789
tri 30554 42523 30851 42820 sw
tri 30851 42523 31148 42820 ne
rect 31148 42729 32831 42820
tri 32831 42729 32922 42820 sw
tri 33120 42729 33211 42820 ne
rect 33211 42730 34900 42820
tri 34900 42730 35190 43020 sw
tri 35190 42730 35480 43020 ne
rect 35480 42732 39428 43020
tri 39428 42732 39722 43026 sw
tri 39722 42732 40016 43026 ne
rect 40016 43020 43684 43026
tri 43684 43020 43972 43308 sw
tri 43972 43020 44260 43308 ne
rect 44260 43173 48121 43308
tri 48121 43173 48351 43403 sw
tri 48418 43173 48648 43403 ne
rect 48648 43273 52499 43403
tri 52499 43273 52792 43566 sw
tri 52792 43273 53085 43566 ne
rect 53085 43384 54662 43566
tri 54662 43384 54954 43676 sw
tri 54954 43384 55246 43676 ne
rect 55246 43461 56891 43676
tri 56891 43461 57149 43719 sw
tri 57178 43461 57436 43719 ne
rect 57436 43461 70613 43719
rect 55246 43384 57149 43461
rect 53085 43273 54954 43384
rect 48648 43173 52792 43273
rect 44260 43020 48351 43173
rect 40016 42732 43972 43020
tri 43972 42732 44260 43020 sw
tri 44260 42732 44548 43020 ne
rect 44548 42876 48351 43020
tri 48351 42876 48648 43173 sw
tri 48648 42876 48945 43173 ne
rect 48945 42980 52792 43173
tri 52792 42980 53085 43273 sw
tri 53085 42980 53378 43273 ne
rect 53378 43092 54954 43273
tri 54954 43092 55246 43384 sw
tri 55246 43092 55538 43384 ne
rect 55538 43174 57149 43384
tri 57149 43174 57436 43461 sw
tri 57436 43174 57723 43461 ne
rect 57723 43174 70613 43461
rect 55538 43092 57436 43174
rect 53378 42980 55246 43092
rect 48945 42876 53085 42980
rect 44548 42732 48648 42876
rect 35480 42730 39722 42732
rect 33211 42729 35190 42730
rect 31148 42523 32922 42729
rect 26623 42507 30851 42523
rect 22232 42372 26341 42507
rect 21648 42080 21940 42372
tri 21940 42080 22232 42372 sw
tri 22232 42080 22524 42372 ne
rect 22524 42225 26341 42372
tri 26341 42225 26623 42507 sw
tri 26623 42225 26905 42507 ne
rect 26905 42226 30851 42507
tri 30851 42226 31148 42523 sw
tri 31148 42226 31445 42523 ne
rect 31445 42440 32922 42523
tri 32922 42440 33211 42729 sw
tri 33211 42440 33500 42729 ne
rect 33500 42440 35190 42729
tri 35190 42440 35480 42730 sw
tri 35480 42440 35770 42730 ne
rect 35770 42440 39722 42730
rect 31445 42226 33211 42440
rect 26905 42225 31148 42226
rect 22524 42184 26623 42225
tri 26623 42184 26664 42225 sw
tri 26905 42184 26946 42225 ne
rect 26946 42184 31148 42225
rect 22524 42080 26664 42184
rect 21648 41788 22232 42080
tri 22232 41788 22524 42080 sw
tri 22524 41788 22816 42080 ne
rect 22816 41902 26664 42080
tri 26664 41902 26946 42184 sw
tri 26946 41902 27228 42184 ne
rect 27228 41929 31148 42184
tri 31148 41929 31445 42226 sw
tri 31445 41929 31742 42226 ne
rect 31742 42151 33211 42226
tri 33211 42151 33500 42440 sw
tri 33500 42151 33789 42440 ne
rect 33789 42151 35480 42440
rect 31742 41929 33500 42151
rect 27228 41902 31445 41929
rect 22816 41788 26946 41902
rect 21648 41496 22524 41788
tri 22524 41496 22816 41788 sw
tri 22816 41496 23108 41788 ne
rect 23108 41620 26946 41788
tri 26946 41620 27228 41902 sw
tri 27228 41620 27510 41902 ne
rect 27510 41731 31445 41902
tri 31445 41731 31643 41929 sw
tri 31742 41731 31940 41929 ne
rect 31940 41862 33500 41929
tri 33500 41862 33789 42151 sw
tri 33789 41862 34078 42151 ne
rect 34078 42150 35480 42151
tri 35480 42150 35770 42440 sw
tri 35770 42150 36060 42440 ne
rect 36060 42438 39722 42440
tri 39722 42438 40016 42732 sw
tri 40016 42438 40310 42732 ne
rect 40310 42444 44260 42732
tri 44260 42444 44548 42732 sw
tri 44548 42444 44836 42732 ne
rect 44836 42579 48648 42732
tri 48648 42579 48945 42876 sw
tri 48945 42579 49242 42876 ne
rect 49242 42687 53085 42876
tri 53085 42687 53378 42980 sw
tri 53378 42687 53671 42980 ne
rect 53671 42800 55246 42980
tri 55246 42800 55538 43092 sw
tri 55538 42800 55830 43092 ne
rect 55830 42887 57436 43092
tri 57436 42887 57723 43174 sw
tri 57723 42887 58010 43174 ne
rect 58010 42887 70613 43174
rect 55830 42800 57723 42887
rect 53671 42687 55538 42800
rect 49242 42579 53378 42687
rect 44836 42444 48945 42579
rect 40310 42438 44548 42444
rect 36060 42150 40016 42438
rect 34078 41910 35770 42150
tri 35770 41910 36010 42150 sw
tri 36060 41910 36300 42150 ne
rect 36300 42144 40016 42150
tri 40016 42144 40310 42438 sw
tri 40310 42144 40604 42438 ne
rect 40604 42264 44548 42438
tri 44548 42264 44728 42444 sw
tri 44836 42264 45016 42444 ne
rect 45016 42282 48945 42444
tri 48945 42282 49242 42579 sw
tri 49242 42282 49539 42579 ne
rect 49539 42394 53378 42579
tri 53378 42394 53671 42687 sw
tri 53671 42394 53964 42687 ne
rect 53964 42600 55538 42687
tri 55538 42600 55738 42800 sw
tri 55830 42600 56030 42800 ne
rect 56030 42600 57723 42800
tri 57723 42600 58010 42887 sw
tri 58010 42800 58097 42887 ne
rect 58097 42875 70613 42887
rect 70669 42875 71000 45739
rect 58097 42800 71000 42875
rect 53964 42394 55738 42600
rect 49539 42282 53671 42394
rect 45016 42264 49242 42282
rect 40604 42144 44728 42264
rect 36300 41910 40310 42144
rect 34078 41862 36010 41910
rect 31940 41731 33789 41862
rect 27510 41620 31643 41731
rect 23108 41496 27228 41620
rect 21648 41204 22816 41496
tri 22816 41204 23108 41496 sw
tri 23108 41204 23400 41496 ne
rect 23400 41338 27228 41496
tri 27228 41338 27510 41620 sw
tri 27510 41338 27792 41620 ne
rect 27792 41434 31643 41620
tri 31643 41434 31940 41731 sw
tri 31940 41434 32237 41731 ne
rect 32237 41573 33789 41731
tri 33789 41573 34078 41862 sw
tri 34078 41573 34367 41862 ne
rect 34367 41620 36010 41862
tri 36010 41620 36300 41910 sw
tri 36300 41620 36590 41910 ne
rect 36590 41850 40310 41910
tri 40310 41850 40604 42144 sw
tri 40604 41850 40898 42144 ne
rect 40898 41976 44728 42144
tri 44728 41976 45016 42264 sw
tri 45016 41976 45304 42264 ne
rect 45304 41985 49242 42264
tri 49242 41985 49539 42282 sw
tri 49539 41985 49836 42282 ne
rect 49836 42101 53671 42282
tri 53671 42101 53964 42394 sw
tri 53964 42101 54257 42394 ne
rect 54257 42308 55738 42394
tri 55738 42308 56030 42600 sw
tri 56030 42308 56322 42600 ne
rect 56322 42497 71000 42600
rect 56322 42308 70613 42497
rect 54257 42101 56030 42308
rect 49836 41985 53964 42101
rect 45304 41976 49539 41985
rect 40898 41850 45016 41976
rect 36590 41620 40604 41850
rect 34367 41573 36300 41620
rect 32237 41434 34078 41573
rect 27792 41338 31940 41434
rect 23400 41204 27510 41338
rect 21648 40924 23108 41204
tri 23108 40924 23388 41204 sw
tri 23400 40924 23680 41204 ne
rect 23680 41056 27510 41204
tri 27510 41056 27792 41338 sw
tri 27792 41056 28074 41338 ne
rect 28074 41137 31940 41338
tri 31940 41137 32237 41434 sw
tri 32237 41137 32534 41434 ne
rect 32534 41297 34078 41434
tri 34078 41297 34354 41573 sw
tri 34367 41297 34643 41573 ne
rect 34643 41330 36300 41573
tri 36300 41330 36590 41620 sw
tri 36590 41330 36880 41620 ne
rect 36880 41556 40604 41620
tri 40604 41556 40898 41850 sw
tri 40898 41556 41192 41850 ne
rect 41192 41688 45016 41850
tri 45016 41688 45304 41976 sw
tri 45304 41688 45592 41976 ne
rect 45592 41688 49539 41976
tri 49539 41688 49836 41985 sw
tri 49836 41688 50133 41985 ne
rect 50133 41879 53964 41985
tri 53964 41879 54186 42101 sw
tri 54257 41879 54479 42101 ne
rect 54479 42016 56030 42101
tri 56030 42016 56322 42308 sw
tri 56322 42016 56614 42308 ne
rect 56614 42016 70613 42308
rect 54479 41879 56322 42016
rect 50133 41688 54186 41879
rect 41192 41556 45304 41688
rect 36880 41330 40898 41556
rect 34643 41297 36590 41330
rect 32534 41137 34354 41297
rect 28074 41056 32237 41137
rect 23680 40924 27792 41056
rect 21648 40632 23388 40924
tri 23388 40632 23680 40924 sw
tri 23680 40632 23972 40924 ne
rect 23972 40774 27792 40924
tri 27792 40774 28074 41056 sw
tri 28074 40774 28356 41056 ne
rect 28356 40840 32237 41056
tri 32237 40840 32534 41137 sw
tri 32534 40840 32831 41137 ne
rect 32831 41129 34354 41137
tri 34354 41129 34522 41297 sw
tri 34643 41129 34811 41297 ne
rect 34811 41129 36590 41297
rect 32831 40840 34522 41129
tri 34522 40840 34811 41129 sw
tri 34811 40840 35100 41129 ne
rect 35100 41040 36590 41129
tri 36590 41040 36880 41330 sw
tri 36880 41040 37170 41330 ne
rect 37170 41262 40898 41330
tri 40898 41262 41192 41556 sw
tri 41192 41262 41486 41556 ne
rect 41486 41400 45304 41556
tri 45304 41400 45592 41688 sw
tri 45592 41400 45880 41688 ne
rect 45880 41400 49836 41688
rect 41486 41262 45592 41400
rect 37170 41040 41192 41262
rect 35100 40840 36880 41040
rect 28356 40774 32534 40840
rect 23972 40632 28074 40774
rect 21648 40340 23680 40632
tri 23680 40340 23972 40632 sw
tri 23972 40340 24264 40632 ne
rect 24264 40492 28074 40632
tri 28074 40492 28356 40774 sw
tri 28356 40492 28638 40774 ne
rect 28638 40543 32534 40774
tri 32534 40543 32831 40840 sw
tri 32831 40543 33128 40840 ne
rect 33128 40749 34811 40840
tri 34811 40749 34902 40840 sw
tri 35100 40749 35191 40840 ne
rect 35191 40750 36880 40840
tri 36880 40750 37170 41040 sw
tri 37170 40750 37460 41040 ne
rect 37460 41002 41192 41040
tri 41192 41002 41452 41262 sw
tri 41486 41002 41746 41262 ne
rect 41746 41112 45592 41262
tri 45592 41112 45880 41400 sw
tri 45880 41112 46168 41400 ne
rect 46168 41391 49836 41400
tri 49836 41391 50133 41688 sw
tri 50133 41391 50430 41688 ne
rect 50430 41586 54186 41688
tri 54186 41586 54479 41879 sw
tri 54479 41586 54772 41879 ne
rect 54772 41784 56322 41879
tri 56322 41784 56554 42016 sw
tri 56614 41784 56846 42016 ne
rect 56846 41784 70613 42016
rect 54772 41586 56554 41784
rect 50430 41391 54479 41586
rect 46168 41238 50133 41391
tri 50133 41238 50286 41391 sw
tri 50430 41238 50583 41391 ne
rect 50583 41293 54479 41391
tri 54479 41293 54772 41586 sw
tri 54772 41293 55065 41586 ne
rect 55065 41492 56554 41586
tri 56554 41492 56846 41784 sw
tri 56846 41492 57138 41784 ne
rect 57138 41492 70613 41784
rect 55065 41293 56846 41492
rect 50583 41238 54772 41293
rect 46168 41112 50286 41238
rect 41746 41002 45880 41112
rect 37460 40750 41452 41002
rect 35191 40749 37170 40750
rect 33128 40543 34902 40749
rect 28638 40492 32831 40543
rect 24264 40340 28356 40492
rect 21648 40048 23972 40340
tri 23972 40048 24264 40340 sw
tri 24264 40048 24556 40340 ne
rect 24556 40210 28356 40340
tri 28356 40210 28638 40492 sw
tri 28638 40210 28920 40492 ne
rect 28920 40246 32831 40492
tri 32831 40246 33128 40543 sw
tri 33128 40246 33425 40543 ne
rect 33425 40460 34902 40543
tri 34902 40460 35191 40749 sw
tri 35191 40460 35480 40749 ne
rect 35480 40460 37170 40749
tri 37170 40460 37460 40750 sw
tri 37460 40460 37750 40750 ne
rect 37750 40708 41452 40750
tri 41452 40708 41746 41002 sw
tri 41746 40708 42040 41002 ne
rect 42040 40824 45880 41002
tri 45880 40824 46168 41112 sw
tri 46168 40824 46456 41112 ne
rect 46456 40941 50286 41112
tri 50286 40941 50583 41238 sw
tri 50583 40941 50880 41238 ne
rect 50880 41000 54772 41238
tri 54772 41000 55065 41293 sw
tri 55065 41000 55358 41293 ne
rect 55358 41200 56846 41293
tri 56846 41200 57138 41492 sw
tri 57138 41200 57430 41492 ne
rect 57430 41297 70613 41492
rect 70669 41297 71000 42497
rect 57430 41200 71000 41297
rect 55358 41000 57138 41200
tri 57138 41000 57338 41200 sw
rect 50880 40941 55065 41000
rect 46456 40824 50583 40941
rect 42040 40708 46168 40824
rect 37750 40460 41746 40708
rect 33425 40246 35191 40460
rect 28920 40210 33128 40246
rect 24556 40048 28638 40210
rect 21648 39756 24264 40048
tri 24264 39756 24556 40048 sw
tri 24556 39756 24848 40048 ne
rect 24848 39928 28638 40048
tri 28638 39928 28920 40210 sw
tri 28920 39928 29202 40210 ne
rect 29202 39949 33128 40210
tri 33128 39949 33425 40246 sw
tri 33425 39949 33722 40246 ne
rect 33722 40171 35191 40246
tri 35191 40171 35480 40460 sw
tri 35480 40171 35769 40460 ne
rect 35769 40171 37460 40460
rect 33722 39949 35480 40171
rect 29202 39928 33425 39949
rect 24848 39830 28920 39928
tri 28920 39830 29018 39928 sw
tri 29202 39830 29300 39928 ne
rect 29300 39830 33425 39928
rect 24848 39756 29018 39830
rect 21648 39464 24556 39756
tri 24556 39464 24848 39756 sw
tri 24848 39464 25140 39756 ne
rect 25140 39548 29018 39756
tri 29018 39548 29300 39830 sw
tri 29300 39548 29582 39830 ne
rect 29582 39751 33425 39830
tri 33425 39751 33623 39949 sw
tri 33722 39751 33920 39949 ne
rect 33920 39882 35480 39949
tri 35480 39882 35769 40171 sw
tri 35769 39882 36058 40171 ne
rect 36058 40170 37460 40171
tri 37460 40170 37750 40460 sw
tri 37750 40170 38040 40460 ne
rect 38040 40414 41746 40460
tri 41746 40414 42040 40708 sw
tri 42040 40414 42334 40708 ne
rect 42334 40536 46168 40708
tri 46168 40536 46456 40824 sw
tri 46456 40536 46744 40824 ne
rect 46744 40644 50583 40824
tri 50583 40644 50880 40941 sw
tri 50880 40644 51177 40941 ne
rect 51177 40707 55065 40941
tri 55065 40707 55358 41000 sw
tri 55358 40707 55651 41000 ne
rect 55651 40707 71000 41000
rect 51177 40644 55358 40707
rect 46744 40536 50880 40644
rect 42334 40414 46456 40536
rect 38040 40170 42040 40414
rect 36058 39882 37750 40170
rect 33920 39751 35769 39882
rect 29582 39548 33623 39751
rect 25140 39464 29300 39548
rect 21648 39172 24848 39464
tri 24848 39172 25140 39464 sw
tri 25140 39172 25432 39464 ne
rect 25432 39266 29300 39464
tri 29300 39266 29582 39548 sw
tri 29582 39266 29864 39548 ne
rect 29864 39454 33623 39548
tri 33623 39454 33920 39751 sw
tri 33920 39454 34217 39751 ne
rect 34217 39593 35769 39751
tri 35769 39593 36058 39882 sw
tri 36058 39593 36347 39882 ne
rect 36347 39880 37750 39882
tri 37750 39880 38040 40170 sw
tri 38040 39880 38330 40170 ne
rect 38330 40120 42040 40170
tri 42040 40120 42334 40414 sw
tri 42334 40120 42628 40414 ne
rect 42628 40248 46456 40414
tri 46456 40248 46744 40536 sw
tri 46744 40248 47032 40536 ne
rect 47032 40347 50880 40536
tri 50880 40347 51177 40644 sw
tri 51177 40347 51474 40644 ne
rect 51474 40414 55358 40644
tri 55358 40414 55651 40707 sw
tri 55651 40414 55944 40707 ne
rect 55944 40414 71000 40707
rect 51474 40347 55651 40414
rect 47032 40248 51177 40347
rect 42628 40120 46744 40248
rect 38330 39880 42334 40120
rect 36347 39822 38040 39880
tri 38040 39822 38098 39880 sw
tri 38330 39822 38388 39880 ne
rect 38388 39826 42334 39880
tri 42334 39826 42628 40120 sw
tri 42628 39826 42922 40120 ne
rect 42922 39960 46744 40120
tri 46744 39960 47032 40248 sw
tri 47032 39960 47320 40248 ne
rect 47320 40050 51177 40248
tri 51177 40050 51474 40347 sw
tri 51474 40050 51771 40347 ne
rect 51771 40186 55651 40347
tri 55651 40186 55879 40414 sw
tri 55944 40186 56172 40414 ne
rect 56172 40186 71000 40414
rect 51771 40050 55879 40186
rect 47320 39960 51474 40050
rect 42922 39928 47032 39960
tri 47032 39928 47064 39960 sw
tri 47320 39928 47352 39960 ne
rect 47352 39928 51474 39960
rect 42922 39826 47064 39928
rect 38388 39822 42628 39826
rect 36347 39593 38098 39822
rect 34217 39454 36058 39593
rect 29864 39266 33920 39454
rect 25432 39172 29582 39266
rect 21648 39004 25140 39172
tri 25140 39004 25308 39172 sw
tri 25432 39004 25600 39172 ne
rect 25600 39004 29582 39172
rect 21648 38712 25308 39004
tri 25308 38712 25600 39004 sw
tri 25600 38712 25892 39004 ne
rect 25892 38984 29582 39004
tri 29582 38984 29864 39266 sw
tri 29864 38984 30146 39266 ne
rect 30146 39157 33920 39266
tri 33920 39157 34217 39454 sw
tri 34217 39157 34514 39454 ne
rect 34514 39332 36058 39454
tri 36058 39332 36319 39593 sw
tri 36347 39332 36608 39593 ne
rect 36608 39532 38098 39593
tri 38098 39532 38388 39822 sw
tri 38388 39532 38678 39822 ne
rect 38678 39532 42628 39822
tri 42628 39532 42922 39826 sw
tri 42922 39532 43216 39826 ne
rect 43216 39640 47064 39826
tri 47064 39640 47352 39928 sw
tri 47352 39640 47640 39928 ne
rect 47640 39753 51474 39928
tri 51474 39753 51771 40050 sw
tri 51771 39753 52068 40050 ne
rect 52068 39893 55879 40050
tri 55879 39893 56172 40186 sw
tri 56172 39893 56465 40186 ne
rect 56465 39893 71000 40186
rect 52068 39753 56172 39893
rect 47640 39640 51771 39753
rect 43216 39532 47352 39640
rect 36608 39332 38388 39532
rect 34514 39157 36319 39332
rect 30146 38984 34217 39157
rect 25892 38712 29864 38984
rect 21648 38420 25600 38712
tri 25600 38420 25892 38712 sw
tri 25892 38420 26184 38712 ne
rect 26184 38702 29864 38712
tri 29864 38702 30146 38984 sw
tri 30146 38702 30428 38984 ne
rect 30428 38860 34217 38984
tri 34217 38860 34514 39157 sw
tri 34514 38860 34811 39157 ne
rect 34811 39149 36319 39157
tri 36319 39149 36502 39332 sw
tri 36608 39149 36791 39332 ne
rect 36791 39242 38388 39332
tri 38388 39242 38678 39532 sw
tri 38678 39242 38968 39532 ne
rect 38968 39242 42922 39532
rect 36791 39149 38678 39242
rect 34811 38860 36502 39149
tri 36502 38860 36791 39149 sw
tri 36791 38860 37080 39149 ne
rect 37080 39060 38678 39149
tri 38678 39060 38860 39242 sw
tri 38968 39060 39150 39242 ne
rect 39150 39238 42922 39242
tri 42922 39238 43216 39532 sw
tri 43216 39238 43510 39532 ne
rect 43510 39352 47352 39532
tri 47352 39352 47640 39640 sw
tri 47640 39352 47928 39640 ne
rect 47928 39456 51771 39640
tri 51771 39456 52068 39753 sw
tri 52068 39456 52365 39753 ne
rect 52365 39600 56172 39753
tri 56172 39600 56465 39893 sw
tri 56465 39600 56758 39893 ne
rect 56758 39600 71000 39893
rect 52365 39456 56465 39600
rect 47928 39352 52068 39456
rect 43510 39238 47640 39352
rect 39150 39076 43216 39238
tri 43216 39076 43378 39238 sw
tri 43510 39076 43672 39238 ne
rect 43672 39076 47640 39238
rect 39150 39060 43378 39076
rect 37080 38860 38860 39060
rect 30428 38702 34514 38860
rect 26184 38420 30146 38702
tri 30146 38420 30428 38702 sw
tri 30428 38420 30710 38702 ne
rect 30710 38563 34514 38702
tri 34514 38563 34811 38860 sw
tri 34811 38563 35108 38860 ne
rect 35108 38769 36791 38860
tri 36791 38769 36882 38860 sw
tri 37080 38769 37171 38860 ne
rect 37171 38770 38860 38860
tri 38860 38770 39150 39060 sw
tri 39150 38770 39440 39060 ne
rect 39440 38782 43378 39060
tri 43378 38782 43672 39076 sw
tri 43672 38782 43966 39076 ne
rect 43966 39064 47640 39076
tri 47640 39064 47928 39352 sw
tri 47928 39064 48216 39352 ne
rect 48216 39159 52068 39352
tri 52068 39159 52365 39456 sw
tri 52365 39159 52662 39456 ne
rect 52662 39400 56465 39456
tri 56465 39400 56665 39600 sw
rect 52662 39332 71000 39400
rect 52662 39159 70613 39332
rect 48216 39064 52365 39159
rect 43966 38782 47928 39064
rect 39440 38770 43672 38782
rect 37171 38769 39150 38770
rect 35108 38563 36882 38769
rect 30710 38420 34811 38563
tri 21648 34176 25892 38420 ne
tri 25892 38128 26184 38420 sw
tri 26184 38128 26476 38420 ne
rect 26476 38138 30428 38420
tri 30428 38138 30710 38420 sw
tri 30710 38138 30992 38420 ne
rect 30992 38266 34811 38420
tri 34811 38266 35108 38563 sw
tri 35108 38266 35405 38563 ne
rect 35405 38480 36882 38563
tri 36882 38480 37171 38769 sw
tri 37171 38480 37460 38769 ne
rect 37460 38480 39150 38769
tri 39150 38480 39440 38770 sw
tri 39440 38480 39730 38770 ne
rect 39730 38488 43672 38770
tri 43672 38488 43966 38782 sw
tri 43966 38488 44260 38782 ne
rect 44260 38776 47928 38782
tri 47928 38776 48216 39064 sw
tri 48216 38776 48504 39064 ne
rect 48504 38929 52365 39064
tri 52365 38929 52595 39159 sw
tri 52662 38929 52892 39159 ne
rect 52892 38929 70613 39159
rect 48504 38776 52595 38929
rect 44260 38488 48216 38776
tri 48216 38488 48504 38776 sw
tri 48504 38488 48792 38776 ne
rect 48792 38632 52595 38776
tri 52595 38632 52892 38929 sw
tri 52892 38632 53189 38929 ne
rect 53189 38632 70613 38929
rect 48792 38488 52892 38632
rect 39730 38480 43966 38488
rect 35405 38266 37171 38480
rect 30992 38138 35108 38266
rect 26476 38128 30710 38138
rect 25892 37836 26184 38128
tri 26184 37836 26476 38128 sw
tri 26476 37836 26768 38128 ne
rect 26768 37940 30710 38128
tri 30710 37940 30908 38138 sw
tri 30992 37940 31190 38138 ne
rect 31190 37969 35108 38138
tri 35108 37969 35405 38266 sw
tri 35405 37969 35702 38266 ne
rect 35702 38191 37171 38266
tri 37171 38191 37460 38480 sw
tri 37460 38191 37749 38480 ne
rect 37749 38191 39440 38480
rect 35702 37969 37460 38191
rect 31190 37940 35405 37969
rect 26768 37836 30908 37940
rect 25892 37544 26476 37836
tri 26476 37544 26768 37836 sw
tri 26768 37544 27060 37836 ne
rect 27060 37658 30908 37836
tri 30908 37658 31190 37940 sw
tri 31190 37658 31472 37940 ne
rect 31472 37771 35405 37940
tri 35405 37771 35603 37969 sw
tri 35702 37771 35900 37969 ne
rect 35900 37902 37460 37969
tri 37460 37902 37749 38191 sw
tri 37749 37902 38038 38191 ne
rect 38038 38190 39440 38191
tri 39440 38190 39730 38480 sw
tri 39730 38190 40020 38480 ne
rect 40020 38194 43966 38480
tri 43966 38194 44260 38488 sw
tri 44260 38194 44554 38488 ne
rect 44554 38200 48504 38488
tri 48504 38200 48792 38488 sw
tri 48792 38200 49080 38488 ne
rect 49080 38335 52892 38488
tri 52892 38335 53189 38632 sw
tri 53189 38335 53486 38632 ne
rect 53486 38335 70613 38632
rect 49080 38200 53189 38335
rect 44554 38194 48792 38200
rect 40020 38190 44260 38194
rect 38038 37902 39730 38190
rect 35900 37771 37749 37902
rect 31472 37658 35603 37771
rect 27060 37544 31190 37658
rect 25892 37252 26768 37544
tri 26768 37252 27060 37544 sw
tri 27060 37252 27352 37544 ne
rect 27352 37376 31190 37544
tri 31190 37376 31472 37658 sw
tri 31472 37376 31754 37658 ne
rect 31754 37474 35603 37658
tri 35603 37474 35900 37771 sw
tri 35900 37474 36197 37771 ne
rect 36197 37613 37749 37771
tri 37749 37613 38038 37902 sw
tri 38038 37613 38327 37902 ne
rect 38327 37900 39730 37902
tri 39730 37900 40020 38190 sw
tri 40020 37900 40310 38190 ne
rect 40310 37900 44260 38190
tri 44260 37900 44554 38194 sw
tri 44554 37900 44848 38194 ne
rect 44848 38020 48792 38194
tri 48792 38020 48972 38200 sw
tri 49080 38020 49260 38200 ne
rect 49260 38038 53189 38200
tri 53189 38038 53486 38335 sw
tri 53486 38038 53783 38335 ne
rect 53783 38038 70613 38335
rect 49260 38020 53486 38038
rect 44848 37900 48972 38020
rect 38327 37666 40020 37900
tri 40020 37666 40254 37900 sw
tri 40310 37666 40544 37900 ne
rect 40544 37666 44554 37900
rect 38327 37613 40254 37666
rect 36197 37474 38038 37613
rect 31754 37376 35900 37474
rect 27352 37252 31472 37376
rect 25892 36960 27060 37252
tri 27060 36960 27352 37252 sw
tri 27352 36960 27644 37252 ne
rect 27644 37094 31472 37252
tri 31472 37094 31754 37376 sw
tri 31754 37094 32036 37376 ne
rect 32036 37177 35900 37376
tri 35900 37177 36197 37474 sw
tri 36197 37177 36494 37474 ne
rect 36494 37458 38038 37474
tri 38038 37458 38193 37613 sw
tri 38327 37458 38482 37613 ne
rect 38482 37458 40254 37613
rect 36494 37177 38193 37458
rect 32036 37094 36197 37177
rect 27644 36960 31754 37094
rect 25892 36680 27352 36960
tri 27352 36680 27632 36960 sw
tri 27644 36680 27924 36960 ne
rect 27924 36812 31754 36960
tri 31754 36812 32036 37094 sw
tri 32036 36812 32318 37094 ne
rect 32318 36880 36197 37094
tri 36197 36880 36494 37177 sw
tri 36494 36880 36791 37177 ne
rect 36791 37169 38193 37177
tri 38193 37169 38482 37458 sw
tri 38482 37169 38771 37458 ne
rect 38771 37376 40254 37458
tri 40254 37376 40544 37666 sw
tri 40544 37376 40834 37666 ne
rect 40834 37606 44554 37666
tri 44554 37606 44848 37900 sw
tri 44848 37606 45142 37900 ne
rect 45142 37732 48972 37900
tri 48972 37732 49260 38020 sw
tri 49260 37732 49548 38020 ne
rect 49548 37741 53486 38020
tri 53486 37741 53783 38038 sw
tri 53783 37741 54080 38038 ne
rect 54080 37741 70613 38038
rect 49548 37732 53783 37741
rect 45142 37606 49260 37732
rect 40834 37376 44848 37606
rect 38771 37169 40544 37376
rect 36791 36880 38482 37169
tri 38482 36880 38771 37169 sw
tri 38771 36880 39060 37169 ne
rect 39060 37086 40544 37169
tri 40544 37086 40834 37376 sw
tri 40834 37086 41124 37376 ne
rect 41124 37312 44848 37376
tri 44848 37312 45142 37606 sw
tri 45142 37312 45436 37606 ne
rect 45436 37444 49260 37606
tri 49260 37444 49548 37732 sw
tri 49548 37444 49836 37732 ne
rect 49836 37444 53783 37732
tri 53783 37444 54080 37741 sw
tri 54080 37444 54377 37741 ne
rect 54377 37444 70613 37741
rect 45436 37312 49548 37444
rect 41124 37086 45142 37312
rect 39060 36880 40834 37086
tri 40834 36880 41040 37086 sw
tri 41124 36880 41330 37086 ne
rect 41330 37018 45142 37086
tri 45142 37018 45436 37312 sw
tri 45436 37018 45730 37312 ne
rect 45730 37156 49548 37312
tri 49548 37156 49836 37444 sw
tri 49836 37156 50124 37444 ne
rect 50124 37156 54080 37444
rect 45730 37018 49836 37156
rect 41330 36880 45436 37018
rect 32318 36812 36494 36880
rect 27924 36680 32036 36812
rect 25892 36388 27632 36680
tri 27632 36388 27924 36680 sw
tri 27924 36388 28216 36680 ne
rect 28216 36530 32036 36680
tri 32036 36530 32318 36812 sw
tri 32318 36530 32600 36812 ne
rect 32600 36583 36494 36812
tri 36494 36583 36791 36880 sw
tri 36791 36583 37088 36880 ne
rect 37088 36789 38771 36880
tri 38771 36789 38862 36880 sw
tri 39060 36789 39151 36880 ne
rect 39151 36790 41040 36880
tri 41040 36790 41130 36880 sw
tri 41330 36790 41420 36880 ne
rect 41420 36790 45436 36880
rect 39151 36789 41130 36790
rect 37088 36583 38862 36789
rect 32600 36530 36791 36583
rect 28216 36388 32318 36530
rect 25892 36096 27924 36388
tri 27924 36096 28216 36388 sw
tri 28216 36096 28508 36388 ne
rect 28508 36248 32318 36388
tri 32318 36248 32600 36530 sw
tri 32600 36248 32882 36530 ne
rect 32882 36286 36791 36530
tri 36791 36286 37088 36583 sw
tri 37088 36286 37385 36583 ne
rect 37385 36500 38862 36583
tri 38862 36500 39151 36789 sw
tri 39151 36500 39440 36789 ne
rect 39440 36500 41130 36789
tri 41130 36500 41420 36790 sw
tri 41420 36500 41710 36790 ne
rect 41710 36758 45436 36790
tri 45436 36758 45696 37018 sw
tri 45730 36758 45990 37018 ne
rect 45990 36868 49836 37018
tri 49836 36868 50124 37156 sw
tri 50124 36868 50412 37156 ne
rect 50412 37147 54080 37156
tri 54080 37147 54377 37444 sw
tri 54377 37147 54674 37444 ne
rect 54674 37147 70613 37444
rect 50412 36994 54377 37147
tri 54377 36994 54530 37147 sw
tri 54674 36994 54827 37147 ne
rect 54827 36994 70613 37147
rect 50412 36868 54530 36994
rect 45990 36758 50124 36868
rect 41710 36500 45696 36758
rect 37385 36286 39151 36500
rect 32882 36248 37088 36286
rect 28508 36096 32600 36248
rect 25892 35804 28216 36096
tri 28216 35804 28508 36096 sw
tri 28508 35804 28800 36096 ne
rect 28800 35966 32600 36096
tri 32600 35966 32882 36248 sw
tri 32882 35966 33164 36248 ne
rect 33164 35989 37088 36248
tri 37088 35989 37385 36286 sw
tri 37385 35989 37682 36286 ne
rect 37682 36211 39151 36286
tri 39151 36211 39440 36500 sw
tri 39440 36211 39729 36500 ne
rect 39729 36211 41420 36500
rect 37682 35989 39440 36211
rect 33164 35966 37385 35989
rect 28800 35804 32882 35966
rect 25892 35512 28508 35804
tri 28508 35512 28800 35804 sw
tri 28800 35512 29092 35804 ne
rect 29092 35684 32882 35804
tri 32882 35684 33164 35966 sw
tri 33164 35684 33446 35966 ne
rect 33446 35791 37385 35966
tri 37385 35791 37583 35989 sw
tri 37682 35791 37880 35989 ne
rect 37880 35922 39440 35989
tri 39440 35922 39729 36211 sw
tri 39729 35922 40018 36211 ne
rect 40018 36210 41420 36211
tri 41420 36210 41710 36500 sw
tri 41710 36210 42000 36500 ne
rect 42000 36464 45696 36500
tri 45696 36464 45990 36758 sw
tri 45990 36464 46284 36758 ne
rect 46284 36580 50124 36758
tri 50124 36580 50412 36868 sw
tri 50412 36580 50700 36868 ne
rect 50700 36697 54530 36868
tri 54530 36697 54827 36994 sw
tri 54827 36697 55124 36994 ne
rect 55124 36697 70613 36994
rect 50700 36580 54827 36697
rect 46284 36464 50412 36580
rect 42000 36210 45990 36464
rect 40018 35922 41710 36210
rect 37880 35791 39729 35922
rect 33446 35684 37583 35791
rect 29092 35586 33164 35684
tri 33164 35586 33262 35684 sw
tri 33446 35586 33544 35684 ne
rect 33544 35586 37583 35684
rect 29092 35512 33262 35586
rect 25892 35220 28800 35512
tri 28800 35220 29092 35512 sw
tri 29092 35220 29384 35512 ne
rect 29384 35304 33262 35512
tri 33262 35304 33544 35586 sw
tri 33544 35304 33826 35586 ne
rect 33826 35494 37583 35586
tri 37583 35494 37880 35791 sw
tri 37880 35494 38177 35791 ne
rect 38177 35633 39729 35791
tri 39729 35633 40018 35922 sw
tri 40018 35633 40307 35922 ne
rect 40307 35920 41710 35922
tri 41710 35920 42000 36210 sw
tri 42000 35920 42290 36210 ne
rect 42290 36170 45990 36210
tri 45990 36170 46284 36464 sw
tri 46284 36170 46578 36464 ne
rect 46578 36292 50412 36464
tri 50412 36292 50700 36580 sw
tri 50700 36292 50988 36580 ne
rect 50988 36400 54827 36580
tri 54827 36400 55124 36697 sw
tri 55124 36400 55421 36697 ne
rect 55421 36468 70613 36697
rect 70669 36468 71000 39332
rect 55421 36400 71000 36468
rect 50988 36292 55124 36400
rect 46578 36170 50700 36292
rect 42290 35920 46284 36170
rect 40307 35868 42000 35920
tri 42000 35868 42052 35920 sw
tri 42290 35868 42342 35920 ne
rect 42342 35876 46284 35920
tri 46284 35876 46578 36170 sw
tri 46578 35876 46872 36170 ne
rect 46872 36004 50700 36170
tri 50700 36004 50988 36292 sw
tri 50988 36004 51276 36292 ne
rect 51276 36200 55124 36292
tri 55124 36200 55324 36400 sw
rect 51276 36132 71000 36200
rect 51276 36004 70613 36132
rect 46872 35876 50988 36004
rect 42342 35868 46578 35876
rect 40307 35633 42052 35868
rect 38177 35494 40018 35633
rect 33826 35304 37880 35494
rect 29384 35220 33544 35304
rect 25892 34928 29092 35220
tri 29092 34928 29384 35220 sw
tri 29384 34928 29676 35220 ne
rect 29676 35022 33544 35220
tri 33544 35022 33826 35304 sw
tri 33826 35022 34108 35304 ne
rect 34108 35197 37880 35304
tri 37880 35197 38177 35494 sw
tri 38177 35197 38474 35494 ne
rect 38474 35478 40018 35494
tri 40018 35478 40173 35633 sw
tri 40307 35478 40462 35633 ne
rect 40462 35578 42052 35633
tri 42052 35578 42342 35868 sw
tri 42342 35578 42632 35868 ne
rect 42632 35582 46578 35868
tri 46578 35582 46872 35876 sw
tri 46872 35582 47166 35876 ne
rect 47166 35716 50988 35876
tri 50988 35716 51276 36004 sw
tri 51276 35716 51564 36004 ne
rect 51564 35716 70613 36004
rect 47166 35684 51276 35716
tri 51276 35684 51308 35716 sw
tri 51564 35684 51596 35716 ne
rect 51596 35684 70613 35716
rect 47166 35582 51308 35684
rect 42632 35578 46872 35582
rect 40462 35478 42342 35578
rect 38474 35197 40173 35478
rect 34108 35022 38177 35197
rect 29676 34928 33826 35022
rect 25892 34760 29384 34928
tri 29384 34760 29552 34928 sw
tri 29676 34760 29844 34928 ne
rect 29844 34760 33826 34928
rect 25892 34468 29552 34760
tri 29552 34468 29844 34760 sw
tri 29844 34468 30136 34760 ne
rect 30136 34740 33826 34760
tri 33826 34740 34108 35022 sw
tri 34108 34740 34390 35022 ne
rect 34390 34900 38177 35022
tri 38177 34900 38474 35197 sw
tri 38474 34900 38771 35197 ne
rect 38771 35189 40173 35197
tri 40173 35189 40462 35478 sw
tri 40462 35189 40751 35478 ne
rect 40751 35288 42342 35478
tri 42342 35288 42632 35578 sw
tri 42632 35288 42922 35578 ne
rect 42922 35288 46872 35578
tri 46872 35288 47166 35582 sw
tri 47166 35288 47460 35582 ne
rect 47460 35396 51308 35582
tri 51308 35396 51596 35684 sw
tri 51596 35396 51884 35684 ne
rect 51884 35396 70613 35684
rect 47460 35288 51596 35396
rect 40751 35189 42632 35288
rect 38771 34900 40462 35189
tri 40462 34900 40751 35189 sw
tri 40751 34900 41040 35189 ne
rect 41040 34998 42632 35189
tri 42632 34998 42922 35288 sw
tri 42922 34998 43212 35288 ne
rect 43212 34998 47166 35288
rect 41040 34900 42922 34998
rect 34390 34740 38474 34900
rect 30136 34468 34108 34740
rect 25892 34176 29844 34468
tri 29844 34176 30136 34468 sw
tri 30136 34176 30428 34468 ne
rect 30428 34458 34108 34468
tri 34108 34458 34390 34740 sw
tri 34390 34458 34672 34740 ne
rect 34672 34603 38474 34740
tri 38474 34603 38771 34900 sw
tri 38771 34603 39068 34900 ne
rect 39068 34809 40751 34900
tri 40751 34809 40842 34900 sw
tri 41040 34809 41131 34900 ne
rect 41131 34810 42922 34900
tri 42922 34810 43110 34998 sw
tri 43212 34810 43400 34998 ne
rect 43400 34994 47166 34998
tri 47166 34994 47460 35288 sw
tri 47460 34994 47754 35288 ne
rect 47754 35108 51596 35288
tri 51596 35108 51884 35396 sw
tri 51884 35108 52172 35396 ne
rect 52172 35108 70613 35396
rect 47754 34994 51884 35108
rect 43400 34832 47460 34994
tri 47460 34832 47622 34994 sw
tri 47754 34832 47916 34994 ne
rect 47916 34832 51884 34994
rect 43400 34810 47622 34832
rect 41131 34809 43110 34810
rect 39068 34603 40842 34809
rect 34672 34458 38771 34603
rect 30428 34176 34390 34458
tri 34390 34176 34672 34458 sw
tri 34672 34176 34954 34458 ne
rect 34954 34306 38771 34458
tri 38771 34306 39068 34603 sw
tri 39068 34306 39365 34603 ne
rect 39365 34520 40842 34603
tri 40842 34520 41131 34809 sw
tri 41131 34520 41420 34809 ne
rect 41420 34520 43110 34809
tri 43110 34520 43400 34810 sw
tri 43400 34520 43690 34810 ne
rect 43690 34538 47622 34810
tri 47622 34538 47916 34832 sw
tri 47916 34538 48210 34832 ne
rect 48210 34820 51884 34832
tri 51884 34820 52172 35108 sw
tri 52172 34820 52460 35108 ne
rect 52460 34820 70613 35108
rect 48210 34538 52172 34820
rect 43690 34520 47916 34538
rect 39365 34306 41131 34520
rect 34954 34176 39068 34306
tri 25892 29932 30136 34176 ne
tri 30136 33884 30428 34176 sw
tri 30428 33884 30720 34176 ne
rect 30720 33894 34672 34176
tri 34672 33894 34954 34176 sw
tri 34954 33894 35236 34176 ne
rect 35236 34009 39068 34176
tri 39068 34009 39365 34306 sw
tri 39365 34009 39662 34306 ne
rect 39662 34231 41131 34306
tri 41131 34231 41420 34520 sw
tri 41420 34231 41709 34520 ne
rect 41709 34244 43400 34520
tri 43400 34244 43676 34520 sw
tri 43690 34244 43966 34520 ne
rect 43966 34244 47916 34520
tri 47916 34244 48210 34538 sw
tri 48210 34244 48504 34538 ne
rect 48504 34532 52172 34538
tri 52172 34532 52460 34820 sw
tri 52460 34532 52748 34820 ne
rect 52748 34532 70613 34820
rect 48504 34244 52460 34532
tri 52460 34244 52748 34532 sw
tri 52748 34244 53036 34532 ne
rect 53036 34244 70613 34532
rect 41709 34231 43676 34244
rect 39662 34009 41420 34231
rect 35236 33894 39365 34009
rect 30720 33884 34954 33894
rect 30136 33592 30428 33884
tri 30428 33592 30720 33884 sw
tri 30720 33592 31012 33884 ne
rect 31012 33696 34954 33884
tri 34954 33696 35152 33894 sw
tri 35236 33696 35434 33894 ne
rect 35434 33811 39365 33894
tri 39365 33811 39563 34009 sw
tri 39662 33811 39860 34009 ne
rect 39860 33942 41420 34009
tri 41420 33942 41709 34231 sw
tri 41709 33942 41998 34231 ne
rect 41998 33954 43676 34231
tri 43676 33954 43966 34244 sw
tri 43966 33954 44256 34244 ne
rect 44256 33954 48210 34244
rect 41998 33942 43966 33954
rect 39860 33811 41709 33942
rect 35434 33696 39563 33811
rect 31012 33592 35152 33696
rect 30136 33300 30720 33592
tri 30720 33300 31012 33592 sw
tri 31012 33300 31304 33592 ne
rect 31304 33414 35152 33592
tri 35152 33414 35434 33696 sw
tri 35434 33414 35716 33696 ne
rect 35716 33514 39563 33696
tri 39563 33514 39860 33811 sw
tri 39860 33514 40157 33811 ne
rect 40157 33653 41709 33811
tri 41709 33653 41998 33942 sw
tri 41998 33653 42287 33942 ne
rect 42287 33664 43966 33942
tri 43966 33664 44256 33954 sw
tri 44256 33664 44546 33954 ne
rect 44546 33950 48210 33954
tri 48210 33950 48504 34244 sw
tri 48504 33950 48798 34244 ne
rect 48798 33956 52748 34244
tri 52748 33956 53036 34244 sw
tri 53036 33956 53324 34244 ne
rect 53324 33956 70613 34244
rect 48798 33950 53036 33956
rect 44546 33664 48504 33950
rect 42287 33653 44256 33664
rect 40157 33514 41998 33653
rect 35716 33414 39860 33514
rect 31304 33300 35434 33414
rect 30136 33008 31012 33300
tri 31012 33008 31304 33300 sw
tri 31304 33008 31596 33300 ne
rect 31596 33132 35434 33300
tri 35434 33132 35716 33414 sw
tri 35716 33132 35998 33414 ne
rect 35998 33217 39860 33414
tri 39860 33217 40157 33514 sw
tri 40157 33217 40454 33514 ne
rect 40454 33498 41998 33514
tri 41998 33498 42153 33653 sw
tri 42287 33498 42442 33653 ne
rect 42442 33498 44256 33653
rect 40454 33217 42153 33498
rect 35998 33132 40157 33217
rect 31596 33008 35716 33132
rect 30136 32716 31304 33008
tri 31304 32716 31596 33008 sw
tri 31596 32716 31888 33008 ne
rect 31888 32850 35716 33008
tri 35716 32850 35998 33132 sw
tri 35998 32850 36280 33132 ne
rect 36280 32920 40157 33132
tri 40157 32920 40454 33217 sw
tri 40454 32920 40751 33217 ne
rect 40751 33209 42153 33217
tri 42153 33209 42442 33498 sw
tri 42442 33209 42731 33498 ne
rect 42731 33422 44256 33498
tri 44256 33422 44498 33664 sw
tri 44546 33422 44788 33664 ne
rect 44788 33656 48504 33664
tri 48504 33656 48798 33950 sw
tri 48798 33656 49092 33950 ne
rect 49092 33776 53036 33950
tri 53036 33776 53216 33956 sw
tri 53324 33776 53504 33956 ne
rect 53504 33776 70613 33956
rect 49092 33656 53216 33776
rect 44788 33422 48798 33656
rect 42731 33209 44498 33422
rect 40751 32920 42442 33209
tri 42442 32920 42731 33209 sw
tri 42731 32920 43020 33209 ne
rect 43020 33132 44498 33209
tri 44498 33132 44788 33422 sw
tri 44788 33132 45078 33422 ne
rect 45078 33362 48798 33422
tri 48798 33362 49092 33656 sw
tri 49092 33362 49386 33656 ne
rect 49386 33488 53216 33656
tri 53216 33488 53504 33776 sw
tri 53504 33488 53792 33776 ne
rect 53792 33488 70613 33776
rect 49386 33362 53504 33488
rect 45078 33132 49092 33362
rect 43020 32920 44788 33132
rect 36280 32850 40454 32920
rect 31888 32716 35998 32850
rect 30136 32436 31596 32716
tri 31596 32436 31876 32716 sw
tri 31888 32436 32168 32716 ne
rect 32168 32568 35998 32716
tri 35998 32568 36280 32850 sw
tri 36280 32568 36562 32850 ne
rect 36562 32623 40454 32850
tri 40454 32623 40751 32920 sw
tri 40751 32623 41048 32920 ne
rect 41048 32829 42731 32920
tri 42731 32829 42822 32920 sw
tri 43020 32829 43111 32920 ne
rect 43111 32842 44788 32920
tri 44788 32842 45078 33132 sw
tri 45078 32842 45368 33132 ne
rect 45368 33068 49092 33132
tri 49092 33068 49386 33362 sw
tri 49386 33068 49680 33362 ne
rect 49680 33200 53504 33362
tri 53504 33200 53792 33488 sw
tri 53792 33200 54080 33488 ne
rect 54080 33268 70613 33488
rect 70669 33268 71000 36132
rect 54080 33200 71000 33268
rect 49680 33068 53792 33200
rect 45368 32842 49386 33068
rect 43111 32830 45078 32842
tri 45078 32830 45090 32842 sw
tri 45368 32830 45380 32842 ne
rect 45380 32830 49386 32842
rect 43111 32829 45090 32830
rect 41048 32623 42822 32829
rect 36562 32568 40751 32623
rect 32168 32436 36280 32568
rect 30136 32144 31876 32436
tri 31876 32144 32168 32436 sw
tri 32168 32144 32460 32436 ne
rect 32460 32286 36280 32436
tri 36280 32286 36562 32568 sw
tri 36562 32286 36844 32568 ne
rect 36844 32326 40751 32568
tri 40751 32326 41048 32623 sw
tri 41048 32326 41345 32623 ne
rect 41345 32540 42822 32623
tri 42822 32540 43111 32829 sw
tri 43111 32540 43400 32829 ne
rect 43400 32540 45090 32829
tri 45090 32540 45380 32830 sw
tri 45380 32540 45670 32830 ne
rect 45670 32774 49386 32830
tri 49386 32774 49680 33068 sw
tri 49680 32774 49974 33068 ne
rect 49974 33000 53792 33068
tri 53792 33000 53992 33200 sw
rect 49974 32920 71000 33000
rect 49974 32774 70613 32920
rect 45670 32540 49680 32774
rect 41345 32326 43111 32540
rect 36844 32286 41048 32326
rect 32460 32144 36562 32286
rect 30136 31852 32168 32144
tri 32168 31852 32460 32144 sw
tri 32460 31852 32752 32144 ne
rect 32752 32004 36562 32144
tri 36562 32004 36844 32286 sw
tri 36844 32004 37126 32286 ne
rect 37126 32029 41048 32286
tri 41048 32029 41345 32326 sw
tri 41345 32029 41642 32326 ne
rect 41642 32251 43111 32326
tri 43111 32251 43400 32540 sw
tri 43400 32251 43689 32540 ne
rect 43689 32251 45380 32540
rect 41642 32029 43400 32251
rect 37126 32004 41345 32029
rect 32752 31852 36844 32004
rect 30136 31560 32460 31852
tri 32460 31560 32752 31852 sw
tri 32752 31560 33044 31852 ne
rect 33044 31722 36844 31852
tri 36844 31722 37126 32004 sw
tri 37126 31722 37408 32004 ne
rect 37408 31831 41345 32004
tri 41345 31831 41543 32029 sw
tri 41642 31831 41840 32029 ne
rect 41840 31962 43400 32029
tri 43400 31962 43689 32251 sw
tri 43689 31962 43978 32251 ne
rect 43978 32250 45380 32251
tri 45380 32250 45670 32540 sw
tri 45670 32250 45960 32540 ne
rect 45960 32514 49680 32540
tri 49680 32514 49940 32774 sw
tri 49974 32514 50234 32774 ne
rect 50234 32514 70613 32774
rect 45960 32250 49940 32514
rect 43978 31962 45670 32250
rect 41840 31831 43689 31962
rect 37408 31722 41543 31831
rect 33044 31560 37126 31722
rect 30136 31268 32752 31560
tri 32752 31268 33044 31560 sw
tri 33044 31268 33336 31560 ne
rect 33336 31440 37126 31560
tri 37126 31440 37408 31722 sw
tri 37408 31440 37690 31722 ne
rect 37690 31534 41543 31722
tri 41543 31534 41840 31831 sw
tri 41840 31534 42137 31831 ne
rect 42137 31673 43689 31831
tri 43689 31673 43978 31962 sw
tri 43978 31673 44267 31962 ne
rect 44267 31960 45670 31962
tri 45670 31960 45960 32250 sw
tri 45960 31960 46250 32250 ne
rect 46250 32220 49940 32250
tri 49940 32220 50234 32514 sw
tri 50234 32220 50528 32514 ne
rect 50528 32220 70613 32514
rect 46250 31960 50234 32220
rect 44267 31673 45960 31960
rect 42137 31534 43978 31673
rect 37690 31440 41840 31534
rect 33336 31342 37408 31440
tri 37408 31342 37506 31440 sw
tri 37690 31342 37788 31440 ne
rect 37788 31342 41840 31440
rect 33336 31268 37506 31342
rect 30136 30976 33044 31268
tri 33044 30976 33336 31268 sw
tri 33336 30976 33628 31268 ne
rect 33628 31060 37506 31268
tri 37506 31060 37788 31342 sw
tri 37788 31060 38070 31342 ne
rect 38070 31237 41840 31342
tri 41840 31237 42137 31534 sw
tri 42137 31237 42434 31534 ne
rect 42434 31518 43978 31534
tri 43978 31518 44133 31673 sw
tri 44267 31518 44422 31673 ne
rect 44422 31670 45960 31673
tri 45960 31670 46250 31960 sw
tri 46250 31670 46540 31960 ne
rect 46540 31926 50234 31960
tri 50234 31926 50528 32220 sw
tri 50528 31926 50822 32220 ne
rect 50822 31926 70613 32220
rect 46540 31670 50528 31926
rect 44422 31624 46250 31670
tri 46250 31624 46296 31670 sw
tri 46540 31624 46586 31670 ne
rect 46586 31632 50528 31670
tri 50528 31632 50822 31926 sw
tri 50822 31632 51116 31926 ne
rect 51116 31632 70613 31926
rect 46586 31624 50822 31632
rect 44422 31518 46296 31624
rect 42434 31237 44133 31518
rect 38070 31060 42137 31237
rect 33628 30976 37788 31060
rect 30136 30684 33336 30976
tri 33336 30684 33628 30976 sw
tri 33628 30684 33920 30976 ne
rect 33920 30778 37788 30976
tri 37788 30778 38070 31060 sw
tri 38070 30778 38352 31060 ne
rect 38352 30940 42137 31060
tri 42137 30940 42434 31237 sw
tri 42434 30940 42731 31237 ne
rect 42731 31229 44133 31237
tri 44133 31229 44422 31518 sw
tri 44422 31229 44711 31518 ne
rect 44711 31334 46296 31518
tri 46296 31334 46586 31624 sw
tri 46586 31334 46876 31624 ne
rect 46876 31338 50822 31624
tri 50822 31338 51116 31632 sw
tri 51116 31338 51410 31632 ne
rect 51410 31338 70613 31632
rect 46876 31334 51116 31338
rect 44711 31229 46586 31334
rect 42731 30940 44422 31229
tri 44422 30940 44711 31229 sw
tri 44711 30940 45000 31229 ne
rect 45000 31044 46586 31229
tri 46586 31044 46876 31334 sw
tri 46876 31044 47166 31334 ne
rect 47166 31044 51116 31334
tri 51116 31044 51410 31338 sw
tri 51410 31044 51704 31338 ne
rect 51704 31044 70613 31338
rect 45000 30940 46876 31044
rect 38352 30778 42434 30940
rect 33920 30684 38070 30778
rect 30136 30516 33628 30684
tri 33628 30516 33796 30684 sw
tri 33920 30516 34088 30684 ne
rect 34088 30516 38070 30684
rect 30136 30224 33796 30516
tri 33796 30224 34088 30516 sw
tri 34088 30224 34380 30516 ne
rect 34380 30496 38070 30516
tri 38070 30496 38352 30778 sw
tri 38352 30496 38634 30778 ne
rect 38634 30643 42434 30778
tri 42434 30643 42731 30940 sw
tri 42731 30643 43028 30940 ne
rect 43028 30849 44711 30940
tri 44711 30849 44802 30940 sw
tri 45000 30849 45091 30940 ne
rect 45091 30850 46876 30940
tri 46876 30850 47070 31044 sw
tri 47166 30850 47360 31044 ne
rect 47360 30850 51410 31044
rect 45091 30849 47070 30850
rect 43028 30643 44802 30849
rect 38634 30496 42731 30643
rect 34380 30224 38352 30496
rect 30136 29932 34088 30224
tri 34088 29932 34380 30224 sw
tri 34380 29932 34672 30224 ne
rect 34672 30214 38352 30224
tri 38352 30214 38634 30496 sw
tri 38634 30214 38916 30496 ne
rect 38916 30346 42731 30496
tri 42731 30346 43028 30643 sw
tri 43028 30346 43325 30643 ne
rect 43325 30560 44802 30643
tri 44802 30560 45091 30849 sw
tri 45091 30560 45380 30849 ne
rect 45380 30560 47070 30849
tri 47070 30560 47360 30850 sw
tri 47360 30560 47650 30850 ne
rect 47650 30750 51410 30850
tri 51410 30750 51704 31044 sw
tri 51704 30750 51998 31044 ne
rect 51998 30750 70613 31044
rect 47650 30588 51704 30750
tri 51704 30588 51866 30750 sw
tri 51998 30588 52160 30750 ne
rect 52160 30588 70613 30750
rect 47650 30560 51866 30588
rect 43325 30346 45091 30560
rect 38916 30214 43028 30346
rect 34672 29932 38634 30214
tri 38634 29932 38916 30214 sw
tri 38916 29932 39198 30214 ne
rect 39198 30049 43028 30214
tri 43028 30049 43325 30346 sw
tri 43325 30049 43622 30346 ne
rect 43622 30271 45091 30346
tri 45091 30271 45380 30560 sw
tri 45380 30271 45669 30560 ne
rect 45669 30271 47360 30560
rect 43622 30049 45380 30271
rect 39198 29932 43325 30049
tri 30136 25688 34380 29932 ne
tri 34380 29640 34672 29932 sw
tri 34672 29640 34964 29932 ne
rect 34964 29650 38916 29932
tri 38916 29650 39198 29932 sw
tri 39198 29650 39480 29932 ne
rect 39480 29752 43325 29932
tri 43325 29752 43622 30049 sw
tri 43622 29752 43919 30049 ne
rect 43919 29982 45380 30049
tri 45380 29982 45669 30271 sw
tri 45669 29982 45958 30271 ne
rect 45958 30270 47360 30271
tri 47360 30270 47650 30560 sw
tri 47650 30270 47940 30560 ne
rect 47940 30294 51866 30560
tri 51866 30294 52160 30588 sw
tri 52160 30294 52454 30588 ne
rect 52454 30294 70613 30588
rect 47940 30270 52160 30294
rect 45958 30000 47650 30270
tri 47650 30000 47920 30270 sw
tri 47940 30000 48210 30270 ne
rect 48210 30000 52160 30270
tri 52160 30000 52454 30294 sw
tri 52454 30000 52748 30294 ne
rect 52748 30056 70613 30294
rect 70669 30056 71000 32920
rect 52748 30000 71000 30056
rect 45958 29982 47920 30000
rect 43919 29752 45669 29982
rect 39480 29650 43622 29752
rect 34964 29640 39198 29650
rect 34380 29348 34672 29640
tri 34672 29348 34964 29640 sw
tri 34964 29348 35256 29640 ne
rect 35256 29452 39198 29640
tri 39198 29452 39396 29650 sw
tri 39480 29452 39678 29650 ne
rect 39678 29554 43622 29650
tri 43622 29554 43820 29752 sw
tri 43919 29554 44117 29752 ne
rect 44117 29693 45669 29752
tri 45669 29693 45958 29982 sw
tri 45958 29693 46247 29982 ne
rect 46247 29710 47920 29982
tri 47920 29710 48210 30000 sw
tri 48210 29710 48500 30000 ne
rect 48500 29800 52454 30000
tri 52454 29800 52654 30000 sw
rect 48500 29752 71000 29800
rect 48500 29710 70613 29752
rect 46247 29693 48210 29710
rect 44117 29554 45958 29693
rect 39678 29452 43820 29554
rect 35256 29348 39396 29452
rect 34380 29056 34964 29348
tri 34964 29056 35256 29348 sw
tri 35256 29056 35548 29348 ne
rect 35548 29170 39396 29348
tri 39396 29170 39678 29452 sw
tri 39678 29170 39960 29452 ne
rect 39960 29257 43820 29452
tri 43820 29257 44117 29554 sw
tri 44117 29257 44414 29554 ne
rect 44414 29466 45958 29554
tri 45958 29466 46185 29693 sw
tri 46247 29466 46474 29693 ne
rect 46474 29466 48210 29693
rect 44414 29257 46185 29466
rect 39960 29170 44117 29257
rect 35548 29056 39678 29170
rect 34380 28764 35256 29056
tri 35256 28764 35548 29056 sw
tri 35548 28764 35840 29056 ne
rect 35840 28888 39678 29056
tri 39678 28888 39960 29170 sw
tri 39960 28888 40242 29170 ne
rect 40242 28960 44117 29170
tri 44117 28960 44414 29257 sw
tri 44414 28960 44711 29257 ne
rect 44711 29177 46185 29257
tri 46185 29177 46474 29466 sw
tri 46474 29177 46763 29466 ne
rect 46763 29420 48210 29466
tri 48210 29420 48500 29710 sw
tri 48500 29420 48790 29710 ne
rect 48790 29420 70613 29710
rect 46763 29178 48500 29420
tri 48500 29178 48742 29420 sw
tri 48790 29178 49032 29420 ne
rect 49032 29178 70613 29420
rect 46763 29177 48742 29178
rect 44711 28960 46474 29177
rect 40242 28888 44414 28960
rect 35840 28764 39960 28888
rect 34380 28472 35548 28764
tri 35548 28472 35840 28764 sw
tri 35840 28472 36132 28764 ne
rect 36132 28606 39960 28764
tri 39960 28606 40242 28888 sw
tri 40242 28606 40524 28888 ne
rect 40524 28663 44414 28888
tri 44414 28663 44711 28960 sw
tri 44711 28663 45008 28960 ne
rect 45008 28888 46474 28960
tri 46474 28888 46763 29177 sw
tri 46763 28888 47052 29177 ne
rect 47052 28888 48742 29177
tri 48742 28888 49032 29178 sw
tri 49032 28888 49322 29178 ne
rect 49322 28888 70613 29178
rect 45008 28869 46763 28888
tri 46763 28869 46782 28888 sw
tri 47052 28869 47071 28888 ne
rect 47071 28870 49032 28888
tri 49032 28870 49050 28888 sw
tri 49322 28870 49340 28888 ne
rect 49340 28870 70613 28888
rect 47071 28869 49050 28870
rect 45008 28663 46782 28869
rect 40524 28606 44711 28663
rect 36132 28472 40242 28606
rect 34380 28192 35840 28472
tri 35840 28192 36120 28472 sw
tri 36132 28192 36412 28472 ne
rect 36412 28324 40242 28472
tri 40242 28324 40524 28606 sw
tri 40524 28324 40806 28606 ne
rect 40806 28366 44711 28606
tri 44711 28366 45008 28663 sw
tri 45008 28366 45305 28663 ne
rect 45305 28580 46782 28663
tri 46782 28580 47071 28869 sw
tri 47071 28580 47360 28869 ne
rect 47360 28580 49050 28869
tri 49050 28580 49340 28870 sw
tri 49340 28580 49630 28870 ne
rect 49630 28580 70613 28870
rect 45305 28366 47071 28580
rect 40806 28324 45008 28366
rect 36412 28192 40524 28324
rect 34380 27900 36120 28192
tri 36120 27900 36412 28192 sw
tri 36412 27900 36704 28192 ne
rect 36704 28042 40524 28192
tri 40524 28042 40806 28324 sw
tri 40806 28042 41088 28324 ne
rect 41088 28069 45008 28324
tri 45008 28069 45305 28366 sw
tri 45305 28069 45602 28366 ne
rect 45602 28291 47071 28366
tri 47071 28291 47360 28580 sw
tri 47360 28291 47649 28580 ne
rect 47649 28291 49340 28580
rect 45602 28069 47360 28291
rect 41088 28042 45305 28069
rect 36704 27900 40806 28042
rect 34380 27608 36412 27900
tri 36412 27608 36704 27900 sw
tri 36704 27608 36996 27900 ne
rect 36996 27760 40806 27900
tri 40806 27760 41088 28042 sw
tri 41088 27760 41370 28042 ne
rect 41370 27871 45305 28042
tri 45305 27871 45503 28069 sw
tri 45602 27871 45800 28069 ne
rect 45800 28002 47360 28069
tri 47360 28002 47649 28291 sw
tri 47649 28002 47938 28291 ne
rect 47938 28290 49340 28291
tri 49340 28290 49630 28580 sw
tri 49630 28290 49920 28580 ne
rect 49920 28290 70613 28580
rect 47938 28002 49630 28290
rect 45800 27871 47649 28002
rect 41370 27760 45503 27871
rect 36996 27608 41088 27760
rect 34380 27316 36704 27608
tri 36704 27316 36996 27608 sw
tri 36996 27316 37288 27608 ne
rect 37288 27478 41088 27608
tri 41088 27478 41370 27760 sw
tri 41370 27478 41652 27760 ne
rect 41652 27574 45503 27760
tri 45503 27574 45800 27871 sw
tri 45800 27574 46097 27871 ne
rect 46097 27713 47649 27871
tri 47649 27713 47938 28002 sw
tri 47938 27713 48227 28002 ne
rect 48227 28000 49630 28002
tri 49630 28000 49920 28290 sw
tri 49920 28000 50210 28290 ne
rect 50210 28000 70613 28290
rect 48227 27713 49920 28000
rect 46097 27667 47938 27713
tri 47938 27667 47984 27713 sw
tri 48227 27667 48273 27713 ne
rect 48273 27710 49920 27713
tri 49920 27710 50210 28000 sw
tri 50210 27710 50500 28000 ne
rect 50500 27710 70613 28000
rect 48273 27667 50210 27710
rect 46097 27574 47984 27667
rect 41652 27478 45800 27574
rect 37288 27316 41370 27478
rect 34380 27024 36996 27316
tri 36996 27024 37288 27316 sw
tri 37288 27024 37580 27316 ne
rect 37580 27196 41370 27316
tri 41370 27196 41652 27478 sw
tri 41652 27196 41934 27478 ne
rect 41934 27277 45800 27478
tri 45800 27277 46097 27574 sw
tri 46097 27277 46394 27574 ne
rect 46394 27378 47984 27574
tri 47984 27378 48273 27667 sw
tri 48273 27378 48562 27667 ne
rect 48562 27470 50210 27667
tri 50210 27470 50450 27710 sw
tri 50500 27470 50740 27710 ne
rect 50740 27470 70613 27710
rect 48562 27378 50450 27470
rect 46394 27277 48273 27378
rect 41934 27196 46097 27277
rect 37580 27098 41652 27196
tri 41652 27098 41750 27196 sw
tri 41934 27098 42032 27196 ne
rect 42032 27098 46097 27196
rect 37580 27024 41750 27098
rect 34380 26732 37288 27024
tri 37288 26732 37580 27024 sw
tri 37580 26732 37872 27024 ne
rect 37872 26816 41750 27024
tri 41750 26816 42032 27098 sw
tri 42032 26816 42314 27098 ne
rect 42314 26980 46097 27098
tri 46097 26980 46394 27277 sw
tri 46394 26980 46691 27277 ne
rect 46691 27089 48273 27277
tri 48273 27089 48562 27378 sw
tri 48562 27089 48851 27378 ne
rect 48851 27180 50450 27378
tri 50450 27180 50740 27470 sw
tri 50740 27180 51030 27470 ne
rect 51030 27180 70613 27470
rect 48851 27089 50740 27180
rect 46691 26980 48562 27089
rect 42314 26816 46394 26980
rect 37872 26732 42032 26816
rect 34380 26440 37580 26732
tri 37580 26440 37872 26732 sw
tri 37872 26440 38164 26732 ne
rect 38164 26534 42032 26732
tri 42032 26534 42314 26816 sw
tri 42314 26534 42596 26816 ne
rect 42596 26683 46394 26816
tri 46394 26683 46691 26980 sw
tri 46691 26683 46988 26980 ne
rect 46988 26800 48562 26980
tri 48562 26800 48851 27089 sw
tri 48851 26800 49140 27089 ne
rect 49140 26890 50740 27089
tri 50740 26890 51030 27180 sw
tri 51030 26890 51320 27180 ne
rect 51320 26890 70613 27180
rect 49140 26800 51030 26890
rect 46988 26683 48851 26800
rect 42596 26534 46691 26683
rect 38164 26440 42314 26534
rect 34380 26272 37872 26440
tri 37872 26272 38040 26440 sw
tri 38164 26272 38332 26440 ne
rect 38332 26272 42314 26440
rect 34380 25980 38040 26272
tri 38040 25980 38332 26272 sw
tri 38332 25980 38624 26272 ne
rect 38624 26252 42314 26272
tri 42314 26252 42596 26534 sw
tri 42596 26252 42878 26534 ne
rect 42878 26386 46691 26534
tri 46691 26386 46988 26683 sw
tri 46988 26386 47285 26683 ne
rect 47285 26600 48851 26683
tri 48851 26600 49051 26800 sw
tri 49140 26600 49340 26800 ne
rect 49340 26600 51030 26800
tri 51030 26600 51320 26890 sw
tri 51320 26800 51410 26890 ne
rect 51410 26888 70613 26890
rect 70669 26888 71000 29752
rect 51410 26800 71000 26888
rect 47285 26386 49051 26600
rect 42878 26252 46988 26386
rect 38624 25980 42596 26252
rect 34380 25688 38332 25980
tri 38332 25688 38624 25980 sw
tri 38624 25688 38916 25980 ne
rect 38916 25970 42596 25980
tri 42596 25970 42878 26252 sw
tri 42878 25970 43160 26252 ne
rect 43160 26089 46988 26252
tri 46988 26089 47285 26386 sw
tri 47285 26089 47582 26386 ne
rect 47582 26311 49051 26386
tri 49051 26311 49340 26600 sw
tri 49340 26311 49629 26600 ne
rect 49629 26311 71000 26600
rect 47582 26089 49340 26311
rect 43160 25970 47285 26089
rect 38916 25688 42878 25970
tri 42878 25688 43160 25970 sw
tri 43160 25688 43442 25970 ne
rect 43442 25891 47285 25970
tri 47285 25891 47483 26089 sw
tri 47582 25891 47780 26089 ne
rect 47780 26022 49340 26089
tri 49340 26022 49629 26311 sw
tri 49629 26022 49918 26311 ne
rect 49918 26022 71000 26311
rect 47780 25891 49629 26022
rect 43442 25688 47483 25891
tri 34380 21444 38624 25688 ne
tri 38624 25396 38916 25688 sw
tri 38916 25396 39208 25688 ne
rect 39208 25406 43160 25688
tri 43160 25406 43442 25688 sw
tri 43442 25406 43724 25688 ne
rect 43724 25594 47483 25688
tri 47483 25594 47780 25891 sw
tri 47780 25594 48077 25891 ne
rect 48077 25778 49629 25891
tri 49629 25778 49873 26022 sw
tri 49918 25778 50162 26022 ne
rect 50162 25778 71000 26022
rect 48077 25594 49873 25778
rect 43724 25406 47780 25594
rect 39208 25396 43442 25406
rect 38624 25104 38916 25396
tri 38916 25104 39208 25396 sw
tri 39208 25104 39500 25396 ne
rect 39500 25208 43442 25396
tri 43442 25208 43640 25406 sw
tri 43724 25208 43922 25406 ne
rect 43922 25297 47780 25406
tri 47780 25297 48077 25594 sw
tri 48077 25297 48374 25594 ne
rect 48374 25489 49873 25594
tri 49873 25489 50162 25778 sw
tri 50162 25489 50451 25778 ne
rect 50451 25489 71000 25778
rect 48374 25297 50162 25489
rect 43922 25208 48077 25297
rect 39500 25104 43640 25208
rect 38624 24812 39208 25104
tri 39208 24812 39500 25104 sw
tri 39500 24812 39792 25104 ne
rect 39792 24926 43640 25104
tri 43640 24926 43922 25208 sw
tri 43922 24926 44204 25208 ne
rect 44204 25000 48077 25208
tri 48077 25000 48374 25297 sw
tri 48374 25000 48671 25297 ne
rect 48671 25200 50162 25297
tri 50162 25200 50451 25489 sw
tri 50451 25200 50740 25489 ne
rect 50740 25200 71000 25489
rect 48671 25000 50451 25200
tri 50451 25000 50651 25200 sw
rect 44204 24926 48374 25000
rect 39792 24812 43922 24926
rect 38624 24520 39500 24812
tri 39500 24520 39792 24812 sw
tri 39792 24520 40084 24812 ne
rect 40084 24644 43922 24812
tri 43922 24644 44204 24926 sw
tri 44204 24644 44486 24926 ne
rect 44486 24703 48374 24926
tri 48374 24703 48671 25000 sw
tri 48671 24703 48968 25000 ne
rect 48968 24906 71000 25000
rect 48968 24703 70613 24906
rect 44486 24644 48671 24703
rect 40084 24520 44204 24644
rect 38624 24228 39792 24520
tri 39792 24228 40084 24520 sw
tri 40084 24228 40376 24520 ne
rect 40376 24362 44204 24520
tri 44204 24362 44486 24644 sw
tri 44486 24362 44768 24644 ne
rect 44768 24406 48671 24644
tri 48671 24406 48968 24703 sw
tri 48968 24406 49265 24703 ne
rect 49265 24406 70613 24703
rect 44768 24362 48968 24406
rect 40376 24228 44486 24362
rect 38624 23948 40084 24228
tri 40084 23948 40364 24228 sw
tri 40376 23948 40656 24228 ne
rect 40656 24080 44486 24228
tri 44486 24080 44768 24362 sw
tri 44768 24080 45050 24362 ne
rect 45050 24194 48968 24362
tri 48968 24194 49180 24406 sw
tri 49265 24194 49477 24406 ne
rect 49477 24194 70613 24406
rect 45050 24080 49180 24194
rect 40656 23948 44768 24080
rect 38624 23656 40364 23948
tri 40364 23656 40656 23948 sw
tri 40656 23656 40948 23948 ne
rect 40948 23798 44768 23948
tri 44768 23798 45050 24080 sw
tri 45050 23798 45332 24080 ne
rect 45332 23897 49180 24080
tri 49180 23897 49477 24194 sw
tri 49477 23897 49774 24194 ne
rect 49774 23897 70613 24194
rect 45332 23798 49477 23897
rect 40948 23656 45050 23798
rect 38624 23364 40656 23656
tri 40656 23364 40948 23656 sw
tri 40948 23364 41240 23656 ne
rect 41240 23516 45050 23656
tri 45050 23516 45332 23798 sw
tri 45332 23516 45614 23798 ne
rect 45614 23600 49477 23798
tri 49477 23600 49774 23897 sw
tri 49774 23600 50071 23897 ne
rect 50071 23706 70613 23897
rect 70669 23706 71000 24906
rect 50071 23600 71000 23706
rect 45614 23516 49774 23600
rect 41240 23364 45332 23516
rect 38624 23072 40948 23364
tri 40948 23072 41240 23364 sw
tri 41240 23072 41532 23364 ne
rect 41532 23234 45332 23364
tri 45332 23234 45614 23516 sw
tri 45614 23234 45896 23516 ne
rect 45896 23400 49774 23516
tri 49774 23400 49974 23600 sw
rect 45896 23234 71000 23400
rect 41532 23072 45614 23234
rect 38624 22780 41240 23072
tri 41240 22780 41532 23072 sw
tri 41532 22780 41824 23072 ne
rect 41824 22952 45614 23072
tri 45614 22952 45896 23234 sw
tri 45896 22952 46178 23234 ne
rect 46178 22952 71000 23234
rect 41824 22854 45896 22952
tri 45896 22854 45994 22952 sw
tri 46178 22854 46276 22952 ne
rect 46276 22854 71000 22952
rect 41824 22780 45994 22854
rect 38624 22488 41532 22780
tri 41532 22488 41824 22780 sw
tri 41824 22488 42116 22780 ne
rect 42116 22572 45994 22780
tri 45994 22572 46276 22854 sw
tri 46276 22572 46558 22854 ne
rect 46558 22572 71000 22854
rect 42116 22488 46276 22572
rect 38624 22196 41824 22488
tri 41824 22196 42116 22488 sw
tri 42116 22196 42408 22488 ne
rect 42408 22290 46276 22488
tri 46276 22290 46558 22572 sw
tri 46558 22290 46840 22572 ne
rect 46840 22290 71000 22572
rect 42408 22196 46558 22290
rect 38624 22028 42116 22196
tri 42116 22028 42284 22196 sw
tri 42408 22028 42576 22196 ne
rect 42576 22028 46558 22196
rect 38624 21736 42284 22028
tri 42284 21736 42576 22028 sw
tri 42576 21736 42868 22028 ne
rect 42868 22008 46558 22028
tri 46558 22008 46840 22290 sw
tri 46840 22008 47122 22290 ne
rect 47122 22008 71000 22290
rect 42868 21736 46840 22008
rect 38624 21444 42576 21736
tri 42576 21444 42868 21736 sw
tri 42868 21444 43160 21736 ne
rect 43160 21726 46840 21736
tri 46840 21726 47122 22008 sw
tri 47122 21726 47404 22008 ne
rect 47404 21726 71000 22008
rect 43160 21444 47122 21726
tri 47122 21444 47404 21726 sw
tri 47404 21444 47686 21726 ne
rect 47686 21444 71000 21726
tri 38624 17200 42868 21444 ne
tri 42868 21152 43160 21444 sw
tri 43160 21152 43452 21444 ne
rect 43452 21162 47404 21444
tri 47404 21162 47686 21444 sw
tri 47686 21162 47968 21444 ne
rect 47968 21162 71000 21444
rect 43452 21152 47686 21162
rect 42868 20860 43160 21152
tri 43160 20860 43452 21152 sw
tri 43452 20860 43744 21152 ne
rect 43744 20964 47686 21152
tri 47686 20964 47884 21162 sw
tri 47968 20964 48166 21162 ne
rect 48166 20964 71000 21162
rect 43744 20860 47884 20964
rect 42868 20568 43452 20860
tri 43452 20568 43744 20860 sw
tri 43744 20568 44036 20860 ne
rect 44036 20682 47884 20860
tri 47884 20682 48166 20964 sw
tri 48166 20682 48448 20964 ne
rect 48448 20682 71000 20964
rect 44036 20568 48166 20682
rect 42868 20276 43744 20568
tri 43744 20276 44036 20568 sw
tri 44036 20276 44328 20568 ne
rect 44328 20400 48166 20568
tri 48166 20400 48448 20682 sw
tri 48448 20400 48730 20682 ne
rect 48730 20400 71000 20682
rect 44328 20276 48448 20400
rect 42868 19984 44036 20276
tri 44036 19984 44328 20276 sw
tri 44328 19984 44620 20276 ne
rect 44620 20200 48448 20276
tri 48448 20200 48648 20400 sw
rect 44620 19984 71000 20200
rect 42868 19704 44328 19984
tri 44328 19704 44608 19984 sw
tri 44620 19704 44900 19984 ne
rect 44900 19704 71000 19984
rect 42868 19412 44608 19704
tri 44608 19412 44900 19704 sw
tri 44900 19412 45192 19704 ne
rect 45192 19412 71000 19704
rect 42868 19120 44900 19412
tri 44900 19120 45192 19412 sw
tri 45192 19120 45484 19412 ne
rect 45484 19120 71000 19412
rect 42868 18828 45192 19120
tri 45192 18828 45484 19120 sw
tri 45484 18828 45776 19120 ne
rect 45776 18828 71000 19120
rect 42868 18536 45484 18828
tri 45484 18536 45776 18828 sw
tri 45776 18536 46068 18828 ne
rect 46068 18536 71000 18828
rect 42868 18244 45776 18536
tri 45776 18244 46068 18536 sw
tri 46068 18244 46360 18536 ne
rect 46360 18244 71000 18536
rect 42868 17952 46068 18244
tri 46068 17952 46360 18244 sw
tri 46360 17952 46652 18244 ne
rect 46652 17952 71000 18244
rect 42868 17784 46360 17952
tri 46360 17784 46528 17952 sw
tri 46652 17784 46820 17952 ne
rect 46820 17784 71000 17952
rect 42868 17492 46528 17784
tri 46528 17492 46820 17784 sw
tri 46820 17492 47112 17784 ne
rect 47112 17492 71000 17784
rect 42868 17200 46820 17492
tri 46820 17200 47112 17492 sw
tri 47112 17200 47404 17492 ne
rect 47404 17200 71000 17492
tri 42868 14000 46068 17200 ne
rect 46068 17000 47112 17200
tri 47112 17000 47312 17200 sw
rect 46068 14000 71000 17000
<< labels >>
rlabel metal3 s 70454 64211 70454 64211 4 VSS
port 1 nsew
rlabel metal3 s 70454 62776 70454 62776 4 VDD
port 2 nsew
rlabel metal3 s 70454 61011 70454 61011 4 DVSS
port 3 nsew
rlabel metal3 s 70454 65976 70454 65976 4 DVSS
port 3 nsew
rlabel metal3 s 70454 69002 70454 69002 4 DVSS
port 3 nsew
rlabel metal3 s 70454 67411 70454 67411 4 DVDD
port 4 nsew
rlabel metal3 s 70454 59576 70454 59576 4 DVDD
port 4 nsew
rlabel metal3 s 70454 57811 70454 57811 4 DVSS
port 3 nsew
rlabel metal3 s 70454 56376 70454 56376 4 DVDD
port 4 nsew
rlabel metal3 s 70454 54611 70454 54611 4 DVDD
port 4 nsew
rlabel metal3 s 70454 53176 70454 53176 4 DVDD
port 4 nsew
rlabel metal3 s 70559 51411 70559 51411 4 VDD
port 2 nsew
rlabel metal3 s 70559 49976 70559 49976 4 VSS
port 1 nsew
rlabel metal3 s 70454 47548 70454 47548 4 DVSS
port 3 nsew
rlabel metal3 s 70454 44321 70454 44321 4 DVDD
port 4 nsew
rlabel metal3 s 70454 40295 70454 40295 4 DVSS
port 3 nsew
rlabel metal3 s 70454 41930 70454 41930 4 DVDD
port 4 nsew
rlabel metal3 s 70454 37912 70454 37912 4 DVDD
port 4 nsew
rlabel metal3 s 70454 34676 70454 34676 4 DVDD
port 4 nsew
rlabel metal3 s 70454 31562 70454 31562 4 DVDD
port 4 nsew
rlabel metal3 s 70454 28347 70454 28347 4 DVDD
port 4 nsew
rlabel metal3 s 70454 26053 70454 26053 4 DVSS
port 3 nsew
rlabel metal3 s 70454 24237 70454 24237 4 DVDD
port 4 nsew
rlabel metal3 s 70454 21860 70454 21860 4 DVSS
port 3 nsew
rlabel metal3 s 70385 18874 70385 18874 4 DVSS
port 3 nsew
rlabel metal3 s 70432 15703 70432 15703 4 DVSS
port 3 nsew
<< properties >>
string FIXED_BBOX 0 0 71000 71000
<< end >>
