magic
tech gf180mcuD
magscale 1 10
timestamp 1764347740
<< nwell >>
rect -1730 9497 11766 10481
rect -1730 -15 -500 9497
rect 10573 -15 11766 9497
rect -1730 -583 11766 -15
<< psubdiff >>
rect -458 8756 10536 9430
rect -458 8300 -118 8756
rect -458 54 -396 8300
rect -150 322 -118 8300
rect 10146 8322 10536 8756
rect 10146 8300 10541 8322
rect 10146 322 10173 8300
rect -150 300 10173 322
rect -150 54 11 300
rect 10057 54 10173 300
rect 10519 54 10541 8300
rect -458 32 10541 54
<< nsubdiff >>
rect -1647 10376 11683 10398
rect -1647 9602 -436 10376
rect 10510 9602 11683 10376
rect -1647 9580 11683 9602
rect -1647 8368 -583 9580
rect -1647 -478 -1587 8368
rect -605 -98 -583 8368
rect 10656 8368 11683 9580
rect 10656 -98 10678 8368
rect -605 -120 10678 -98
rect -605 -478 -436 -120
rect 10510 -478 10678 -120
rect 11660 -478 11683 8368
rect -1647 -500 11683 -478
<< psubdiffcont >>
rect -396 54 -150 8300
rect 11 54 10057 300
rect 10173 54 10519 8300
<< nsubdiffcont >>
rect -436 9602 10510 10376
rect -1587 -478 -605 8368
rect -436 -478 10510 -120
rect 10678 -478 11660 8368
<< metal1 >>
rect -447 10376 10521 10387
rect -447 9602 -436 10376
rect 10510 9602 10521 10376
rect -447 9591 10521 9602
rect -1598 8368 -594 8388
rect -1598 -478 -1587 8368
rect -605 -109 -594 8368
rect -457 8300 111 8396
rect -457 54 -396 8300
rect -150 311 111 8300
rect 9962 8300 10530 8397
rect 9962 311 10173 8300
rect -150 300 10173 311
rect -150 54 11 300
rect 10057 54 10173 300
rect 10519 54 10530 8300
rect -457 43 10530 54
rect 10666 8368 11670 8410
rect 10666 -109 10678 8368
rect -605 -120 10678 -109
rect -605 -478 -436 -120
rect 10510 -478 10678 -120
rect 11660 -478 11670 8368
rect -1598 -489 11670 -478
<< end >>
