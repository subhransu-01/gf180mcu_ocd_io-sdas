magic
tech gf180mcuD
magscale 1 10
timestamp 1764277317
<< nwell >>
rect 2167 27624 10795 29168
<< hvnmos >>
rect 4129 26006 4269 27006
rect 5191 26006 5331 27006
rect 5435 26006 5575 27006
rect 5679 26006 5819 27006
rect 5923 26006 6063 27006
rect 6167 26006 6307 27006
rect 6411 26006 6551 27006
rect 6655 26006 6795 27006
rect 6899 26006 7039 27006
rect 7143 26006 7283 27006
rect 7387 26006 7527 27006
rect 7631 26006 7771 27006
rect 7875 26006 8015 27006
<< hvpmos >>
rect 2665 27789 2805 28789
rect 2909 27789 3049 28789
rect 3153 27789 3293 28789
rect 3397 27789 3537 28789
rect 3641 27789 3781 28789
rect 3885 27789 4025 28789
rect 4129 27789 4269 28789
rect 4545 27789 4685 28789
rect 4789 27789 4929 28789
rect 5033 27789 5173 28789
rect 5277 27789 5417 28789
rect 5521 27789 5661 28789
rect 5765 27789 5905 28789
rect 6009 27789 6149 28789
rect 6253 27789 6393 28789
rect 6497 27789 6637 28789
rect 6741 27789 6881 28789
rect 6985 27789 7125 28789
rect 7229 27789 7369 28789
rect 7473 27789 7613 28789
rect 7717 27789 7857 28789
rect 7961 27789 8101 28789
rect 8205 27789 8345 28789
rect 8449 27789 8589 28789
rect 8693 27789 8833 28789
rect 8937 27789 9077 28789
rect 9181 27789 9321 28789
rect 9425 27789 9565 28789
rect 9669 27789 9809 28789
rect 9913 27789 10053 28789
rect 10157 27789 10297 28789
<< mvndiff >>
rect 4041 26993 4129 27006
rect 4041 26947 4054 26993
rect 4100 26947 4129 26993
rect 4041 26890 4129 26947
rect 4041 26844 4054 26890
rect 4100 26844 4129 26890
rect 4041 26787 4129 26844
rect 4041 26741 4054 26787
rect 4100 26741 4129 26787
rect 4041 26684 4129 26741
rect 4041 26638 4054 26684
rect 4100 26638 4129 26684
rect 4041 26581 4129 26638
rect 4041 26535 4054 26581
rect 4100 26535 4129 26581
rect 4041 26478 4129 26535
rect 4041 26432 4054 26478
rect 4100 26432 4129 26478
rect 4041 26375 4129 26432
rect 4041 26329 4054 26375
rect 4100 26329 4129 26375
rect 4041 26272 4129 26329
rect 4041 26226 4054 26272
rect 4100 26226 4129 26272
rect 4041 26169 4129 26226
rect 4041 26123 4054 26169
rect 4100 26123 4129 26169
rect 4041 26065 4129 26123
rect 4041 26019 4054 26065
rect 4100 26019 4129 26065
rect 4041 26006 4129 26019
rect 4269 26993 4357 27006
rect 4269 26947 4298 26993
rect 4344 26947 4357 26993
rect 4269 26890 4357 26947
rect 4269 26844 4298 26890
rect 4344 26844 4357 26890
rect 4269 26787 4357 26844
rect 4269 26741 4298 26787
rect 4344 26741 4357 26787
rect 4269 26684 4357 26741
rect 4269 26638 4298 26684
rect 4344 26638 4357 26684
rect 4269 26581 4357 26638
rect 4269 26535 4298 26581
rect 4344 26535 4357 26581
rect 4269 26478 4357 26535
rect 4269 26432 4298 26478
rect 4344 26432 4357 26478
rect 4269 26375 4357 26432
rect 4269 26329 4298 26375
rect 4344 26329 4357 26375
rect 4269 26272 4357 26329
rect 4269 26226 4298 26272
rect 4344 26226 4357 26272
rect 4269 26169 4357 26226
rect 4269 26123 4298 26169
rect 4344 26123 4357 26169
rect 4269 26065 4357 26123
rect 4269 26019 4298 26065
rect 4344 26019 4357 26065
rect 4269 26006 4357 26019
rect 5103 26993 5191 27006
rect 5103 26947 5116 26993
rect 5162 26947 5191 26993
rect 5103 26890 5191 26947
rect 5103 26844 5116 26890
rect 5162 26844 5191 26890
rect 5103 26787 5191 26844
rect 5103 26741 5116 26787
rect 5162 26741 5191 26787
rect 5103 26684 5191 26741
rect 5103 26638 5116 26684
rect 5162 26638 5191 26684
rect 5103 26581 5191 26638
rect 5103 26535 5116 26581
rect 5162 26535 5191 26581
rect 5103 26478 5191 26535
rect 5103 26432 5116 26478
rect 5162 26432 5191 26478
rect 5103 26375 5191 26432
rect 5103 26329 5116 26375
rect 5162 26329 5191 26375
rect 5103 26272 5191 26329
rect 5103 26226 5116 26272
rect 5162 26226 5191 26272
rect 5103 26169 5191 26226
rect 5103 26123 5116 26169
rect 5162 26123 5191 26169
rect 5103 26065 5191 26123
rect 5103 26019 5116 26065
rect 5162 26019 5191 26065
rect 5103 26006 5191 26019
rect 5331 26993 5435 27006
rect 5331 26947 5360 26993
rect 5406 26947 5435 26993
rect 5331 26890 5435 26947
rect 5331 26844 5360 26890
rect 5406 26844 5435 26890
rect 5331 26787 5435 26844
rect 5331 26741 5360 26787
rect 5406 26741 5435 26787
rect 5331 26684 5435 26741
rect 5331 26638 5360 26684
rect 5406 26638 5435 26684
rect 5331 26581 5435 26638
rect 5331 26535 5360 26581
rect 5406 26535 5435 26581
rect 5331 26478 5435 26535
rect 5331 26432 5360 26478
rect 5406 26432 5435 26478
rect 5331 26375 5435 26432
rect 5331 26329 5360 26375
rect 5406 26329 5435 26375
rect 5331 26272 5435 26329
rect 5331 26226 5360 26272
rect 5406 26226 5435 26272
rect 5331 26169 5435 26226
rect 5331 26123 5360 26169
rect 5406 26123 5435 26169
rect 5331 26065 5435 26123
rect 5331 26019 5360 26065
rect 5406 26019 5435 26065
rect 5331 26006 5435 26019
rect 5575 26993 5679 27006
rect 5575 26947 5604 26993
rect 5650 26947 5679 26993
rect 5575 26890 5679 26947
rect 5575 26844 5604 26890
rect 5650 26844 5679 26890
rect 5575 26787 5679 26844
rect 5575 26741 5604 26787
rect 5650 26741 5679 26787
rect 5575 26684 5679 26741
rect 5575 26638 5604 26684
rect 5650 26638 5679 26684
rect 5575 26581 5679 26638
rect 5575 26535 5604 26581
rect 5650 26535 5679 26581
rect 5575 26478 5679 26535
rect 5575 26432 5604 26478
rect 5650 26432 5679 26478
rect 5575 26375 5679 26432
rect 5575 26329 5604 26375
rect 5650 26329 5679 26375
rect 5575 26272 5679 26329
rect 5575 26226 5604 26272
rect 5650 26226 5679 26272
rect 5575 26169 5679 26226
rect 5575 26123 5604 26169
rect 5650 26123 5679 26169
rect 5575 26065 5679 26123
rect 5575 26019 5604 26065
rect 5650 26019 5679 26065
rect 5575 26006 5679 26019
rect 5819 26993 5923 27006
rect 5819 26947 5848 26993
rect 5894 26947 5923 26993
rect 5819 26890 5923 26947
rect 5819 26844 5848 26890
rect 5894 26844 5923 26890
rect 5819 26787 5923 26844
rect 5819 26741 5848 26787
rect 5894 26741 5923 26787
rect 5819 26684 5923 26741
rect 5819 26638 5848 26684
rect 5894 26638 5923 26684
rect 5819 26581 5923 26638
rect 5819 26535 5848 26581
rect 5894 26535 5923 26581
rect 5819 26478 5923 26535
rect 5819 26432 5848 26478
rect 5894 26432 5923 26478
rect 5819 26375 5923 26432
rect 5819 26329 5848 26375
rect 5894 26329 5923 26375
rect 5819 26272 5923 26329
rect 5819 26226 5848 26272
rect 5894 26226 5923 26272
rect 5819 26169 5923 26226
rect 5819 26123 5848 26169
rect 5894 26123 5923 26169
rect 5819 26065 5923 26123
rect 5819 26019 5848 26065
rect 5894 26019 5923 26065
rect 5819 26006 5923 26019
rect 6063 26993 6167 27006
rect 6063 26947 6092 26993
rect 6138 26947 6167 26993
rect 6063 26890 6167 26947
rect 6063 26844 6092 26890
rect 6138 26844 6167 26890
rect 6063 26787 6167 26844
rect 6063 26741 6092 26787
rect 6138 26741 6167 26787
rect 6063 26684 6167 26741
rect 6063 26638 6092 26684
rect 6138 26638 6167 26684
rect 6063 26581 6167 26638
rect 6063 26535 6092 26581
rect 6138 26535 6167 26581
rect 6063 26478 6167 26535
rect 6063 26432 6092 26478
rect 6138 26432 6167 26478
rect 6063 26375 6167 26432
rect 6063 26329 6092 26375
rect 6138 26329 6167 26375
rect 6063 26272 6167 26329
rect 6063 26226 6092 26272
rect 6138 26226 6167 26272
rect 6063 26169 6167 26226
rect 6063 26123 6092 26169
rect 6138 26123 6167 26169
rect 6063 26065 6167 26123
rect 6063 26019 6092 26065
rect 6138 26019 6167 26065
rect 6063 26006 6167 26019
rect 6307 26993 6411 27006
rect 6307 26947 6336 26993
rect 6382 26947 6411 26993
rect 6307 26890 6411 26947
rect 6307 26844 6336 26890
rect 6382 26844 6411 26890
rect 6307 26787 6411 26844
rect 6307 26741 6336 26787
rect 6382 26741 6411 26787
rect 6307 26684 6411 26741
rect 6307 26638 6336 26684
rect 6382 26638 6411 26684
rect 6307 26581 6411 26638
rect 6307 26535 6336 26581
rect 6382 26535 6411 26581
rect 6307 26478 6411 26535
rect 6307 26432 6336 26478
rect 6382 26432 6411 26478
rect 6307 26375 6411 26432
rect 6307 26329 6336 26375
rect 6382 26329 6411 26375
rect 6307 26272 6411 26329
rect 6307 26226 6336 26272
rect 6382 26226 6411 26272
rect 6307 26169 6411 26226
rect 6307 26123 6336 26169
rect 6382 26123 6411 26169
rect 6307 26065 6411 26123
rect 6307 26019 6336 26065
rect 6382 26019 6411 26065
rect 6307 26006 6411 26019
rect 6551 26993 6655 27006
rect 6551 26947 6580 26993
rect 6626 26947 6655 26993
rect 6551 26890 6655 26947
rect 6551 26844 6580 26890
rect 6626 26844 6655 26890
rect 6551 26787 6655 26844
rect 6551 26741 6580 26787
rect 6626 26741 6655 26787
rect 6551 26684 6655 26741
rect 6551 26638 6580 26684
rect 6626 26638 6655 26684
rect 6551 26581 6655 26638
rect 6551 26535 6580 26581
rect 6626 26535 6655 26581
rect 6551 26478 6655 26535
rect 6551 26432 6580 26478
rect 6626 26432 6655 26478
rect 6551 26375 6655 26432
rect 6551 26329 6580 26375
rect 6626 26329 6655 26375
rect 6551 26272 6655 26329
rect 6551 26226 6580 26272
rect 6626 26226 6655 26272
rect 6551 26169 6655 26226
rect 6551 26123 6580 26169
rect 6626 26123 6655 26169
rect 6551 26065 6655 26123
rect 6551 26019 6580 26065
rect 6626 26019 6655 26065
rect 6551 26006 6655 26019
rect 6795 26993 6899 27006
rect 6795 26947 6824 26993
rect 6870 26947 6899 26993
rect 6795 26890 6899 26947
rect 6795 26844 6824 26890
rect 6870 26844 6899 26890
rect 6795 26787 6899 26844
rect 6795 26741 6824 26787
rect 6870 26741 6899 26787
rect 6795 26684 6899 26741
rect 6795 26638 6824 26684
rect 6870 26638 6899 26684
rect 6795 26581 6899 26638
rect 6795 26535 6824 26581
rect 6870 26535 6899 26581
rect 6795 26478 6899 26535
rect 6795 26432 6824 26478
rect 6870 26432 6899 26478
rect 6795 26375 6899 26432
rect 6795 26329 6824 26375
rect 6870 26329 6899 26375
rect 6795 26272 6899 26329
rect 6795 26226 6824 26272
rect 6870 26226 6899 26272
rect 6795 26169 6899 26226
rect 6795 26123 6824 26169
rect 6870 26123 6899 26169
rect 6795 26065 6899 26123
rect 6795 26019 6824 26065
rect 6870 26019 6899 26065
rect 6795 26006 6899 26019
rect 7039 26993 7143 27006
rect 7039 26947 7068 26993
rect 7114 26947 7143 26993
rect 7039 26890 7143 26947
rect 7039 26844 7068 26890
rect 7114 26844 7143 26890
rect 7039 26787 7143 26844
rect 7039 26741 7068 26787
rect 7114 26741 7143 26787
rect 7039 26684 7143 26741
rect 7039 26638 7068 26684
rect 7114 26638 7143 26684
rect 7039 26581 7143 26638
rect 7039 26535 7068 26581
rect 7114 26535 7143 26581
rect 7039 26478 7143 26535
rect 7039 26432 7068 26478
rect 7114 26432 7143 26478
rect 7039 26375 7143 26432
rect 7039 26329 7068 26375
rect 7114 26329 7143 26375
rect 7039 26272 7143 26329
rect 7039 26226 7068 26272
rect 7114 26226 7143 26272
rect 7039 26169 7143 26226
rect 7039 26123 7068 26169
rect 7114 26123 7143 26169
rect 7039 26065 7143 26123
rect 7039 26019 7068 26065
rect 7114 26019 7143 26065
rect 7039 26006 7143 26019
rect 7283 26993 7387 27006
rect 7283 26947 7312 26993
rect 7358 26947 7387 26993
rect 7283 26890 7387 26947
rect 7283 26844 7312 26890
rect 7358 26844 7387 26890
rect 7283 26787 7387 26844
rect 7283 26741 7312 26787
rect 7358 26741 7387 26787
rect 7283 26684 7387 26741
rect 7283 26638 7312 26684
rect 7358 26638 7387 26684
rect 7283 26581 7387 26638
rect 7283 26535 7312 26581
rect 7358 26535 7387 26581
rect 7283 26478 7387 26535
rect 7283 26432 7312 26478
rect 7358 26432 7387 26478
rect 7283 26375 7387 26432
rect 7283 26329 7312 26375
rect 7358 26329 7387 26375
rect 7283 26272 7387 26329
rect 7283 26226 7312 26272
rect 7358 26226 7387 26272
rect 7283 26169 7387 26226
rect 7283 26123 7312 26169
rect 7358 26123 7387 26169
rect 7283 26065 7387 26123
rect 7283 26019 7312 26065
rect 7358 26019 7387 26065
rect 7283 26006 7387 26019
rect 7527 26993 7631 27006
rect 7527 26947 7556 26993
rect 7602 26947 7631 26993
rect 7527 26890 7631 26947
rect 7527 26844 7556 26890
rect 7602 26844 7631 26890
rect 7527 26787 7631 26844
rect 7527 26741 7556 26787
rect 7602 26741 7631 26787
rect 7527 26684 7631 26741
rect 7527 26638 7556 26684
rect 7602 26638 7631 26684
rect 7527 26581 7631 26638
rect 7527 26535 7556 26581
rect 7602 26535 7631 26581
rect 7527 26478 7631 26535
rect 7527 26432 7556 26478
rect 7602 26432 7631 26478
rect 7527 26375 7631 26432
rect 7527 26329 7556 26375
rect 7602 26329 7631 26375
rect 7527 26272 7631 26329
rect 7527 26226 7556 26272
rect 7602 26226 7631 26272
rect 7527 26169 7631 26226
rect 7527 26123 7556 26169
rect 7602 26123 7631 26169
rect 7527 26065 7631 26123
rect 7527 26019 7556 26065
rect 7602 26019 7631 26065
rect 7527 26006 7631 26019
rect 7771 26993 7875 27006
rect 7771 26947 7800 26993
rect 7846 26947 7875 26993
rect 7771 26890 7875 26947
rect 7771 26844 7800 26890
rect 7846 26844 7875 26890
rect 7771 26787 7875 26844
rect 7771 26741 7800 26787
rect 7846 26741 7875 26787
rect 7771 26684 7875 26741
rect 7771 26638 7800 26684
rect 7846 26638 7875 26684
rect 7771 26581 7875 26638
rect 7771 26535 7800 26581
rect 7846 26535 7875 26581
rect 7771 26478 7875 26535
rect 7771 26432 7800 26478
rect 7846 26432 7875 26478
rect 7771 26375 7875 26432
rect 7771 26329 7800 26375
rect 7846 26329 7875 26375
rect 7771 26272 7875 26329
rect 7771 26226 7800 26272
rect 7846 26226 7875 26272
rect 7771 26169 7875 26226
rect 7771 26123 7800 26169
rect 7846 26123 7875 26169
rect 7771 26065 7875 26123
rect 7771 26019 7800 26065
rect 7846 26019 7875 26065
rect 7771 26006 7875 26019
rect 8015 26993 8103 27006
rect 8015 26947 8044 26993
rect 8090 26947 8103 26993
rect 8015 26890 8103 26947
rect 8015 26844 8044 26890
rect 8090 26844 8103 26890
rect 8015 26787 8103 26844
rect 8015 26741 8044 26787
rect 8090 26741 8103 26787
rect 8015 26684 8103 26741
rect 8015 26638 8044 26684
rect 8090 26638 8103 26684
rect 8015 26581 8103 26638
rect 8015 26535 8044 26581
rect 8090 26535 8103 26581
rect 8015 26478 8103 26535
rect 8015 26432 8044 26478
rect 8090 26432 8103 26478
rect 8015 26375 8103 26432
rect 8015 26329 8044 26375
rect 8090 26329 8103 26375
rect 8015 26272 8103 26329
rect 8015 26226 8044 26272
rect 8090 26226 8103 26272
rect 8015 26169 8103 26226
rect 8015 26123 8044 26169
rect 8090 26123 8103 26169
rect 8015 26065 8103 26123
rect 8015 26019 8044 26065
rect 8090 26019 8103 26065
rect 8015 26006 8103 26019
<< mvpdiff >>
rect 2577 28776 2665 28789
rect 2577 28730 2590 28776
rect 2636 28730 2665 28776
rect 2577 28673 2665 28730
rect 2577 28627 2590 28673
rect 2636 28627 2665 28673
rect 2577 28570 2665 28627
rect 2577 28524 2590 28570
rect 2636 28524 2665 28570
rect 2577 28467 2665 28524
rect 2577 28421 2590 28467
rect 2636 28421 2665 28467
rect 2577 28364 2665 28421
rect 2577 28318 2590 28364
rect 2636 28318 2665 28364
rect 2577 28261 2665 28318
rect 2577 28215 2590 28261
rect 2636 28215 2665 28261
rect 2577 28158 2665 28215
rect 2577 28112 2590 28158
rect 2636 28112 2665 28158
rect 2577 28055 2665 28112
rect 2577 28009 2590 28055
rect 2636 28009 2665 28055
rect 2577 27952 2665 28009
rect 2577 27906 2590 27952
rect 2636 27906 2665 27952
rect 2577 27848 2665 27906
rect 2577 27802 2590 27848
rect 2636 27802 2665 27848
rect 2577 27789 2665 27802
rect 2805 28776 2909 28789
rect 2805 28730 2834 28776
rect 2880 28730 2909 28776
rect 2805 28673 2909 28730
rect 2805 28627 2834 28673
rect 2880 28627 2909 28673
rect 2805 28570 2909 28627
rect 2805 28524 2834 28570
rect 2880 28524 2909 28570
rect 2805 28467 2909 28524
rect 2805 28421 2834 28467
rect 2880 28421 2909 28467
rect 2805 28364 2909 28421
rect 2805 28318 2834 28364
rect 2880 28318 2909 28364
rect 2805 28261 2909 28318
rect 2805 28215 2834 28261
rect 2880 28215 2909 28261
rect 2805 28158 2909 28215
rect 2805 28112 2834 28158
rect 2880 28112 2909 28158
rect 2805 28055 2909 28112
rect 2805 28009 2834 28055
rect 2880 28009 2909 28055
rect 2805 27952 2909 28009
rect 2805 27906 2834 27952
rect 2880 27906 2909 27952
rect 2805 27848 2909 27906
rect 2805 27802 2834 27848
rect 2880 27802 2909 27848
rect 2805 27789 2909 27802
rect 3049 28776 3153 28789
rect 3049 28730 3078 28776
rect 3124 28730 3153 28776
rect 3049 28673 3153 28730
rect 3049 28627 3078 28673
rect 3124 28627 3153 28673
rect 3049 28570 3153 28627
rect 3049 28524 3078 28570
rect 3124 28524 3153 28570
rect 3049 28467 3153 28524
rect 3049 28421 3078 28467
rect 3124 28421 3153 28467
rect 3049 28364 3153 28421
rect 3049 28318 3078 28364
rect 3124 28318 3153 28364
rect 3049 28261 3153 28318
rect 3049 28215 3078 28261
rect 3124 28215 3153 28261
rect 3049 28158 3153 28215
rect 3049 28112 3078 28158
rect 3124 28112 3153 28158
rect 3049 28055 3153 28112
rect 3049 28009 3078 28055
rect 3124 28009 3153 28055
rect 3049 27952 3153 28009
rect 3049 27906 3078 27952
rect 3124 27906 3153 27952
rect 3049 27848 3153 27906
rect 3049 27802 3078 27848
rect 3124 27802 3153 27848
rect 3049 27789 3153 27802
rect 3293 28776 3397 28789
rect 3293 28730 3322 28776
rect 3368 28730 3397 28776
rect 3293 28673 3397 28730
rect 3293 28627 3322 28673
rect 3368 28627 3397 28673
rect 3293 28570 3397 28627
rect 3293 28524 3322 28570
rect 3368 28524 3397 28570
rect 3293 28467 3397 28524
rect 3293 28421 3322 28467
rect 3368 28421 3397 28467
rect 3293 28364 3397 28421
rect 3293 28318 3322 28364
rect 3368 28318 3397 28364
rect 3293 28261 3397 28318
rect 3293 28215 3322 28261
rect 3368 28215 3397 28261
rect 3293 28158 3397 28215
rect 3293 28112 3322 28158
rect 3368 28112 3397 28158
rect 3293 28055 3397 28112
rect 3293 28009 3322 28055
rect 3368 28009 3397 28055
rect 3293 27952 3397 28009
rect 3293 27906 3322 27952
rect 3368 27906 3397 27952
rect 3293 27848 3397 27906
rect 3293 27802 3322 27848
rect 3368 27802 3397 27848
rect 3293 27789 3397 27802
rect 3537 28776 3641 28789
rect 3537 28730 3566 28776
rect 3612 28730 3641 28776
rect 3537 28673 3641 28730
rect 3537 28627 3566 28673
rect 3612 28627 3641 28673
rect 3537 28570 3641 28627
rect 3537 28524 3566 28570
rect 3612 28524 3641 28570
rect 3537 28467 3641 28524
rect 3537 28421 3566 28467
rect 3612 28421 3641 28467
rect 3537 28364 3641 28421
rect 3537 28318 3566 28364
rect 3612 28318 3641 28364
rect 3537 28261 3641 28318
rect 3537 28215 3566 28261
rect 3612 28215 3641 28261
rect 3537 28158 3641 28215
rect 3537 28112 3566 28158
rect 3612 28112 3641 28158
rect 3537 28055 3641 28112
rect 3537 28009 3566 28055
rect 3612 28009 3641 28055
rect 3537 27952 3641 28009
rect 3537 27906 3566 27952
rect 3612 27906 3641 27952
rect 3537 27848 3641 27906
rect 3537 27802 3566 27848
rect 3612 27802 3641 27848
rect 3537 27789 3641 27802
rect 3781 28776 3885 28789
rect 3781 28730 3810 28776
rect 3856 28730 3885 28776
rect 3781 28673 3885 28730
rect 3781 28627 3810 28673
rect 3856 28627 3885 28673
rect 3781 28570 3885 28627
rect 3781 28524 3810 28570
rect 3856 28524 3885 28570
rect 3781 28467 3885 28524
rect 3781 28421 3810 28467
rect 3856 28421 3885 28467
rect 3781 28364 3885 28421
rect 3781 28318 3810 28364
rect 3856 28318 3885 28364
rect 3781 28261 3885 28318
rect 3781 28215 3810 28261
rect 3856 28215 3885 28261
rect 3781 28158 3885 28215
rect 3781 28112 3810 28158
rect 3856 28112 3885 28158
rect 3781 28055 3885 28112
rect 3781 28009 3810 28055
rect 3856 28009 3885 28055
rect 3781 27952 3885 28009
rect 3781 27906 3810 27952
rect 3856 27906 3885 27952
rect 3781 27848 3885 27906
rect 3781 27802 3810 27848
rect 3856 27802 3885 27848
rect 3781 27789 3885 27802
rect 4025 28776 4129 28789
rect 4025 28730 4054 28776
rect 4100 28730 4129 28776
rect 4025 28673 4129 28730
rect 4025 28627 4054 28673
rect 4100 28627 4129 28673
rect 4025 28570 4129 28627
rect 4025 28524 4054 28570
rect 4100 28524 4129 28570
rect 4025 28467 4129 28524
rect 4025 28421 4054 28467
rect 4100 28421 4129 28467
rect 4025 28364 4129 28421
rect 4025 28318 4054 28364
rect 4100 28318 4129 28364
rect 4025 28261 4129 28318
rect 4025 28215 4054 28261
rect 4100 28215 4129 28261
rect 4025 28158 4129 28215
rect 4025 28112 4054 28158
rect 4100 28112 4129 28158
rect 4025 28055 4129 28112
rect 4025 28009 4054 28055
rect 4100 28009 4129 28055
rect 4025 27952 4129 28009
rect 4025 27906 4054 27952
rect 4100 27906 4129 27952
rect 4025 27848 4129 27906
rect 4025 27802 4054 27848
rect 4100 27802 4129 27848
rect 4025 27789 4129 27802
rect 4269 28776 4357 28789
rect 4269 28730 4298 28776
rect 4344 28730 4357 28776
rect 4269 28673 4357 28730
rect 4269 28627 4298 28673
rect 4344 28627 4357 28673
rect 4269 28570 4357 28627
rect 4269 28524 4298 28570
rect 4344 28524 4357 28570
rect 4269 28467 4357 28524
rect 4269 28421 4298 28467
rect 4344 28421 4357 28467
rect 4269 28364 4357 28421
rect 4269 28318 4298 28364
rect 4344 28318 4357 28364
rect 4269 28261 4357 28318
rect 4269 28215 4298 28261
rect 4344 28215 4357 28261
rect 4269 28158 4357 28215
rect 4269 28112 4298 28158
rect 4344 28112 4357 28158
rect 4269 28055 4357 28112
rect 4269 28009 4298 28055
rect 4344 28009 4357 28055
rect 4269 27952 4357 28009
rect 4269 27906 4298 27952
rect 4344 27906 4357 27952
rect 4269 27848 4357 27906
rect 4269 27802 4298 27848
rect 4344 27802 4357 27848
rect 4269 27789 4357 27802
rect 4457 28776 4545 28789
rect 4457 28730 4470 28776
rect 4516 28730 4545 28776
rect 4457 28673 4545 28730
rect 4457 28627 4470 28673
rect 4516 28627 4545 28673
rect 4457 28570 4545 28627
rect 4457 28524 4470 28570
rect 4516 28524 4545 28570
rect 4457 28467 4545 28524
rect 4457 28421 4470 28467
rect 4516 28421 4545 28467
rect 4457 28364 4545 28421
rect 4457 28318 4470 28364
rect 4516 28318 4545 28364
rect 4457 28261 4545 28318
rect 4457 28215 4470 28261
rect 4516 28215 4545 28261
rect 4457 28158 4545 28215
rect 4457 28112 4470 28158
rect 4516 28112 4545 28158
rect 4457 28055 4545 28112
rect 4457 28009 4470 28055
rect 4516 28009 4545 28055
rect 4457 27952 4545 28009
rect 4457 27906 4470 27952
rect 4516 27906 4545 27952
rect 4457 27848 4545 27906
rect 4457 27802 4470 27848
rect 4516 27802 4545 27848
rect 4457 27789 4545 27802
rect 4685 28776 4789 28789
rect 4685 28730 4714 28776
rect 4760 28730 4789 28776
rect 4685 28673 4789 28730
rect 4685 28627 4714 28673
rect 4760 28627 4789 28673
rect 4685 28570 4789 28627
rect 4685 28524 4714 28570
rect 4760 28524 4789 28570
rect 4685 28467 4789 28524
rect 4685 28421 4714 28467
rect 4760 28421 4789 28467
rect 4685 28364 4789 28421
rect 4685 28318 4714 28364
rect 4760 28318 4789 28364
rect 4685 28261 4789 28318
rect 4685 28215 4714 28261
rect 4760 28215 4789 28261
rect 4685 28158 4789 28215
rect 4685 28112 4714 28158
rect 4760 28112 4789 28158
rect 4685 28055 4789 28112
rect 4685 28009 4714 28055
rect 4760 28009 4789 28055
rect 4685 27952 4789 28009
rect 4685 27906 4714 27952
rect 4760 27906 4789 27952
rect 4685 27848 4789 27906
rect 4685 27802 4714 27848
rect 4760 27802 4789 27848
rect 4685 27789 4789 27802
rect 4929 28776 5033 28789
rect 4929 28730 4958 28776
rect 5004 28730 5033 28776
rect 4929 28673 5033 28730
rect 4929 28627 4958 28673
rect 5004 28627 5033 28673
rect 4929 28570 5033 28627
rect 4929 28524 4958 28570
rect 5004 28524 5033 28570
rect 4929 28467 5033 28524
rect 4929 28421 4958 28467
rect 5004 28421 5033 28467
rect 4929 28364 5033 28421
rect 4929 28318 4958 28364
rect 5004 28318 5033 28364
rect 4929 28261 5033 28318
rect 4929 28215 4958 28261
rect 5004 28215 5033 28261
rect 4929 28158 5033 28215
rect 4929 28112 4958 28158
rect 5004 28112 5033 28158
rect 4929 28055 5033 28112
rect 4929 28009 4958 28055
rect 5004 28009 5033 28055
rect 4929 27952 5033 28009
rect 4929 27906 4958 27952
rect 5004 27906 5033 27952
rect 4929 27848 5033 27906
rect 4929 27802 4958 27848
rect 5004 27802 5033 27848
rect 4929 27789 5033 27802
rect 5173 28776 5277 28789
rect 5173 28730 5202 28776
rect 5248 28730 5277 28776
rect 5173 28673 5277 28730
rect 5173 28627 5202 28673
rect 5248 28627 5277 28673
rect 5173 28570 5277 28627
rect 5173 28524 5202 28570
rect 5248 28524 5277 28570
rect 5173 28467 5277 28524
rect 5173 28421 5202 28467
rect 5248 28421 5277 28467
rect 5173 28364 5277 28421
rect 5173 28318 5202 28364
rect 5248 28318 5277 28364
rect 5173 28261 5277 28318
rect 5173 28215 5202 28261
rect 5248 28215 5277 28261
rect 5173 28158 5277 28215
rect 5173 28112 5202 28158
rect 5248 28112 5277 28158
rect 5173 28055 5277 28112
rect 5173 28009 5202 28055
rect 5248 28009 5277 28055
rect 5173 27952 5277 28009
rect 5173 27906 5202 27952
rect 5248 27906 5277 27952
rect 5173 27848 5277 27906
rect 5173 27802 5202 27848
rect 5248 27802 5277 27848
rect 5173 27789 5277 27802
rect 5417 28776 5521 28789
rect 5417 28730 5446 28776
rect 5492 28730 5521 28776
rect 5417 28673 5521 28730
rect 5417 28627 5446 28673
rect 5492 28627 5521 28673
rect 5417 28570 5521 28627
rect 5417 28524 5446 28570
rect 5492 28524 5521 28570
rect 5417 28467 5521 28524
rect 5417 28421 5446 28467
rect 5492 28421 5521 28467
rect 5417 28364 5521 28421
rect 5417 28318 5446 28364
rect 5492 28318 5521 28364
rect 5417 28261 5521 28318
rect 5417 28215 5446 28261
rect 5492 28215 5521 28261
rect 5417 28158 5521 28215
rect 5417 28112 5446 28158
rect 5492 28112 5521 28158
rect 5417 28055 5521 28112
rect 5417 28009 5446 28055
rect 5492 28009 5521 28055
rect 5417 27952 5521 28009
rect 5417 27906 5446 27952
rect 5492 27906 5521 27952
rect 5417 27848 5521 27906
rect 5417 27802 5446 27848
rect 5492 27802 5521 27848
rect 5417 27789 5521 27802
rect 5661 28776 5765 28789
rect 5661 28730 5690 28776
rect 5736 28730 5765 28776
rect 5661 28673 5765 28730
rect 5661 28627 5690 28673
rect 5736 28627 5765 28673
rect 5661 28570 5765 28627
rect 5661 28524 5690 28570
rect 5736 28524 5765 28570
rect 5661 28467 5765 28524
rect 5661 28421 5690 28467
rect 5736 28421 5765 28467
rect 5661 28364 5765 28421
rect 5661 28318 5690 28364
rect 5736 28318 5765 28364
rect 5661 28261 5765 28318
rect 5661 28215 5690 28261
rect 5736 28215 5765 28261
rect 5661 28158 5765 28215
rect 5661 28112 5690 28158
rect 5736 28112 5765 28158
rect 5661 28055 5765 28112
rect 5661 28009 5690 28055
rect 5736 28009 5765 28055
rect 5661 27952 5765 28009
rect 5661 27906 5690 27952
rect 5736 27906 5765 27952
rect 5661 27848 5765 27906
rect 5661 27802 5690 27848
rect 5736 27802 5765 27848
rect 5661 27789 5765 27802
rect 5905 28776 6009 28789
rect 5905 28730 5934 28776
rect 5980 28730 6009 28776
rect 5905 28673 6009 28730
rect 5905 28627 5934 28673
rect 5980 28627 6009 28673
rect 5905 28570 6009 28627
rect 5905 28524 5934 28570
rect 5980 28524 6009 28570
rect 5905 28467 6009 28524
rect 5905 28421 5934 28467
rect 5980 28421 6009 28467
rect 5905 28364 6009 28421
rect 5905 28318 5934 28364
rect 5980 28318 6009 28364
rect 5905 28261 6009 28318
rect 5905 28215 5934 28261
rect 5980 28215 6009 28261
rect 5905 28158 6009 28215
rect 5905 28112 5934 28158
rect 5980 28112 6009 28158
rect 5905 28055 6009 28112
rect 5905 28009 5934 28055
rect 5980 28009 6009 28055
rect 5905 27952 6009 28009
rect 5905 27906 5934 27952
rect 5980 27906 6009 27952
rect 5905 27848 6009 27906
rect 5905 27802 5934 27848
rect 5980 27802 6009 27848
rect 5905 27789 6009 27802
rect 6149 28776 6253 28789
rect 6149 28730 6178 28776
rect 6224 28730 6253 28776
rect 6149 28673 6253 28730
rect 6149 28627 6178 28673
rect 6224 28627 6253 28673
rect 6149 28570 6253 28627
rect 6149 28524 6178 28570
rect 6224 28524 6253 28570
rect 6149 28467 6253 28524
rect 6149 28421 6178 28467
rect 6224 28421 6253 28467
rect 6149 28364 6253 28421
rect 6149 28318 6178 28364
rect 6224 28318 6253 28364
rect 6149 28261 6253 28318
rect 6149 28215 6178 28261
rect 6224 28215 6253 28261
rect 6149 28158 6253 28215
rect 6149 28112 6178 28158
rect 6224 28112 6253 28158
rect 6149 28055 6253 28112
rect 6149 28009 6178 28055
rect 6224 28009 6253 28055
rect 6149 27952 6253 28009
rect 6149 27906 6178 27952
rect 6224 27906 6253 27952
rect 6149 27848 6253 27906
rect 6149 27802 6178 27848
rect 6224 27802 6253 27848
rect 6149 27789 6253 27802
rect 6393 28776 6497 28789
rect 6393 28730 6422 28776
rect 6468 28730 6497 28776
rect 6393 28673 6497 28730
rect 6393 28627 6422 28673
rect 6468 28627 6497 28673
rect 6393 28570 6497 28627
rect 6393 28524 6422 28570
rect 6468 28524 6497 28570
rect 6393 28467 6497 28524
rect 6393 28421 6422 28467
rect 6468 28421 6497 28467
rect 6393 28364 6497 28421
rect 6393 28318 6422 28364
rect 6468 28318 6497 28364
rect 6393 28261 6497 28318
rect 6393 28215 6422 28261
rect 6468 28215 6497 28261
rect 6393 28158 6497 28215
rect 6393 28112 6422 28158
rect 6468 28112 6497 28158
rect 6393 28055 6497 28112
rect 6393 28009 6422 28055
rect 6468 28009 6497 28055
rect 6393 27952 6497 28009
rect 6393 27906 6422 27952
rect 6468 27906 6497 27952
rect 6393 27848 6497 27906
rect 6393 27802 6422 27848
rect 6468 27802 6497 27848
rect 6393 27789 6497 27802
rect 6637 28776 6741 28789
rect 6637 28730 6666 28776
rect 6712 28730 6741 28776
rect 6637 28673 6741 28730
rect 6637 28627 6666 28673
rect 6712 28627 6741 28673
rect 6637 28570 6741 28627
rect 6637 28524 6666 28570
rect 6712 28524 6741 28570
rect 6637 28467 6741 28524
rect 6637 28421 6666 28467
rect 6712 28421 6741 28467
rect 6637 28364 6741 28421
rect 6637 28318 6666 28364
rect 6712 28318 6741 28364
rect 6637 28261 6741 28318
rect 6637 28215 6666 28261
rect 6712 28215 6741 28261
rect 6637 28158 6741 28215
rect 6637 28112 6666 28158
rect 6712 28112 6741 28158
rect 6637 28055 6741 28112
rect 6637 28009 6666 28055
rect 6712 28009 6741 28055
rect 6637 27952 6741 28009
rect 6637 27906 6666 27952
rect 6712 27906 6741 27952
rect 6637 27848 6741 27906
rect 6637 27802 6666 27848
rect 6712 27802 6741 27848
rect 6637 27789 6741 27802
rect 6881 28776 6985 28789
rect 6881 28730 6910 28776
rect 6956 28730 6985 28776
rect 6881 28673 6985 28730
rect 6881 28627 6910 28673
rect 6956 28627 6985 28673
rect 6881 28570 6985 28627
rect 6881 28524 6910 28570
rect 6956 28524 6985 28570
rect 6881 28467 6985 28524
rect 6881 28421 6910 28467
rect 6956 28421 6985 28467
rect 6881 28364 6985 28421
rect 6881 28318 6910 28364
rect 6956 28318 6985 28364
rect 6881 28261 6985 28318
rect 6881 28215 6910 28261
rect 6956 28215 6985 28261
rect 6881 28158 6985 28215
rect 6881 28112 6910 28158
rect 6956 28112 6985 28158
rect 6881 28055 6985 28112
rect 6881 28009 6910 28055
rect 6956 28009 6985 28055
rect 6881 27952 6985 28009
rect 6881 27906 6910 27952
rect 6956 27906 6985 27952
rect 6881 27848 6985 27906
rect 6881 27802 6910 27848
rect 6956 27802 6985 27848
rect 6881 27789 6985 27802
rect 7125 28776 7229 28789
rect 7125 28730 7154 28776
rect 7200 28730 7229 28776
rect 7125 28673 7229 28730
rect 7125 28627 7154 28673
rect 7200 28627 7229 28673
rect 7125 28570 7229 28627
rect 7125 28524 7154 28570
rect 7200 28524 7229 28570
rect 7125 28467 7229 28524
rect 7125 28421 7154 28467
rect 7200 28421 7229 28467
rect 7125 28364 7229 28421
rect 7125 28318 7154 28364
rect 7200 28318 7229 28364
rect 7125 28261 7229 28318
rect 7125 28215 7154 28261
rect 7200 28215 7229 28261
rect 7125 28158 7229 28215
rect 7125 28112 7154 28158
rect 7200 28112 7229 28158
rect 7125 28055 7229 28112
rect 7125 28009 7154 28055
rect 7200 28009 7229 28055
rect 7125 27952 7229 28009
rect 7125 27906 7154 27952
rect 7200 27906 7229 27952
rect 7125 27848 7229 27906
rect 7125 27802 7154 27848
rect 7200 27802 7229 27848
rect 7125 27789 7229 27802
rect 7369 28776 7473 28789
rect 7369 28730 7398 28776
rect 7444 28730 7473 28776
rect 7369 28673 7473 28730
rect 7369 28627 7398 28673
rect 7444 28627 7473 28673
rect 7369 28570 7473 28627
rect 7369 28524 7398 28570
rect 7444 28524 7473 28570
rect 7369 28467 7473 28524
rect 7369 28421 7398 28467
rect 7444 28421 7473 28467
rect 7369 28364 7473 28421
rect 7369 28318 7398 28364
rect 7444 28318 7473 28364
rect 7369 28261 7473 28318
rect 7369 28215 7398 28261
rect 7444 28215 7473 28261
rect 7369 28158 7473 28215
rect 7369 28112 7398 28158
rect 7444 28112 7473 28158
rect 7369 28055 7473 28112
rect 7369 28009 7398 28055
rect 7444 28009 7473 28055
rect 7369 27952 7473 28009
rect 7369 27906 7398 27952
rect 7444 27906 7473 27952
rect 7369 27848 7473 27906
rect 7369 27802 7398 27848
rect 7444 27802 7473 27848
rect 7369 27789 7473 27802
rect 7613 28776 7717 28789
rect 7613 28730 7642 28776
rect 7688 28730 7717 28776
rect 7613 28673 7717 28730
rect 7613 28627 7642 28673
rect 7688 28627 7717 28673
rect 7613 28570 7717 28627
rect 7613 28524 7642 28570
rect 7688 28524 7717 28570
rect 7613 28467 7717 28524
rect 7613 28421 7642 28467
rect 7688 28421 7717 28467
rect 7613 28364 7717 28421
rect 7613 28318 7642 28364
rect 7688 28318 7717 28364
rect 7613 28261 7717 28318
rect 7613 28215 7642 28261
rect 7688 28215 7717 28261
rect 7613 28158 7717 28215
rect 7613 28112 7642 28158
rect 7688 28112 7717 28158
rect 7613 28055 7717 28112
rect 7613 28009 7642 28055
rect 7688 28009 7717 28055
rect 7613 27952 7717 28009
rect 7613 27906 7642 27952
rect 7688 27906 7717 27952
rect 7613 27848 7717 27906
rect 7613 27802 7642 27848
rect 7688 27802 7717 27848
rect 7613 27789 7717 27802
rect 7857 28776 7961 28789
rect 7857 28730 7886 28776
rect 7932 28730 7961 28776
rect 7857 28673 7961 28730
rect 7857 28627 7886 28673
rect 7932 28627 7961 28673
rect 7857 28570 7961 28627
rect 7857 28524 7886 28570
rect 7932 28524 7961 28570
rect 7857 28467 7961 28524
rect 7857 28421 7886 28467
rect 7932 28421 7961 28467
rect 7857 28364 7961 28421
rect 7857 28318 7886 28364
rect 7932 28318 7961 28364
rect 7857 28261 7961 28318
rect 7857 28215 7886 28261
rect 7932 28215 7961 28261
rect 7857 28158 7961 28215
rect 7857 28112 7886 28158
rect 7932 28112 7961 28158
rect 7857 28055 7961 28112
rect 7857 28009 7886 28055
rect 7932 28009 7961 28055
rect 7857 27952 7961 28009
rect 7857 27906 7886 27952
rect 7932 27906 7961 27952
rect 7857 27848 7961 27906
rect 7857 27802 7886 27848
rect 7932 27802 7961 27848
rect 7857 27789 7961 27802
rect 8101 28776 8205 28789
rect 8101 28730 8130 28776
rect 8176 28730 8205 28776
rect 8101 28673 8205 28730
rect 8101 28627 8130 28673
rect 8176 28627 8205 28673
rect 8101 28570 8205 28627
rect 8101 28524 8130 28570
rect 8176 28524 8205 28570
rect 8101 28467 8205 28524
rect 8101 28421 8130 28467
rect 8176 28421 8205 28467
rect 8101 28364 8205 28421
rect 8101 28318 8130 28364
rect 8176 28318 8205 28364
rect 8101 28261 8205 28318
rect 8101 28215 8130 28261
rect 8176 28215 8205 28261
rect 8101 28158 8205 28215
rect 8101 28112 8130 28158
rect 8176 28112 8205 28158
rect 8101 28055 8205 28112
rect 8101 28009 8130 28055
rect 8176 28009 8205 28055
rect 8101 27952 8205 28009
rect 8101 27906 8130 27952
rect 8176 27906 8205 27952
rect 8101 27848 8205 27906
rect 8101 27802 8130 27848
rect 8176 27802 8205 27848
rect 8101 27789 8205 27802
rect 8345 28776 8449 28789
rect 8345 28730 8374 28776
rect 8420 28730 8449 28776
rect 8345 28673 8449 28730
rect 8345 28627 8374 28673
rect 8420 28627 8449 28673
rect 8345 28570 8449 28627
rect 8345 28524 8374 28570
rect 8420 28524 8449 28570
rect 8345 28467 8449 28524
rect 8345 28421 8374 28467
rect 8420 28421 8449 28467
rect 8345 28364 8449 28421
rect 8345 28318 8374 28364
rect 8420 28318 8449 28364
rect 8345 28261 8449 28318
rect 8345 28215 8374 28261
rect 8420 28215 8449 28261
rect 8345 28158 8449 28215
rect 8345 28112 8374 28158
rect 8420 28112 8449 28158
rect 8345 28055 8449 28112
rect 8345 28009 8374 28055
rect 8420 28009 8449 28055
rect 8345 27952 8449 28009
rect 8345 27906 8374 27952
rect 8420 27906 8449 27952
rect 8345 27848 8449 27906
rect 8345 27802 8374 27848
rect 8420 27802 8449 27848
rect 8345 27789 8449 27802
rect 8589 28776 8693 28789
rect 8589 28730 8618 28776
rect 8664 28730 8693 28776
rect 8589 28673 8693 28730
rect 8589 28627 8618 28673
rect 8664 28627 8693 28673
rect 8589 28570 8693 28627
rect 8589 28524 8618 28570
rect 8664 28524 8693 28570
rect 8589 28467 8693 28524
rect 8589 28421 8618 28467
rect 8664 28421 8693 28467
rect 8589 28364 8693 28421
rect 8589 28318 8618 28364
rect 8664 28318 8693 28364
rect 8589 28261 8693 28318
rect 8589 28215 8618 28261
rect 8664 28215 8693 28261
rect 8589 28158 8693 28215
rect 8589 28112 8618 28158
rect 8664 28112 8693 28158
rect 8589 28055 8693 28112
rect 8589 28009 8618 28055
rect 8664 28009 8693 28055
rect 8589 27952 8693 28009
rect 8589 27906 8618 27952
rect 8664 27906 8693 27952
rect 8589 27848 8693 27906
rect 8589 27802 8618 27848
rect 8664 27802 8693 27848
rect 8589 27789 8693 27802
rect 8833 28776 8937 28789
rect 8833 28730 8862 28776
rect 8908 28730 8937 28776
rect 8833 28673 8937 28730
rect 8833 28627 8862 28673
rect 8908 28627 8937 28673
rect 8833 28570 8937 28627
rect 8833 28524 8862 28570
rect 8908 28524 8937 28570
rect 8833 28467 8937 28524
rect 8833 28421 8862 28467
rect 8908 28421 8937 28467
rect 8833 28364 8937 28421
rect 8833 28318 8862 28364
rect 8908 28318 8937 28364
rect 8833 28261 8937 28318
rect 8833 28215 8862 28261
rect 8908 28215 8937 28261
rect 8833 28158 8937 28215
rect 8833 28112 8862 28158
rect 8908 28112 8937 28158
rect 8833 28055 8937 28112
rect 8833 28009 8862 28055
rect 8908 28009 8937 28055
rect 8833 27952 8937 28009
rect 8833 27906 8862 27952
rect 8908 27906 8937 27952
rect 8833 27848 8937 27906
rect 8833 27802 8862 27848
rect 8908 27802 8937 27848
rect 8833 27789 8937 27802
rect 9077 28776 9181 28789
rect 9077 28730 9106 28776
rect 9152 28730 9181 28776
rect 9077 28673 9181 28730
rect 9077 28627 9106 28673
rect 9152 28627 9181 28673
rect 9077 28570 9181 28627
rect 9077 28524 9106 28570
rect 9152 28524 9181 28570
rect 9077 28467 9181 28524
rect 9077 28421 9106 28467
rect 9152 28421 9181 28467
rect 9077 28364 9181 28421
rect 9077 28318 9106 28364
rect 9152 28318 9181 28364
rect 9077 28261 9181 28318
rect 9077 28215 9106 28261
rect 9152 28215 9181 28261
rect 9077 28158 9181 28215
rect 9077 28112 9106 28158
rect 9152 28112 9181 28158
rect 9077 28055 9181 28112
rect 9077 28009 9106 28055
rect 9152 28009 9181 28055
rect 9077 27952 9181 28009
rect 9077 27906 9106 27952
rect 9152 27906 9181 27952
rect 9077 27848 9181 27906
rect 9077 27802 9106 27848
rect 9152 27802 9181 27848
rect 9077 27789 9181 27802
rect 9321 28776 9425 28789
rect 9321 28730 9350 28776
rect 9396 28730 9425 28776
rect 9321 28673 9425 28730
rect 9321 28627 9350 28673
rect 9396 28627 9425 28673
rect 9321 28570 9425 28627
rect 9321 28524 9350 28570
rect 9396 28524 9425 28570
rect 9321 28467 9425 28524
rect 9321 28421 9350 28467
rect 9396 28421 9425 28467
rect 9321 28364 9425 28421
rect 9321 28318 9350 28364
rect 9396 28318 9425 28364
rect 9321 28261 9425 28318
rect 9321 28215 9350 28261
rect 9396 28215 9425 28261
rect 9321 28158 9425 28215
rect 9321 28112 9350 28158
rect 9396 28112 9425 28158
rect 9321 28055 9425 28112
rect 9321 28009 9350 28055
rect 9396 28009 9425 28055
rect 9321 27952 9425 28009
rect 9321 27906 9350 27952
rect 9396 27906 9425 27952
rect 9321 27848 9425 27906
rect 9321 27802 9350 27848
rect 9396 27802 9425 27848
rect 9321 27789 9425 27802
rect 9565 28776 9669 28789
rect 9565 28730 9594 28776
rect 9640 28730 9669 28776
rect 9565 28673 9669 28730
rect 9565 28627 9594 28673
rect 9640 28627 9669 28673
rect 9565 28570 9669 28627
rect 9565 28524 9594 28570
rect 9640 28524 9669 28570
rect 9565 28467 9669 28524
rect 9565 28421 9594 28467
rect 9640 28421 9669 28467
rect 9565 28364 9669 28421
rect 9565 28318 9594 28364
rect 9640 28318 9669 28364
rect 9565 28261 9669 28318
rect 9565 28215 9594 28261
rect 9640 28215 9669 28261
rect 9565 28158 9669 28215
rect 9565 28112 9594 28158
rect 9640 28112 9669 28158
rect 9565 28055 9669 28112
rect 9565 28009 9594 28055
rect 9640 28009 9669 28055
rect 9565 27952 9669 28009
rect 9565 27906 9594 27952
rect 9640 27906 9669 27952
rect 9565 27848 9669 27906
rect 9565 27802 9594 27848
rect 9640 27802 9669 27848
rect 9565 27789 9669 27802
rect 9809 28776 9913 28789
rect 9809 28730 9838 28776
rect 9884 28730 9913 28776
rect 9809 28673 9913 28730
rect 9809 28627 9838 28673
rect 9884 28627 9913 28673
rect 9809 28570 9913 28627
rect 9809 28524 9838 28570
rect 9884 28524 9913 28570
rect 9809 28467 9913 28524
rect 9809 28421 9838 28467
rect 9884 28421 9913 28467
rect 9809 28364 9913 28421
rect 9809 28318 9838 28364
rect 9884 28318 9913 28364
rect 9809 28261 9913 28318
rect 9809 28215 9838 28261
rect 9884 28215 9913 28261
rect 9809 28158 9913 28215
rect 9809 28112 9838 28158
rect 9884 28112 9913 28158
rect 9809 28055 9913 28112
rect 9809 28009 9838 28055
rect 9884 28009 9913 28055
rect 9809 27952 9913 28009
rect 9809 27906 9838 27952
rect 9884 27906 9913 27952
rect 9809 27848 9913 27906
rect 9809 27802 9838 27848
rect 9884 27802 9913 27848
rect 9809 27789 9913 27802
rect 10053 28776 10157 28789
rect 10053 28730 10082 28776
rect 10128 28730 10157 28776
rect 10053 28673 10157 28730
rect 10053 28627 10082 28673
rect 10128 28627 10157 28673
rect 10053 28570 10157 28627
rect 10053 28524 10082 28570
rect 10128 28524 10157 28570
rect 10053 28467 10157 28524
rect 10053 28421 10082 28467
rect 10128 28421 10157 28467
rect 10053 28364 10157 28421
rect 10053 28318 10082 28364
rect 10128 28318 10157 28364
rect 10053 28261 10157 28318
rect 10053 28215 10082 28261
rect 10128 28215 10157 28261
rect 10053 28158 10157 28215
rect 10053 28112 10082 28158
rect 10128 28112 10157 28158
rect 10053 28055 10157 28112
rect 10053 28009 10082 28055
rect 10128 28009 10157 28055
rect 10053 27952 10157 28009
rect 10053 27906 10082 27952
rect 10128 27906 10157 27952
rect 10053 27848 10157 27906
rect 10053 27802 10082 27848
rect 10128 27802 10157 27848
rect 10053 27789 10157 27802
rect 10297 28776 10385 28789
rect 10297 28730 10326 28776
rect 10372 28730 10385 28776
rect 10297 28673 10385 28730
rect 10297 28627 10326 28673
rect 10372 28627 10385 28673
rect 10297 28570 10385 28627
rect 10297 28524 10326 28570
rect 10372 28524 10385 28570
rect 10297 28467 10385 28524
rect 10297 28421 10326 28467
rect 10372 28421 10385 28467
rect 10297 28364 10385 28421
rect 10297 28318 10326 28364
rect 10372 28318 10385 28364
rect 10297 28261 10385 28318
rect 10297 28215 10326 28261
rect 10372 28215 10385 28261
rect 10297 28158 10385 28215
rect 10297 28112 10326 28158
rect 10372 28112 10385 28158
rect 10297 28055 10385 28112
rect 10297 28009 10326 28055
rect 10372 28009 10385 28055
rect 10297 27952 10385 28009
rect 10297 27906 10326 27952
rect 10372 27906 10385 27952
rect 10297 27848 10385 27906
rect 10297 27802 10326 27848
rect 10372 27802 10385 27848
rect 10297 27789 10385 27802
<< mvndiffc >>
rect 4054 26947 4100 26993
rect 4054 26844 4100 26890
rect 4054 26741 4100 26787
rect 4054 26638 4100 26684
rect 4054 26535 4100 26581
rect 4054 26432 4100 26478
rect 4054 26329 4100 26375
rect 4054 26226 4100 26272
rect 4054 26123 4100 26169
rect 4054 26019 4100 26065
rect 4298 26947 4344 26993
rect 4298 26844 4344 26890
rect 4298 26741 4344 26787
rect 4298 26638 4344 26684
rect 4298 26535 4344 26581
rect 4298 26432 4344 26478
rect 4298 26329 4344 26375
rect 4298 26226 4344 26272
rect 4298 26123 4344 26169
rect 4298 26019 4344 26065
rect 5116 26947 5162 26993
rect 5116 26844 5162 26890
rect 5116 26741 5162 26787
rect 5116 26638 5162 26684
rect 5116 26535 5162 26581
rect 5116 26432 5162 26478
rect 5116 26329 5162 26375
rect 5116 26226 5162 26272
rect 5116 26123 5162 26169
rect 5116 26019 5162 26065
rect 5360 26947 5406 26993
rect 5360 26844 5406 26890
rect 5360 26741 5406 26787
rect 5360 26638 5406 26684
rect 5360 26535 5406 26581
rect 5360 26432 5406 26478
rect 5360 26329 5406 26375
rect 5360 26226 5406 26272
rect 5360 26123 5406 26169
rect 5360 26019 5406 26065
rect 5604 26947 5650 26993
rect 5604 26844 5650 26890
rect 5604 26741 5650 26787
rect 5604 26638 5650 26684
rect 5604 26535 5650 26581
rect 5604 26432 5650 26478
rect 5604 26329 5650 26375
rect 5604 26226 5650 26272
rect 5604 26123 5650 26169
rect 5604 26019 5650 26065
rect 5848 26947 5894 26993
rect 5848 26844 5894 26890
rect 5848 26741 5894 26787
rect 5848 26638 5894 26684
rect 5848 26535 5894 26581
rect 5848 26432 5894 26478
rect 5848 26329 5894 26375
rect 5848 26226 5894 26272
rect 5848 26123 5894 26169
rect 5848 26019 5894 26065
rect 6092 26947 6138 26993
rect 6092 26844 6138 26890
rect 6092 26741 6138 26787
rect 6092 26638 6138 26684
rect 6092 26535 6138 26581
rect 6092 26432 6138 26478
rect 6092 26329 6138 26375
rect 6092 26226 6138 26272
rect 6092 26123 6138 26169
rect 6092 26019 6138 26065
rect 6336 26947 6382 26993
rect 6336 26844 6382 26890
rect 6336 26741 6382 26787
rect 6336 26638 6382 26684
rect 6336 26535 6382 26581
rect 6336 26432 6382 26478
rect 6336 26329 6382 26375
rect 6336 26226 6382 26272
rect 6336 26123 6382 26169
rect 6336 26019 6382 26065
rect 6580 26947 6626 26993
rect 6580 26844 6626 26890
rect 6580 26741 6626 26787
rect 6580 26638 6626 26684
rect 6580 26535 6626 26581
rect 6580 26432 6626 26478
rect 6580 26329 6626 26375
rect 6580 26226 6626 26272
rect 6580 26123 6626 26169
rect 6580 26019 6626 26065
rect 6824 26947 6870 26993
rect 6824 26844 6870 26890
rect 6824 26741 6870 26787
rect 6824 26638 6870 26684
rect 6824 26535 6870 26581
rect 6824 26432 6870 26478
rect 6824 26329 6870 26375
rect 6824 26226 6870 26272
rect 6824 26123 6870 26169
rect 6824 26019 6870 26065
rect 7068 26947 7114 26993
rect 7068 26844 7114 26890
rect 7068 26741 7114 26787
rect 7068 26638 7114 26684
rect 7068 26535 7114 26581
rect 7068 26432 7114 26478
rect 7068 26329 7114 26375
rect 7068 26226 7114 26272
rect 7068 26123 7114 26169
rect 7068 26019 7114 26065
rect 7312 26947 7358 26993
rect 7312 26844 7358 26890
rect 7312 26741 7358 26787
rect 7312 26638 7358 26684
rect 7312 26535 7358 26581
rect 7312 26432 7358 26478
rect 7312 26329 7358 26375
rect 7312 26226 7358 26272
rect 7312 26123 7358 26169
rect 7312 26019 7358 26065
rect 7556 26947 7602 26993
rect 7556 26844 7602 26890
rect 7556 26741 7602 26787
rect 7556 26638 7602 26684
rect 7556 26535 7602 26581
rect 7556 26432 7602 26478
rect 7556 26329 7602 26375
rect 7556 26226 7602 26272
rect 7556 26123 7602 26169
rect 7556 26019 7602 26065
rect 7800 26947 7846 26993
rect 7800 26844 7846 26890
rect 7800 26741 7846 26787
rect 7800 26638 7846 26684
rect 7800 26535 7846 26581
rect 7800 26432 7846 26478
rect 7800 26329 7846 26375
rect 7800 26226 7846 26272
rect 7800 26123 7846 26169
rect 7800 26019 7846 26065
rect 8044 26947 8090 26993
rect 8044 26844 8090 26890
rect 8044 26741 8090 26787
rect 8044 26638 8090 26684
rect 8044 26535 8090 26581
rect 8044 26432 8090 26478
rect 8044 26329 8090 26375
rect 8044 26226 8090 26272
rect 8044 26123 8090 26169
rect 8044 26019 8090 26065
<< mvpdiffc >>
rect 2590 28730 2636 28776
rect 2590 28627 2636 28673
rect 2590 28524 2636 28570
rect 2590 28421 2636 28467
rect 2590 28318 2636 28364
rect 2590 28215 2636 28261
rect 2590 28112 2636 28158
rect 2590 28009 2636 28055
rect 2590 27906 2636 27952
rect 2590 27802 2636 27848
rect 2834 28730 2880 28776
rect 2834 28627 2880 28673
rect 2834 28524 2880 28570
rect 2834 28421 2880 28467
rect 2834 28318 2880 28364
rect 2834 28215 2880 28261
rect 2834 28112 2880 28158
rect 2834 28009 2880 28055
rect 2834 27906 2880 27952
rect 2834 27802 2880 27848
rect 3078 28730 3124 28776
rect 3078 28627 3124 28673
rect 3078 28524 3124 28570
rect 3078 28421 3124 28467
rect 3078 28318 3124 28364
rect 3078 28215 3124 28261
rect 3078 28112 3124 28158
rect 3078 28009 3124 28055
rect 3078 27906 3124 27952
rect 3078 27802 3124 27848
rect 3322 28730 3368 28776
rect 3322 28627 3368 28673
rect 3322 28524 3368 28570
rect 3322 28421 3368 28467
rect 3322 28318 3368 28364
rect 3322 28215 3368 28261
rect 3322 28112 3368 28158
rect 3322 28009 3368 28055
rect 3322 27906 3368 27952
rect 3322 27802 3368 27848
rect 3566 28730 3612 28776
rect 3566 28627 3612 28673
rect 3566 28524 3612 28570
rect 3566 28421 3612 28467
rect 3566 28318 3612 28364
rect 3566 28215 3612 28261
rect 3566 28112 3612 28158
rect 3566 28009 3612 28055
rect 3566 27906 3612 27952
rect 3566 27802 3612 27848
rect 3810 28730 3856 28776
rect 3810 28627 3856 28673
rect 3810 28524 3856 28570
rect 3810 28421 3856 28467
rect 3810 28318 3856 28364
rect 3810 28215 3856 28261
rect 3810 28112 3856 28158
rect 3810 28009 3856 28055
rect 3810 27906 3856 27952
rect 3810 27802 3856 27848
rect 4054 28730 4100 28776
rect 4054 28627 4100 28673
rect 4054 28524 4100 28570
rect 4054 28421 4100 28467
rect 4054 28318 4100 28364
rect 4054 28215 4100 28261
rect 4054 28112 4100 28158
rect 4054 28009 4100 28055
rect 4054 27906 4100 27952
rect 4054 27802 4100 27848
rect 4298 28730 4344 28776
rect 4298 28627 4344 28673
rect 4298 28524 4344 28570
rect 4298 28421 4344 28467
rect 4298 28318 4344 28364
rect 4298 28215 4344 28261
rect 4298 28112 4344 28158
rect 4298 28009 4344 28055
rect 4298 27906 4344 27952
rect 4298 27802 4344 27848
rect 4470 28730 4516 28776
rect 4470 28627 4516 28673
rect 4470 28524 4516 28570
rect 4470 28421 4516 28467
rect 4470 28318 4516 28364
rect 4470 28215 4516 28261
rect 4470 28112 4516 28158
rect 4470 28009 4516 28055
rect 4470 27906 4516 27952
rect 4470 27802 4516 27848
rect 4714 28730 4760 28776
rect 4714 28627 4760 28673
rect 4714 28524 4760 28570
rect 4714 28421 4760 28467
rect 4714 28318 4760 28364
rect 4714 28215 4760 28261
rect 4714 28112 4760 28158
rect 4714 28009 4760 28055
rect 4714 27906 4760 27952
rect 4714 27802 4760 27848
rect 4958 28730 5004 28776
rect 4958 28627 5004 28673
rect 4958 28524 5004 28570
rect 4958 28421 5004 28467
rect 4958 28318 5004 28364
rect 4958 28215 5004 28261
rect 4958 28112 5004 28158
rect 4958 28009 5004 28055
rect 4958 27906 5004 27952
rect 4958 27802 5004 27848
rect 5202 28730 5248 28776
rect 5202 28627 5248 28673
rect 5202 28524 5248 28570
rect 5202 28421 5248 28467
rect 5202 28318 5248 28364
rect 5202 28215 5248 28261
rect 5202 28112 5248 28158
rect 5202 28009 5248 28055
rect 5202 27906 5248 27952
rect 5202 27802 5248 27848
rect 5446 28730 5492 28776
rect 5446 28627 5492 28673
rect 5446 28524 5492 28570
rect 5446 28421 5492 28467
rect 5446 28318 5492 28364
rect 5446 28215 5492 28261
rect 5446 28112 5492 28158
rect 5446 28009 5492 28055
rect 5446 27906 5492 27952
rect 5446 27802 5492 27848
rect 5690 28730 5736 28776
rect 5690 28627 5736 28673
rect 5690 28524 5736 28570
rect 5690 28421 5736 28467
rect 5690 28318 5736 28364
rect 5690 28215 5736 28261
rect 5690 28112 5736 28158
rect 5690 28009 5736 28055
rect 5690 27906 5736 27952
rect 5690 27802 5736 27848
rect 5934 28730 5980 28776
rect 5934 28627 5980 28673
rect 5934 28524 5980 28570
rect 5934 28421 5980 28467
rect 5934 28318 5980 28364
rect 5934 28215 5980 28261
rect 5934 28112 5980 28158
rect 5934 28009 5980 28055
rect 5934 27906 5980 27952
rect 5934 27802 5980 27848
rect 6178 28730 6224 28776
rect 6178 28627 6224 28673
rect 6178 28524 6224 28570
rect 6178 28421 6224 28467
rect 6178 28318 6224 28364
rect 6178 28215 6224 28261
rect 6178 28112 6224 28158
rect 6178 28009 6224 28055
rect 6178 27906 6224 27952
rect 6178 27802 6224 27848
rect 6422 28730 6468 28776
rect 6422 28627 6468 28673
rect 6422 28524 6468 28570
rect 6422 28421 6468 28467
rect 6422 28318 6468 28364
rect 6422 28215 6468 28261
rect 6422 28112 6468 28158
rect 6422 28009 6468 28055
rect 6422 27906 6468 27952
rect 6422 27802 6468 27848
rect 6666 28730 6712 28776
rect 6666 28627 6712 28673
rect 6666 28524 6712 28570
rect 6666 28421 6712 28467
rect 6666 28318 6712 28364
rect 6666 28215 6712 28261
rect 6666 28112 6712 28158
rect 6666 28009 6712 28055
rect 6666 27906 6712 27952
rect 6666 27802 6712 27848
rect 6910 28730 6956 28776
rect 6910 28627 6956 28673
rect 6910 28524 6956 28570
rect 6910 28421 6956 28467
rect 6910 28318 6956 28364
rect 6910 28215 6956 28261
rect 6910 28112 6956 28158
rect 6910 28009 6956 28055
rect 6910 27906 6956 27952
rect 6910 27802 6956 27848
rect 7154 28730 7200 28776
rect 7154 28627 7200 28673
rect 7154 28524 7200 28570
rect 7154 28421 7200 28467
rect 7154 28318 7200 28364
rect 7154 28215 7200 28261
rect 7154 28112 7200 28158
rect 7154 28009 7200 28055
rect 7154 27906 7200 27952
rect 7154 27802 7200 27848
rect 7398 28730 7444 28776
rect 7398 28627 7444 28673
rect 7398 28524 7444 28570
rect 7398 28421 7444 28467
rect 7398 28318 7444 28364
rect 7398 28215 7444 28261
rect 7398 28112 7444 28158
rect 7398 28009 7444 28055
rect 7398 27906 7444 27952
rect 7398 27802 7444 27848
rect 7642 28730 7688 28776
rect 7642 28627 7688 28673
rect 7642 28524 7688 28570
rect 7642 28421 7688 28467
rect 7642 28318 7688 28364
rect 7642 28215 7688 28261
rect 7642 28112 7688 28158
rect 7642 28009 7688 28055
rect 7642 27906 7688 27952
rect 7642 27802 7688 27848
rect 7886 28730 7932 28776
rect 7886 28627 7932 28673
rect 7886 28524 7932 28570
rect 7886 28421 7932 28467
rect 7886 28318 7932 28364
rect 7886 28215 7932 28261
rect 7886 28112 7932 28158
rect 7886 28009 7932 28055
rect 7886 27906 7932 27952
rect 7886 27802 7932 27848
rect 8130 28730 8176 28776
rect 8130 28627 8176 28673
rect 8130 28524 8176 28570
rect 8130 28421 8176 28467
rect 8130 28318 8176 28364
rect 8130 28215 8176 28261
rect 8130 28112 8176 28158
rect 8130 28009 8176 28055
rect 8130 27906 8176 27952
rect 8130 27802 8176 27848
rect 8374 28730 8420 28776
rect 8374 28627 8420 28673
rect 8374 28524 8420 28570
rect 8374 28421 8420 28467
rect 8374 28318 8420 28364
rect 8374 28215 8420 28261
rect 8374 28112 8420 28158
rect 8374 28009 8420 28055
rect 8374 27906 8420 27952
rect 8374 27802 8420 27848
rect 8618 28730 8664 28776
rect 8618 28627 8664 28673
rect 8618 28524 8664 28570
rect 8618 28421 8664 28467
rect 8618 28318 8664 28364
rect 8618 28215 8664 28261
rect 8618 28112 8664 28158
rect 8618 28009 8664 28055
rect 8618 27906 8664 27952
rect 8618 27802 8664 27848
rect 8862 28730 8908 28776
rect 8862 28627 8908 28673
rect 8862 28524 8908 28570
rect 8862 28421 8908 28467
rect 8862 28318 8908 28364
rect 8862 28215 8908 28261
rect 8862 28112 8908 28158
rect 8862 28009 8908 28055
rect 8862 27906 8908 27952
rect 8862 27802 8908 27848
rect 9106 28730 9152 28776
rect 9106 28627 9152 28673
rect 9106 28524 9152 28570
rect 9106 28421 9152 28467
rect 9106 28318 9152 28364
rect 9106 28215 9152 28261
rect 9106 28112 9152 28158
rect 9106 28009 9152 28055
rect 9106 27906 9152 27952
rect 9106 27802 9152 27848
rect 9350 28730 9396 28776
rect 9350 28627 9396 28673
rect 9350 28524 9396 28570
rect 9350 28421 9396 28467
rect 9350 28318 9396 28364
rect 9350 28215 9396 28261
rect 9350 28112 9396 28158
rect 9350 28009 9396 28055
rect 9350 27906 9396 27952
rect 9350 27802 9396 27848
rect 9594 28730 9640 28776
rect 9594 28627 9640 28673
rect 9594 28524 9640 28570
rect 9594 28421 9640 28467
rect 9594 28318 9640 28364
rect 9594 28215 9640 28261
rect 9594 28112 9640 28158
rect 9594 28009 9640 28055
rect 9594 27906 9640 27952
rect 9594 27802 9640 27848
rect 9838 28730 9884 28776
rect 9838 28627 9884 28673
rect 9838 28524 9884 28570
rect 9838 28421 9884 28467
rect 9838 28318 9884 28364
rect 9838 28215 9884 28261
rect 9838 28112 9884 28158
rect 9838 28009 9884 28055
rect 9838 27906 9884 27952
rect 9838 27802 9884 27848
rect 10082 28730 10128 28776
rect 10082 28627 10128 28673
rect 10082 28524 10128 28570
rect 10082 28421 10128 28467
rect 10082 28318 10128 28364
rect 10082 28215 10128 28261
rect 10082 28112 10128 28158
rect 10082 28009 10128 28055
rect 10082 27906 10128 27952
rect 10082 27802 10128 27848
rect 10326 28730 10372 28776
rect 10326 28627 10372 28673
rect 10326 28524 10372 28570
rect 10326 28421 10372 28467
rect 10326 28318 10372 28364
rect 10326 28215 10372 28261
rect 10326 28112 10372 28158
rect 10326 28009 10372 28055
rect 10326 27906 10372 27952
rect 10326 27802 10372 27848
<< psubdiff >>
rect 2253 27156 2343 27178
rect 2253 25888 2275 27156
rect 2321 25888 2343 27156
rect 10619 27156 10709 27178
rect 2253 25802 2343 25888
rect 10619 25888 10641 27156
rect 10687 25888 10709 27156
rect 10619 25802 10709 25888
rect 2253 25780 10709 25802
rect 2253 25734 2275 25780
rect 6739 25734 6975 25780
rect 7209 25734 7445 25780
rect 7679 25734 8009 25780
rect 10687 25734 10709 25780
rect 2253 25712 10709 25734
<< nsubdiff >>
rect 2253 29060 10709 29082
rect 2253 29014 2275 29060
rect 10687 29014 10709 29060
rect 2253 28992 10709 29014
rect 2253 28906 2343 28992
rect 2253 27732 2275 28906
rect 2321 27732 2343 28906
rect 10619 28906 10709 28992
rect 2253 27710 2343 27732
rect 10619 27732 10641 28906
rect 10687 27732 10709 28906
rect 10619 27710 10709 27732
<< psubdiffcont >>
rect 2275 25888 2321 27156
rect 10641 25888 10687 27156
rect 2275 25734 6739 25780
rect 6975 25734 7209 25780
rect 7445 25734 7679 25780
rect 8009 25734 10687 25780
<< nsubdiffcont >>
rect 2275 29014 10687 29060
rect 2275 27732 2321 28906
rect 10641 27732 10687 28906
<< polysilicon >>
rect 2665 28789 2805 28833
rect 2909 28789 3049 28833
rect 3153 28789 3293 28833
rect 3397 28789 3537 28833
rect 3641 28789 3781 28833
rect 3885 28789 4025 28833
rect 4129 28789 4269 28833
rect 4545 28789 4685 28833
rect 4789 28789 4929 28833
rect 5033 28789 5173 28833
rect 5277 28789 5417 28833
rect 5521 28789 5661 28833
rect 5765 28789 5905 28833
rect 6009 28789 6149 28833
rect 6253 28789 6393 28833
rect 6497 28789 6637 28833
rect 6741 28789 6881 28833
rect 6985 28789 7125 28833
rect 7229 28789 7369 28833
rect 7473 28789 7613 28833
rect 7717 28789 7857 28833
rect 7961 28789 8101 28833
rect 8205 28789 8345 28833
rect 8449 28789 8589 28833
rect 8693 28789 8833 28833
rect 8937 28789 9077 28833
rect 9181 28789 9321 28833
rect 9425 28789 9565 28833
rect 9669 28789 9809 28833
rect 9913 28789 10053 28833
rect 10157 28789 10297 28833
rect 2665 27601 2805 27789
rect 2909 27601 3049 27789
rect 3153 27601 3293 27789
rect 3397 27601 3537 27789
rect 2665 27582 3537 27601
rect 2665 27536 2749 27582
rect 3453 27536 3537 27582
rect 2665 27517 3537 27536
rect 3641 27601 3781 27789
rect 3885 27601 4025 27789
rect 4129 27601 4269 27789
rect 3641 27582 4269 27601
rect 3641 27536 3697 27582
rect 4213 27536 4269 27582
rect 3641 27517 4269 27536
rect 4545 27601 4685 27789
rect 4789 27601 4929 27789
rect 5033 27601 5173 27789
rect 5277 27601 5417 27789
rect 5521 27601 5661 27789
rect 5765 27601 5905 27789
rect 6009 27601 6149 27789
rect 6253 27601 6393 27789
rect 6497 27601 6637 27789
rect 6741 27601 6881 27789
rect 6985 27601 7125 27789
rect 7229 27601 7369 27789
rect 7473 27601 7613 27789
rect 7717 27601 7857 27789
rect 7961 27601 8101 27789
rect 8205 27601 8345 27789
rect 8449 27601 8589 27789
rect 8693 27601 8833 27789
rect 8937 27601 9077 27789
rect 9181 27601 9321 27789
rect 9425 27601 9565 27789
rect 9669 27601 9809 27789
rect 9913 27601 10053 27789
rect 10157 27601 10297 27789
rect 4545 27582 10297 27601
rect 4545 27536 4578 27582
rect 10264 27536 10297 27582
rect 4545 27517 10297 27536
rect 5191 27259 6551 27278
rect 5191 27213 5237 27259
rect 6505 27213 6551 27259
rect 5191 27194 6551 27213
rect 4053 27131 4269 27150
rect 4053 27085 4072 27131
rect 4212 27085 4269 27131
rect 4053 27066 4269 27085
rect 4129 27006 4269 27066
rect 5191 27006 5331 27194
rect 5435 27006 5575 27194
rect 5679 27006 5819 27194
rect 5923 27006 6063 27194
rect 6167 27006 6307 27194
rect 6411 27006 6551 27194
rect 6655 27259 8015 27278
rect 6655 27213 6701 27259
rect 7969 27213 8015 27259
rect 6655 27194 8015 27213
rect 6655 27006 6795 27194
rect 6899 27006 7039 27194
rect 7143 27006 7283 27194
rect 7387 27006 7527 27194
rect 7631 27006 7771 27194
rect 7875 27006 8015 27194
rect 4129 25962 4269 26006
rect 5191 25962 5331 26006
rect 5435 25962 5575 26006
rect 5679 25962 5819 26006
rect 5923 25962 6063 26006
rect 6167 25962 6307 26006
rect 6411 25962 6551 26006
rect 6655 25962 6795 26006
rect 6899 25962 7039 26006
rect 7143 25962 7283 26006
rect 7387 25962 7527 26006
rect 7631 25962 7771 26006
rect 7875 25962 8015 26006
<< polycontact >>
rect 2749 27536 3453 27582
rect 3697 27536 4213 27582
rect 4578 27536 10264 27582
rect 5237 27213 6505 27259
rect 4072 27085 4212 27131
rect 6701 27213 7969 27259
<< metal1 >>
rect -1 27593 67 30038
rect 2264 29060 10698 29071
rect 2264 29014 2275 29060
rect 10687 29014 10698 29060
rect 2264 29003 10698 29014
rect 2264 28906 2332 29003
rect 2264 27732 2275 28906
rect 2321 27732 2332 28906
rect 2575 28776 2651 29003
rect 2575 28730 2590 28776
rect 2636 28730 2651 28776
rect 2575 28673 2651 28730
rect 2575 28627 2590 28673
rect 2636 28627 2651 28673
rect 2575 28570 2651 28627
rect 2575 28524 2590 28570
rect 2636 28524 2651 28570
rect 2575 28467 2651 28524
rect 2575 28421 2590 28467
rect 2636 28421 2651 28467
rect 2575 28364 2651 28421
rect 2575 28318 2590 28364
rect 2636 28318 2651 28364
rect 2575 28261 2651 28318
rect 2575 28215 2590 28261
rect 2636 28215 2651 28261
rect 2575 28158 2651 28215
rect 2575 28112 2590 28158
rect 2636 28112 2651 28158
rect 2575 28055 2651 28112
rect 2575 28009 2590 28055
rect 2636 28009 2651 28055
rect 2575 27952 2651 28009
rect 2575 27906 2590 27952
rect 2636 27906 2651 27952
rect 2575 27848 2651 27906
rect 2575 27802 2590 27848
rect 2636 27802 2651 27848
rect 2575 27789 2651 27802
rect 2819 28776 2895 28789
rect 2819 28730 2834 28776
rect 2880 28730 2895 28776
rect 2819 28673 2895 28730
rect 2819 28627 2834 28673
rect 2880 28627 2895 28673
rect 2819 28570 2895 28627
rect 2819 28524 2834 28570
rect 2880 28524 2895 28570
rect 2819 28467 2895 28524
rect 2819 28421 2834 28467
rect 2880 28421 2895 28467
rect 2819 28364 2895 28421
rect 2819 28318 2834 28364
rect 2880 28318 2895 28364
rect 2819 28261 2895 28318
rect 2819 28215 2834 28261
rect 2880 28215 2895 28261
rect 2819 28158 2895 28215
rect 2819 28112 2834 28158
rect 2880 28112 2895 28158
rect 2819 28055 2895 28112
rect 2819 28009 2834 28055
rect 2880 28009 2895 28055
rect 2819 27952 2895 28009
rect 2819 27906 2834 27952
rect 2880 27906 2895 27952
rect 2819 27848 2895 27906
rect 2819 27802 2834 27848
rect 2880 27802 2895 27848
rect 2264 27721 2332 27732
rect 2819 27729 2895 27802
rect 3063 28776 3139 29003
rect 3063 28730 3078 28776
rect 3124 28730 3139 28776
rect 3063 28673 3139 28730
rect 3063 28627 3078 28673
rect 3124 28627 3139 28673
rect 3063 28570 3139 28627
rect 3063 28524 3078 28570
rect 3124 28524 3139 28570
rect 3063 28467 3139 28524
rect 3063 28421 3078 28467
rect 3124 28421 3139 28467
rect 3063 28364 3139 28421
rect 3063 28318 3078 28364
rect 3124 28318 3139 28364
rect 3063 28261 3139 28318
rect 3063 28215 3078 28261
rect 3124 28215 3139 28261
rect 3063 28158 3139 28215
rect 3063 28112 3078 28158
rect 3124 28112 3139 28158
rect 3063 28055 3139 28112
rect 3063 28009 3078 28055
rect 3124 28009 3139 28055
rect 3063 27952 3139 28009
rect 3063 27906 3078 27952
rect 3124 27906 3139 27952
rect 3063 27848 3139 27906
rect 3063 27802 3078 27848
rect 3124 27802 3139 27848
rect 3063 27789 3139 27802
rect 3307 28776 3383 28789
rect 3307 28730 3322 28776
rect 3368 28730 3383 28776
rect 3307 28673 3383 28730
rect 3307 28627 3322 28673
rect 3368 28627 3383 28673
rect 3307 28570 3383 28627
rect 3307 28524 3322 28570
rect 3368 28524 3383 28570
rect 3307 28467 3383 28524
rect 3307 28421 3322 28467
rect 3368 28421 3383 28467
rect 3307 28364 3383 28421
rect 3307 28318 3322 28364
rect 3368 28318 3383 28364
rect 3307 28261 3383 28318
rect 3307 28215 3322 28261
rect 3368 28215 3383 28261
rect 3307 28158 3383 28215
rect 3307 28112 3322 28158
rect 3368 28112 3383 28158
rect 3307 28055 3383 28112
rect 3307 28009 3322 28055
rect 3368 28009 3383 28055
rect 3307 27952 3383 28009
rect 3307 27906 3322 27952
rect 3368 27906 3383 27952
rect 3307 27848 3383 27906
rect 3307 27802 3322 27848
rect 3368 27802 3383 27848
rect 3307 27729 3383 27802
rect 3551 28776 3627 29003
rect 3551 28730 3566 28776
rect 3612 28730 3627 28776
rect 3551 28673 3627 28730
rect 3551 28627 3566 28673
rect 3612 28627 3627 28673
rect 3551 28570 3627 28627
rect 3551 28524 3566 28570
rect 3612 28524 3627 28570
rect 3551 28467 3627 28524
rect 3551 28421 3566 28467
rect 3612 28421 3627 28467
rect 3551 28364 3627 28421
rect 3551 28318 3566 28364
rect 3612 28318 3627 28364
rect 3551 28261 3627 28318
rect 3551 28215 3566 28261
rect 3612 28215 3627 28261
rect 3551 28158 3627 28215
rect 3551 28112 3566 28158
rect 3612 28112 3627 28158
rect 3551 28055 3627 28112
rect 3551 28009 3566 28055
rect 3612 28009 3627 28055
rect 3551 27952 3627 28009
rect 3551 27906 3566 27952
rect 3612 27906 3627 27952
rect 3551 27848 3627 27906
rect 3551 27802 3566 27848
rect 3612 27802 3627 27848
rect 3551 27789 3627 27802
rect 3795 28776 3871 28789
rect 3795 28730 3810 28776
rect 3856 28730 3871 28776
rect 3795 28673 3871 28730
rect 3795 28627 3810 28673
rect 3856 28627 3871 28673
rect 3795 28570 3871 28627
rect 3795 28524 3810 28570
rect 3856 28524 3871 28570
rect 3795 28467 3871 28524
rect 3795 28421 3810 28467
rect 3856 28421 3871 28467
rect 3795 28364 3871 28421
rect 3795 28318 3810 28364
rect 3856 28318 3871 28364
rect 3795 28261 3871 28318
rect 3795 28215 3810 28261
rect 3856 28215 3871 28261
rect 3795 28158 3871 28215
rect 3795 28112 3810 28158
rect 3856 28112 3871 28158
rect 3795 28055 3871 28112
rect 3795 28009 3810 28055
rect 3856 28009 3871 28055
rect 3795 27952 3871 28009
rect 3795 27906 3810 27952
rect 3856 27906 3871 27952
rect 3795 27848 3871 27906
rect 3795 27802 3810 27848
rect 3856 27802 3871 27848
rect 3795 27729 3871 27802
rect 4039 28776 4115 29003
rect 4039 28730 4054 28776
rect 4100 28730 4115 28776
rect 4039 28673 4115 28730
rect 4039 28627 4054 28673
rect 4100 28627 4115 28673
rect 4039 28570 4115 28627
rect 4039 28524 4054 28570
rect 4100 28524 4115 28570
rect 4039 28467 4115 28524
rect 4039 28421 4054 28467
rect 4100 28421 4115 28467
rect 4039 28364 4115 28421
rect 4039 28318 4054 28364
rect 4100 28318 4115 28364
rect 4039 28261 4115 28318
rect 4039 28215 4054 28261
rect 4100 28215 4115 28261
rect 4039 28158 4115 28215
rect 4039 28112 4054 28158
rect 4100 28112 4115 28158
rect 4039 28055 4115 28112
rect 4039 28009 4054 28055
rect 4100 28009 4115 28055
rect 4039 27952 4115 28009
rect 4039 27906 4054 27952
rect 4100 27906 4115 27952
rect 4039 27848 4115 27906
rect 4039 27802 4054 27848
rect 4100 27802 4115 27848
rect 4039 27789 4115 27802
rect 4283 28776 4359 28789
rect 4283 28730 4298 28776
rect 4344 28730 4359 28776
rect 4283 28673 4359 28730
rect 4283 28627 4298 28673
rect 4344 28627 4359 28673
rect 4283 28570 4359 28627
rect 4283 28524 4298 28570
rect 4344 28524 4359 28570
rect 4283 28467 4359 28524
rect 4283 28421 4298 28467
rect 4344 28421 4359 28467
rect 4283 28364 4359 28421
rect 4283 28318 4298 28364
rect 4344 28318 4359 28364
rect 4283 28261 4359 28318
rect 4283 28215 4298 28261
rect 4344 28215 4359 28261
rect 4283 28158 4359 28215
rect 4283 28112 4298 28158
rect 4344 28112 4359 28158
rect 4283 28055 4359 28112
rect 4283 28009 4298 28055
rect 4344 28009 4359 28055
rect 4283 27952 4359 28009
rect 4283 27906 4298 27952
rect 4344 27906 4359 27952
rect 4283 27848 4359 27906
rect 4283 27802 4298 27848
rect 4344 27802 4359 27848
rect 4283 27729 4359 27802
rect 4455 28776 4531 29003
rect 4455 28730 4470 28776
rect 4516 28730 4531 28776
rect 4455 28673 4531 28730
rect 4455 28627 4470 28673
rect 4516 28627 4531 28673
rect 4455 28570 4531 28627
rect 4455 28524 4470 28570
rect 4516 28524 4531 28570
rect 4455 28467 4531 28524
rect 4455 28421 4470 28467
rect 4516 28421 4531 28467
rect 4455 28364 4531 28421
rect 4455 28318 4470 28364
rect 4516 28318 4531 28364
rect 4455 28261 4531 28318
rect 4455 28215 4470 28261
rect 4516 28215 4531 28261
rect 4455 28158 4531 28215
rect 4455 28112 4470 28158
rect 4516 28112 4531 28158
rect 4455 28055 4531 28112
rect 4455 28009 4470 28055
rect 4516 28009 4531 28055
rect 4455 27952 4531 28009
rect 4455 27906 4470 27952
rect 4516 27906 4531 27952
rect 4455 27848 4531 27906
rect 4455 27802 4470 27848
rect 4516 27802 4531 27848
rect 4455 27789 4531 27802
rect 4699 28776 4775 28789
rect 4699 28730 4714 28776
rect 4760 28730 4775 28776
rect 4699 28673 4775 28730
rect 4699 28627 4714 28673
rect 4760 28627 4775 28673
rect 4699 28570 4775 28627
rect 4699 28524 4714 28570
rect 4760 28524 4775 28570
rect 4699 28467 4775 28524
rect 4699 28421 4714 28467
rect 4760 28421 4775 28467
rect 4699 28364 4775 28421
rect 4699 28318 4714 28364
rect 4760 28318 4775 28364
rect 4699 28261 4775 28318
rect 4699 28215 4714 28261
rect 4760 28215 4775 28261
rect 4699 28158 4775 28215
rect 4699 28112 4714 28158
rect 4760 28112 4775 28158
rect 4699 28055 4775 28112
rect 4699 28009 4714 28055
rect 4760 28009 4775 28055
rect 4699 27952 4775 28009
rect 4699 27906 4714 27952
rect 4760 27906 4775 27952
rect 4699 27848 4775 27906
rect 4699 27802 4714 27848
rect 4760 27802 4775 27848
rect 2819 27653 3627 27729
rect 3795 27653 4359 27729
rect 4699 27729 4775 27802
rect 4943 28776 5019 29003
rect 4943 28730 4958 28776
rect 5004 28730 5019 28776
rect 4943 28673 5019 28730
rect 4943 28627 4958 28673
rect 5004 28627 5019 28673
rect 4943 28570 5019 28627
rect 4943 28524 4958 28570
rect 5004 28524 5019 28570
rect 4943 28467 5019 28524
rect 4943 28421 4958 28467
rect 5004 28421 5019 28467
rect 4943 28364 5019 28421
rect 4943 28318 4958 28364
rect 5004 28318 5019 28364
rect 4943 28261 5019 28318
rect 4943 28215 4958 28261
rect 5004 28215 5019 28261
rect 4943 28158 5019 28215
rect 4943 28112 4958 28158
rect 5004 28112 5019 28158
rect 4943 28055 5019 28112
rect 4943 28009 4958 28055
rect 5004 28009 5019 28055
rect 4943 27952 5019 28009
rect 4943 27906 4958 27952
rect 5004 27906 5019 27952
rect 4943 27848 5019 27906
rect 4943 27802 4958 27848
rect 5004 27802 5019 27848
rect 4943 27789 5019 27802
rect 5187 28776 5263 28789
rect 5187 28730 5202 28776
rect 5248 28730 5263 28776
rect 5187 28673 5263 28730
rect 5187 28627 5202 28673
rect 5248 28627 5263 28673
rect 5187 28570 5263 28627
rect 5187 28524 5202 28570
rect 5248 28524 5263 28570
rect 5187 28467 5263 28524
rect 5187 28421 5202 28467
rect 5248 28421 5263 28467
rect 5187 28364 5263 28421
rect 5187 28318 5202 28364
rect 5248 28318 5263 28364
rect 5187 28261 5263 28318
rect 5187 28215 5202 28261
rect 5248 28215 5263 28261
rect 5187 28158 5263 28215
rect 5187 28112 5202 28158
rect 5248 28112 5263 28158
rect 5187 28055 5263 28112
rect 5187 28009 5202 28055
rect 5248 28009 5263 28055
rect 5187 27952 5263 28009
rect 5187 27906 5202 27952
rect 5248 27906 5263 27952
rect 5187 27848 5263 27906
rect 5187 27802 5202 27848
rect 5248 27802 5263 27848
rect 5187 27729 5263 27802
rect 5431 28776 5507 29003
rect 5431 28730 5446 28776
rect 5492 28730 5507 28776
rect 5431 28673 5507 28730
rect 5431 28627 5446 28673
rect 5492 28627 5507 28673
rect 5431 28570 5507 28627
rect 5431 28524 5446 28570
rect 5492 28524 5507 28570
rect 5431 28467 5507 28524
rect 5431 28421 5446 28467
rect 5492 28421 5507 28467
rect 5431 28364 5507 28421
rect 5431 28318 5446 28364
rect 5492 28318 5507 28364
rect 5431 28261 5507 28318
rect 5431 28215 5446 28261
rect 5492 28215 5507 28261
rect 5431 28158 5507 28215
rect 5431 28112 5446 28158
rect 5492 28112 5507 28158
rect 5431 28055 5507 28112
rect 5431 28009 5446 28055
rect 5492 28009 5507 28055
rect 5431 27952 5507 28009
rect 5431 27906 5446 27952
rect 5492 27906 5507 27952
rect 5431 27848 5507 27906
rect 5431 27802 5446 27848
rect 5492 27802 5507 27848
rect 5431 27789 5507 27802
rect 5675 28776 5751 28789
rect 5675 28730 5690 28776
rect 5736 28730 5751 28776
rect 5675 28673 5751 28730
rect 5675 28627 5690 28673
rect 5736 28627 5751 28673
rect 5675 28570 5751 28627
rect 5675 28524 5690 28570
rect 5736 28524 5751 28570
rect 5675 28467 5751 28524
rect 5675 28421 5690 28467
rect 5736 28421 5751 28467
rect 5675 28364 5751 28421
rect 5675 28318 5690 28364
rect 5736 28318 5751 28364
rect 5675 28261 5751 28318
rect 5675 28215 5690 28261
rect 5736 28215 5751 28261
rect 5675 28158 5751 28215
rect 5675 28112 5690 28158
rect 5736 28112 5751 28158
rect 5675 28055 5751 28112
rect 5675 28009 5690 28055
rect 5736 28009 5751 28055
rect 5675 27952 5751 28009
rect 5675 27906 5690 27952
rect 5736 27906 5751 27952
rect 5675 27848 5751 27906
rect 5675 27802 5690 27848
rect 5736 27802 5751 27848
rect 5675 27729 5751 27802
rect 5919 28776 5995 29003
rect 5919 28730 5934 28776
rect 5980 28730 5995 28776
rect 5919 28673 5995 28730
rect 5919 28627 5934 28673
rect 5980 28627 5995 28673
rect 5919 28570 5995 28627
rect 5919 28524 5934 28570
rect 5980 28524 5995 28570
rect 5919 28467 5995 28524
rect 5919 28421 5934 28467
rect 5980 28421 5995 28467
rect 5919 28364 5995 28421
rect 5919 28318 5934 28364
rect 5980 28318 5995 28364
rect 5919 28261 5995 28318
rect 5919 28215 5934 28261
rect 5980 28215 5995 28261
rect 5919 28158 5995 28215
rect 5919 28112 5934 28158
rect 5980 28112 5995 28158
rect 5919 28055 5995 28112
rect 5919 28009 5934 28055
rect 5980 28009 5995 28055
rect 5919 27952 5995 28009
rect 5919 27906 5934 27952
rect 5980 27906 5995 27952
rect 5919 27848 5995 27906
rect 5919 27802 5934 27848
rect 5980 27802 5995 27848
rect 5919 27789 5995 27802
rect 6163 28776 6239 28789
rect 6163 28730 6178 28776
rect 6224 28730 6239 28776
rect 6163 28673 6239 28730
rect 6163 28627 6178 28673
rect 6224 28627 6239 28673
rect 6163 28570 6239 28627
rect 6163 28524 6178 28570
rect 6224 28524 6239 28570
rect 6163 28467 6239 28524
rect 6163 28421 6178 28467
rect 6224 28421 6239 28467
rect 6163 28364 6239 28421
rect 6163 28318 6178 28364
rect 6224 28318 6239 28364
rect 6163 28261 6239 28318
rect 6163 28215 6178 28261
rect 6224 28215 6239 28261
rect 6163 28158 6239 28215
rect 6163 28112 6178 28158
rect 6224 28112 6239 28158
rect 6163 28055 6239 28112
rect 6163 28009 6178 28055
rect 6224 28009 6239 28055
rect 6163 27952 6239 28009
rect 6163 27906 6178 27952
rect 6224 27906 6239 27952
rect 6163 27848 6239 27906
rect 6163 27802 6178 27848
rect 6224 27802 6239 27848
rect 6163 27729 6239 27802
rect 6407 28776 6483 29003
rect 6407 28730 6422 28776
rect 6468 28730 6483 28776
rect 6407 28673 6483 28730
rect 6407 28627 6422 28673
rect 6468 28627 6483 28673
rect 6407 28570 6483 28627
rect 6407 28524 6422 28570
rect 6468 28524 6483 28570
rect 6407 28467 6483 28524
rect 6407 28421 6422 28467
rect 6468 28421 6483 28467
rect 6407 28364 6483 28421
rect 6407 28318 6422 28364
rect 6468 28318 6483 28364
rect 6407 28261 6483 28318
rect 6407 28215 6422 28261
rect 6468 28215 6483 28261
rect 6407 28158 6483 28215
rect 6407 28112 6422 28158
rect 6468 28112 6483 28158
rect 6407 28055 6483 28112
rect 6407 28009 6422 28055
rect 6468 28009 6483 28055
rect 6407 27952 6483 28009
rect 6407 27906 6422 27952
rect 6468 27906 6483 27952
rect 6407 27848 6483 27906
rect 6407 27802 6422 27848
rect 6468 27802 6483 27848
rect 6407 27789 6483 27802
rect 6651 28776 6727 28789
rect 6651 28730 6666 28776
rect 6712 28730 6727 28776
rect 6651 28673 6727 28730
rect 6651 28627 6666 28673
rect 6712 28627 6727 28673
rect 6651 28570 6727 28627
rect 6651 28524 6666 28570
rect 6712 28524 6727 28570
rect 6651 28467 6727 28524
rect 6651 28421 6666 28467
rect 6712 28421 6727 28467
rect 6651 28364 6727 28421
rect 6651 28318 6666 28364
rect 6712 28318 6727 28364
rect 6651 28261 6727 28318
rect 6651 28215 6666 28261
rect 6712 28215 6727 28261
rect 6651 28158 6727 28215
rect 6651 28112 6666 28158
rect 6712 28112 6727 28158
rect 6651 28055 6727 28112
rect 6651 28009 6666 28055
rect 6712 28009 6727 28055
rect 6651 27952 6727 28009
rect 6651 27906 6666 27952
rect 6712 27906 6727 27952
rect 6651 27848 6727 27906
rect 6651 27802 6666 27848
rect 6712 27802 6727 27848
rect 6651 27729 6727 27802
rect 6895 28776 6971 29003
rect 6895 28730 6910 28776
rect 6956 28730 6971 28776
rect 6895 28673 6971 28730
rect 6895 28627 6910 28673
rect 6956 28627 6971 28673
rect 6895 28570 6971 28627
rect 6895 28524 6910 28570
rect 6956 28524 6971 28570
rect 6895 28467 6971 28524
rect 6895 28421 6910 28467
rect 6956 28421 6971 28467
rect 6895 28364 6971 28421
rect 6895 28318 6910 28364
rect 6956 28318 6971 28364
rect 6895 28261 6971 28318
rect 6895 28215 6910 28261
rect 6956 28215 6971 28261
rect 6895 28158 6971 28215
rect 6895 28112 6910 28158
rect 6956 28112 6971 28158
rect 6895 28055 6971 28112
rect 6895 28009 6910 28055
rect 6956 28009 6971 28055
rect 6895 27952 6971 28009
rect 6895 27906 6910 27952
rect 6956 27906 6971 27952
rect 6895 27848 6971 27906
rect 6895 27802 6910 27848
rect 6956 27802 6971 27848
rect 6895 27789 6971 27802
rect 7139 28776 7215 28789
rect 7139 28730 7154 28776
rect 7200 28730 7215 28776
rect 7139 28673 7215 28730
rect 7139 28627 7154 28673
rect 7200 28627 7215 28673
rect 7139 28570 7215 28627
rect 7139 28524 7154 28570
rect 7200 28524 7215 28570
rect 7139 28467 7215 28524
rect 7139 28421 7154 28467
rect 7200 28421 7215 28467
rect 7139 28364 7215 28421
rect 7139 28318 7154 28364
rect 7200 28318 7215 28364
rect 7139 28261 7215 28318
rect 7139 28215 7154 28261
rect 7200 28215 7215 28261
rect 7139 28158 7215 28215
rect 7139 28112 7154 28158
rect 7200 28112 7215 28158
rect 7139 28055 7215 28112
rect 7139 28009 7154 28055
rect 7200 28009 7215 28055
rect 7139 27952 7215 28009
rect 7139 27906 7154 27952
rect 7200 27906 7215 27952
rect 7139 27848 7215 27906
rect 7139 27802 7154 27848
rect 7200 27802 7215 27848
rect 7139 27729 7215 27802
rect 7383 28776 7459 29003
rect 7383 28730 7398 28776
rect 7444 28730 7459 28776
rect 7383 28673 7459 28730
rect 7383 28627 7398 28673
rect 7444 28627 7459 28673
rect 7383 28570 7459 28627
rect 7383 28524 7398 28570
rect 7444 28524 7459 28570
rect 7383 28467 7459 28524
rect 7383 28421 7398 28467
rect 7444 28421 7459 28467
rect 7383 28364 7459 28421
rect 7383 28318 7398 28364
rect 7444 28318 7459 28364
rect 7383 28261 7459 28318
rect 7383 28215 7398 28261
rect 7444 28215 7459 28261
rect 7383 28158 7459 28215
rect 7383 28112 7398 28158
rect 7444 28112 7459 28158
rect 7383 28055 7459 28112
rect 7383 28009 7398 28055
rect 7444 28009 7459 28055
rect 7383 27952 7459 28009
rect 7383 27906 7398 27952
rect 7444 27906 7459 27952
rect 7383 27848 7459 27906
rect 7383 27802 7398 27848
rect 7444 27802 7459 27848
rect 7383 27789 7459 27802
rect 7627 28776 7703 28789
rect 7627 28730 7642 28776
rect 7688 28730 7703 28776
rect 7627 28673 7703 28730
rect 7627 28627 7642 28673
rect 7688 28627 7703 28673
rect 7627 28570 7703 28627
rect 7627 28524 7642 28570
rect 7688 28524 7703 28570
rect 7627 28467 7703 28524
rect 7627 28421 7642 28467
rect 7688 28421 7703 28467
rect 7627 28364 7703 28421
rect 7627 28318 7642 28364
rect 7688 28318 7703 28364
rect 7627 28261 7703 28318
rect 7627 28215 7642 28261
rect 7688 28215 7703 28261
rect 7627 28158 7703 28215
rect 7627 28112 7642 28158
rect 7688 28112 7703 28158
rect 7627 28055 7703 28112
rect 7627 28009 7642 28055
rect 7688 28009 7703 28055
rect 7627 27952 7703 28009
rect 7627 27906 7642 27952
rect 7688 27906 7703 27952
rect 7627 27848 7703 27906
rect 7627 27802 7642 27848
rect 7688 27802 7703 27848
rect 7627 27729 7703 27802
rect 7871 28776 7947 29003
rect 7871 28730 7886 28776
rect 7932 28730 7947 28776
rect 7871 28673 7947 28730
rect 7871 28627 7886 28673
rect 7932 28627 7947 28673
rect 7871 28570 7947 28627
rect 7871 28524 7886 28570
rect 7932 28524 7947 28570
rect 7871 28467 7947 28524
rect 7871 28421 7886 28467
rect 7932 28421 7947 28467
rect 7871 28364 7947 28421
rect 7871 28318 7886 28364
rect 7932 28318 7947 28364
rect 7871 28261 7947 28318
rect 7871 28215 7886 28261
rect 7932 28215 7947 28261
rect 7871 28158 7947 28215
rect 7871 28112 7886 28158
rect 7932 28112 7947 28158
rect 7871 28055 7947 28112
rect 7871 28009 7886 28055
rect 7932 28009 7947 28055
rect 7871 27952 7947 28009
rect 7871 27906 7886 27952
rect 7932 27906 7947 27952
rect 7871 27848 7947 27906
rect 7871 27802 7886 27848
rect 7932 27802 7947 27848
rect 7871 27789 7947 27802
rect 8115 28776 8191 28789
rect 8115 28730 8130 28776
rect 8176 28730 8191 28776
rect 8115 28673 8191 28730
rect 8115 28627 8130 28673
rect 8176 28627 8191 28673
rect 8115 28570 8191 28627
rect 8115 28524 8130 28570
rect 8176 28524 8191 28570
rect 8115 28467 8191 28524
rect 8115 28421 8130 28467
rect 8176 28421 8191 28467
rect 8115 28364 8191 28421
rect 8115 28318 8130 28364
rect 8176 28318 8191 28364
rect 8115 28261 8191 28318
rect 8115 28215 8130 28261
rect 8176 28215 8191 28261
rect 8115 28158 8191 28215
rect 8115 28112 8130 28158
rect 8176 28112 8191 28158
rect 8115 28055 8191 28112
rect 8115 28009 8130 28055
rect 8176 28009 8191 28055
rect 8115 27952 8191 28009
rect 8115 27906 8130 27952
rect 8176 27906 8191 27952
rect 8115 27848 8191 27906
rect 8115 27802 8130 27848
rect 8176 27802 8191 27848
rect 8115 27729 8191 27802
rect 8359 28776 8435 29003
rect 8359 28730 8374 28776
rect 8420 28730 8435 28776
rect 8359 28673 8435 28730
rect 8359 28627 8374 28673
rect 8420 28627 8435 28673
rect 8359 28570 8435 28627
rect 8359 28524 8374 28570
rect 8420 28524 8435 28570
rect 8359 28467 8435 28524
rect 8359 28421 8374 28467
rect 8420 28421 8435 28467
rect 8359 28364 8435 28421
rect 8359 28318 8374 28364
rect 8420 28318 8435 28364
rect 8359 28261 8435 28318
rect 8359 28215 8374 28261
rect 8420 28215 8435 28261
rect 8359 28158 8435 28215
rect 8359 28112 8374 28158
rect 8420 28112 8435 28158
rect 8359 28055 8435 28112
rect 8359 28009 8374 28055
rect 8420 28009 8435 28055
rect 8359 27952 8435 28009
rect 8359 27906 8374 27952
rect 8420 27906 8435 27952
rect 8359 27848 8435 27906
rect 8359 27802 8374 27848
rect 8420 27802 8435 27848
rect 8359 27789 8435 27802
rect 8603 28776 8679 28789
rect 8603 28730 8618 28776
rect 8664 28730 8679 28776
rect 8603 28673 8679 28730
rect 8603 28627 8618 28673
rect 8664 28627 8679 28673
rect 8603 28570 8679 28627
rect 8603 28524 8618 28570
rect 8664 28524 8679 28570
rect 8603 28467 8679 28524
rect 8603 28421 8618 28467
rect 8664 28421 8679 28467
rect 8603 28364 8679 28421
rect 8603 28318 8618 28364
rect 8664 28318 8679 28364
rect 8603 28261 8679 28318
rect 8603 28215 8618 28261
rect 8664 28215 8679 28261
rect 8603 28158 8679 28215
rect 8603 28112 8618 28158
rect 8664 28112 8679 28158
rect 8603 28055 8679 28112
rect 8603 28009 8618 28055
rect 8664 28009 8679 28055
rect 8603 27952 8679 28009
rect 8603 27906 8618 27952
rect 8664 27906 8679 27952
rect 8603 27848 8679 27906
rect 8603 27802 8618 27848
rect 8664 27802 8679 27848
rect 8603 27729 8679 27802
rect 8847 28776 8923 29003
rect 8847 28730 8862 28776
rect 8908 28730 8923 28776
rect 8847 28673 8923 28730
rect 8847 28627 8862 28673
rect 8908 28627 8923 28673
rect 8847 28570 8923 28627
rect 8847 28524 8862 28570
rect 8908 28524 8923 28570
rect 8847 28467 8923 28524
rect 8847 28421 8862 28467
rect 8908 28421 8923 28467
rect 8847 28364 8923 28421
rect 8847 28318 8862 28364
rect 8908 28318 8923 28364
rect 8847 28261 8923 28318
rect 8847 28215 8862 28261
rect 8908 28215 8923 28261
rect 8847 28158 8923 28215
rect 8847 28112 8862 28158
rect 8908 28112 8923 28158
rect 8847 28055 8923 28112
rect 8847 28009 8862 28055
rect 8908 28009 8923 28055
rect 8847 27952 8923 28009
rect 8847 27906 8862 27952
rect 8908 27906 8923 27952
rect 8847 27848 8923 27906
rect 8847 27802 8862 27848
rect 8908 27802 8923 27848
rect 8847 27789 8923 27802
rect 9091 28776 9167 28789
rect 9091 28730 9106 28776
rect 9152 28730 9167 28776
rect 9091 28673 9167 28730
rect 9091 28627 9106 28673
rect 9152 28627 9167 28673
rect 9091 28570 9167 28627
rect 9091 28524 9106 28570
rect 9152 28524 9167 28570
rect 9091 28467 9167 28524
rect 9091 28421 9106 28467
rect 9152 28421 9167 28467
rect 9091 28364 9167 28421
rect 9091 28318 9106 28364
rect 9152 28318 9167 28364
rect 9091 28261 9167 28318
rect 9091 28215 9106 28261
rect 9152 28215 9167 28261
rect 9091 28158 9167 28215
rect 9091 28112 9106 28158
rect 9152 28112 9167 28158
rect 9091 28055 9167 28112
rect 9091 28009 9106 28055
rect 9152 28009 9167 28055
rect 9091 27952 9167 28009
rect 9091 27906 9106 27952
rect 9152 27906 9167 27952
rect 9091 27848 9167 27906
rect 9091 27802 9106 27848
rect 9152 27802 9167 27848
rect 9091 27729 9167 27802
rect 9335 28776 9411 29003
rect 9335 28730 9350 28776
rect 9396 28730 9411 28776
rect 9335 28673 9411 28730
rect 9335 28627 9350 28673
rect 9396 28627 9411 28673
rect 9335 28570 9411 28627
rect 9335 28524 9350 28570
rect 9396 28524 9411 28570
rect 9335 28467 9411 28524
rect 9335 28421 9350 28467
rect 9396 28421 9411 28467
rect 9335 28364 9411 28421
rect 9335 28318 9350 28364
rect 9396 28318 9411 28364
rect 9335 28261 9411 28318
rect 9335 28215 9350 28261
rect 9396 28215 9411 28261
rect 9335 28158 9411 28215
rect 9335 28112 9350 28158
rect 9396 28112 9411 28158
rect 9335 28055 9411 28112
rect 9335 28009 9350 28055
rect 9396 28009 9411 28055
rect 9335 27952 9411 28009
rect 9335 27906 9350 27952
rect 9396 27906 9411 27952
rect 9335 27848 9411 27906
rect 9335 27802 9350 27848
rect 9396 27802 9411 27848
rect 9335 27789 9411 27802
rect 9579 28776 9655 28789
rect 9579 28730 9594 28776
rect 9640 28730 9655 28776
rect 9579 28673 9655 28730
rect 9579 28627 9594 28673
rect 9640 28627 9655 28673
rect 9579 28570 9655 28627
rect 9579 28524 9594 28570
rect 9640 28524 9655 28570
rect 9579 28467 9655 28524
rect 9579 28421 9594 28467
rect 9640 28421 9655 28467
rect 9579 28364 9655 28421
rect 9579 28318 9594 28364
rect 9640 28318 9655 28364
rect 9579 28261 9655 28318
rect 9579 28215 9594 28261
rect 9640 28215 9655 28261
rect 9579 28158 9655 28215
rect 9579 28112 9594 28158
rect 9640 28112 9655 28158
rect 9579 28055 9655 28112
rect 9579 28009 9594 28055
rect 9640 28009 9655 28055
rect 9579 27952 9655 28009
rect 9579 27906 9594 27952
rect 9640 27906 9655 27952
rect 9579 27848 9655 27906
rect 9579 27802 9594 27848
rect 9640 27802 9655 27848
rect 9579 27729 9655 27802
rect 9823 28776 9899 29003
rect 9823 28730 9838 28776
rect 9884 28730 9899 28776
rect 9823 28673 9899 28730
rect 9823 28627 9838 28673
rect 9884 28627 9899 28673
rect 9823 28570 9899 28627
rect 9823 28524 9838 28570
rect 9884 28524 9899 28570
rect 9823 28467 9899 28524
rect 9823 28421 9838 28467
rect 9884 28421 9899 28467
rect 9823 28364 9899 28421
rect 9823 28318 9838 28364
rect 9884 28318 9899 28364
rect 9823 28261 9899 28318
rect 9823 28215 9838 28261
rect 9884 28215 9899 28261
rect 9823 28158 9899 28215
rect 9823 28112 9838 28158
rect 9884 28112 9899 28158
rect 9823 28055 9899 28112
rect 9823 28009 9838 28055
rect 9884 28009 9899 28055
rect 9823 27952 9899 28009
rect 9823 27906 9838 27952
rect 9884 27906 9899 27952
rect 9823 27848 9899 27906
rect 9823 27802 9838 27848
rect 9884 27802 9899 27848
rect 9823 27789 9899 27802
rect 10067 28776 10143 28789
rect 10067 28730 10082 28776
rect 10128 28730 10143 28776
rect 10067 28673 10143 28730
rect 10067 28627 10082 28673
rect 10128 28627 10143 28673
rect 10067 28570 10143 28627
rect 10067 28524 10082 28570
rect 10128 28524 10143 28570
rect 10067 28467 10143 28524
rect 10067 28421 10082 28467
rect 10128 28421 10143 28467
rect 10067 28364 10143 28421
rect 10067 28318 10082 28364
rect 10128 28318 10143 28364
rect 10067 28261 10143 28318
rect 10067 28215 10082 28261
rect 10128 28215 10143 28261
rect 10067 28158 10143 28215
rect 10067 28112 10082 28158
rect 10128 28112 10143 28158
rect 10067 28055 10143 28112
rect 10067 28009 10082 28055
rect 10128 28009 10143 28055
rect 10067 27952 10143 28009
rect 10067 27906 10082 27952
rect 10128 27906 10143 27952
rect 10067 27848 10143 27906
rect 10067 27802 10082 27848
rect 10128 27802 10143 27848
rect 10067 27729 10143 27802
rect 10311 28776 10387 29003
rect 10311 28730 10326 28776
rect 10372 28730 10387 28776
rect 10311 28673 10387 28730
rect 10311 28627 10326 28673
rect 10372 28627 10387 28673
rect 10311 28570 10387 28627
rect 10311 28524 10326 28570
rect 10372 28524 10387 28570
rect 10311 28467 10387 28524
rect 10311 28421 10326 28467
rect 10372 28421 10387 28467
rect 10311 28364 10387 28421
rect 10311 28318 10326 28364
rect 10372 28318 10387 28364
rect 10311 28261 10387 28318
rect 10311 28215 10326 28261
rect 10372 28215 10387 28261
rect 10311 28158 10387 28215
rect 10311 28112 10326 28158
rect 10372 28112 10387 28158
rect 10311 28055 10387 28112
rect 10311 28009 10326 28055
rect 10372 28009 10387 28055
rect 10311 27952 10387 28009
rect 10311 27906 10326 27952
rect 10372 27906 10387 27952
rect 10311 27848 10387 27906
rect 10311 27802 10326 27848
rect 10372 27802 10387 27848
rect 10311 27789 10387 27802
rect 10630 28906 10698 29003
rect 10630 27732 10641 28906
rect 10687 27732 10698 28906
rect 4699 27653 10433 27729
rect 10630 27721 10698 27732
rect 3551 27597 3627 27653
rect -1 27582 3464 27593
rect -1 27536 2749 27582
rect 3453 27536 3464 27582
rect -1 27393 3464 27536
rect 2264 27156 2332 27167
rect 2264 25888 2275 27156
rect 2321 25888 2332 27156
rect 3388 27146 3464 27393
rect 3551 27582 4224 27597
rect 3551 27536 3697 27582
rect 4213 27536 4224 27582
rect 3551 27521 4224 27536
rect 4283 27593 4359 27653
rect 4283 27582 10275 27593
rect 4283 27536 4578 27582
rect 10264 27536 10275 27582
rect 3551 27274 3627 27521
rect 4283 27517 10275 27536
rect 3551 27259 6516 27274
rect 3551 27213 5237 27259
rect 6505 27213 6516 27259
rect 3551 27198 6516 27213
rect 6652 27270 6728 27517
rect 6652 27259 7980 27270
rect 6652 27213 6701 27259
rect 7969 27213 7980 27259
rect 6652 27202 7980 27213
rect 3388 27131 4223 27146
rect 3388 27085 4072 27131
rect 4212 27085 4223 27131
rect 3388 27070 4223 27085
rect 2264 25791 2332 25888
rect 4039 26993 4115 27006
rect 4039 26947 4054 26993
rect 4100 26947 4115 26993
rect 4039 26890 4115 26947
rect 4039 26844 4054 26890
rect 4100 26844 4115 26890
rect 4039 26787 4115 26844
rect 4039 26741 4054 26787
rect 4100 26741 4115 26787
rect 4039 26684 4115 26741
rect 4039 26638 4054 26684
rect 4100 26638 4115 26684
rect 4039 26581 4115 26638
rect 4039 26535 4054 26581
rect 4100 26535 4115 26581
rect 4039 26478 4115 26535
rect 4039 26432 4054 26478
rect 4100 26432 4115 26478
rect 4039 26375 4115 26432
rect 4039 26329 4054 26375
rect 4100 26329 4115 26375
rect 4039 26272 4115 26329
rect 4039 26226 4054 26272
rect 4100 26226 4115 26272
rect 4039 26169 4115 26226
rect 4039 26123 4054 26169
rect 4100 26123 4115 26169
rect 4039 26065 4115 26123
rect 4039 26019 4054 26065
rect 4100 26019 4115 26065
rect 4039 25791 4115 26019
rect 4283 26993 4359 27198
rect 6652 27142 6728 27202
rect 10357 27142 10433 27653
rect 5345 27066 6728 27142
rect 6809 27066 10433 27142
rect 10630 27156 10698 27167
rect 4283 26947 4298 26993
rect 4344 26947 4359 26993
rect 4283 26890 4359 26947
rect 4283 26844 4298 26890
rect 4344 26844 4359 26890
rect 4283 26787 4359 26844
rect 4283 26741 4298 26787
rect 4344 26741 4359 26787
rect 4283 26684 4359 26741
rect 4283 26638 4298 26684
rect 4344 26638 4359 26684
rect 4283 26581 4359 26638
rect 4283 26535 4298 26581
rect 4344 26535 4359 26581
rect 4283 26478 4359 26535
rect 4283 26432 4298 26478
rect 4344 26432 4359 26478
rect 4283 26375 4359 26432
rect 4283 26329 4298 26375
rect 4344 26329 4359 26375
rect 4283 26272 4359 26329
rect 4283 26226 4298 26272
rect 4344 26226 4359 26272
rect 4283 26169 4359 26226
rect 4283 26123 4298 26169
rect 4344 26123 4359 26169
rect 4283 26065 4359 26123
rect 4283 26019 4298 26065
rect 4344 26019 4359 26065
rect 4283 26006 4359 26019
rect 5101 26993 5177 27006
rect 5101 26947 5116 26993
rect 5162 26947 5177 26993
rect 5101 26890 5177 26947
rect 5101 26844 5116 26890
rect 5162 26844 5177 26890
rect 5101 26787 5177 26844
rect 5101 26741 5116 26787
rect 5162 26741 5177 26787
rect 5101 26684 5177 26741
rect 5101 26638 5116 26684
rect 5162 26638 5177 26684
rect 5101 26581 5177 26638
rect 5101 26535 5116 26581
rect 5162 26535 5177 26581
rect 5101 26478 5177 26535
rect 5101 26432 5116 26478
rect 5162 26432 5177 26478
rect 5101 26375 5177 26432
rect 5101 26329 5116 26375
rect 5162 26329 5177 26375
rect 5101 26272 5177 26329
rect 5101 26226 5116 26272
rect 5162 26226 5177 26272
rect 5101 26169 5177 26226
rect 5101 26123 5116 26169
rect 5162 26123 5177 26169
rect 5101 26065 5177 26123
rect 5101 26019 5116 26065
rect 5162 26019 5177 26065
rect 5101 25791 5177 26019
rect 5345 26993 5421 27066
rect 5345 26947 5360 26993
rect 5406 26947 5421 26993
rect 5345 26890 5421 26947
rect 5345 26844 5360 26890
rect 5406 26844 5421 26890
rect 5345 26787 5421 26844
rect 5345 26741 5360 26787
rect 5406 26741 5421 26787
rect 5345 26684 5421 26741
rect 5345 26638 5360 26684
rect 5406 26638 5421 26684
rect 5345 26581 5421 26638
rect 5345 26535 5360 26581
rect 5406 26535 5421 26581
rect 5345 26478 5421 26535
rect 5345 26432 5360 26478
rect 5406 26432 5421 26478
rect 5345 26375 5421 26432
rect 5345 26329 5360 26375
rect 5406 26329 5421 26375
rect 5345 26272 5421 26329
rect 5345 26226 5360 26272
rect 5406 26226 5421 26272
rect 5345 26169 5421 26226
rect 5345 26123 5360 26169
rect 5406 26123 5421 26169
rect 5345 26065 5421 26123
rect 5345 26019 5360 26065
rect 5406 26019 5421 26065
rect 5345 26006 5421 26019
rect 5589 26993 5665 27006
rect 5589 26947 5604 26993
rect 5650 26947 5665 26993
rect 5589 26890 5665 26947
rect 5589 26844 5604 26890
rect 5650 26844 5665 26890
rect 5589 26787 5665 26844
rect 5589 26741 5604 26787
rect 5650 26741 5665 26787
rect 5589 26684 5665 26741
rect 5589 26638 5604 26684
rect 5650 26638 5665 26684
rect 5589 26581 5665 26638
rect 5589 26535 5604 26581
rect 5650 26535 5665 26581
rect 5589 26478 5665 26535
rect 5589 26432 5604 26478
rect 5650 26432 5665 26478
rect 5589 26375 5665 26432
rect 5589 26329 5604 26375
rect 5650 26329 5665 26375
rect 5589 26272 5665 26329
rect 5589 26226 5604 26272
rect 5650 26226 5665 26272
rect 5589 26169 5665 26226
rect 5589 26123 5604 26169
rect 5650 26123 5665 26169
rect 5589 26065 5665 26123
rect 5589 26019 5604 26065
rect 5650 26019 5665 26065
rect 5589 25791 5665 26019
rect 5833 26993 5909 27066
rect 5833 26947 5848 26993
rect 5894 26947 5909 26993
rect 5833 26890 5909 26947
rect 5833 26844 5848 26890
rect 5894 26844 5909 26890
rect 5833 26787 5909 26844
rect 5833 26741 5848 26787
rect 5894 26741 5909 26787
rect 5833 26684 5909 26741
rect 5833 26638 5848 26684
rect 5894 26638 5909 26684
rect 5833 26581 5909 26638
rect 5833 26535 5848 26581
rect 5894 26535 5909 26581
rect 5833 26478 5909 26535
rect 5833 26432 5848 26478
rect 5894 26432 5909 26478
rect 5833 26375 5909 26432
rect 5833 26329 5848 26375
rect 5894 26329 5909 26375
rect 5833 26272 5909 26329
rect 5833 26226 5848 26272
rect 5894 26226 5909 26272
rect 5833 26169 5909 26226
rect 5833 26123 5848 26169
rect 5894 26123 5909 26169
rect 5833 26065 5909 26123
rect 5833 26019 5848 26065
rect 5894 26019 5909 26065
rect 5833 26006 5909 26019
rect 6077 26993 6153 27006
rect 6077 26947 6092 26993
rect 6138 26947 6153 26993
rect 6077 26890 6153 26947
rect 6077 26844 6092 26890
rect 6138 26844 6153 26890
rect 6077 26787 6153 26844
rect 6077 26741 6092 26787
rect 6138 26741 6153 26787
rect 6077 26684 6153 26741
rect 6077 26638 6092 26684
rect 6138 26638 6153 26684
rect 6077 26581 6153 26638
rect 6077 26535 6092 26581
rect 6138 26535 6153 26581
rect 6077 26478 6153 26535
rect 6077 26432 6092 26478
rect 6138 26432 6153 26478
rect 6077 26375 6153 26432
rect 6077 26329 6092 26375
rect 6138 26329 6153 26375
rect 6077 26272 6153 26329
rect 6077 26226 6092 26272
rect 6138 26226 6153 26272
rect 6077 26169 6153 26226
rect 6077 26123 6092 26169
rect 6138 26123 6153 26169
rect 6077 26065 6153 26123
rect 6077 26019 6092 26065
rect 6138 26019 6153 26065
rect 6077 25791 6153 26019
rect 6321 26993 6397 27066
rect 6321 26947 6336 26993
rect 6382 26947 6397 26993
rect 6321 26890 6397 26947
rect 6321 26844 6336 26890
rect 6382 26844 6397 26890
rect 6321 26787 6397 26844
rect 6321 26741 6336 26787
rect 6382 26741 6397 26787
rect 6321 26684 6397 26741
rect 6321 26638 6336 26684
rect 6382 26638 6397 26684
rect 6321 26581 6397 26638
rect 6321 26535 6336 26581
rect 6382 26535 6397 26581
rect 6321 26478 6397 26535
rect 6321 26432 6336 26478
rect 6382 26432 6397 26478
rect 6321 26375 6397 26432
rect 6321 26329 6336 26375
rect 6382 26329 6397 26375
rect 6321 26272 6397 26329
rect 6321 26226 6336 26272
rect 6382 26226 6397 26272
rect 6321 26169 6397 26226
rect 6321 26123 6336 26169
rect 6382 26123 6397 26169
rect 6321 26065 6397 26123
rect 6321 26019 6336 26065
rect 6382 26019 6397 26065
rect 6321 26006 6397 26019
rect 6565 26993 6641 27006
rect 6565 26947 6580 26993
rect 6626 26947 6641 26993
rect 6565 26890 6641 26947
rect 6565 26844 6580 26890
rect 6626 26844 6641 26890
rect 6565 26787 6641 26844
rect 6565 26741 6580 26787
rect 6626 26741 6641 26787
rect 6565 26684 6641 26741
rect 6565 26638 6580 26684
rect 6626 26638 6641 26684
rect 6565 26581 6641 26638
rect 6565 26535 6580 26581
rect 6626 26535 6641 26581
rect 6565 26478 6641 26535
rect 6565 26432 6580 26478
rect 6626 26432 6641 26478
rect 6565 26375 6641 26432
rect 6565 26329 6580 26375
rect 6626 26329 6641 26375
rect 6565 26272 6641 26329
rect 6565 26226 6580 26272
rect 6626 26226 6641 26272
rect 6565 26169 6641 26226
rect 6565 26123 6580 26169
rect 6626 26123 6641 26169
rect 6565 26065 6641 26123
rect 6565 26019 6580 26065
rect 6626 26019 6641 26065
rect 6565 25791 6641 26019
rect 6809 26993 6885 27066
rect 6809 26947 6824 26993
rect 6870 26947 6885 26993
rect 6809 26890 6885 26947
rect 6809 26844 6824 26890
rect 6870 26844 6885 26890
rect 6809 26787 6885 26844
rect 6809 26741 6824 26787
rect 6870 26741 6885 26787
rect 6809 26684 6885 26741
rect 6809 26638 6824 26684
rect 6870 26638 6885 26684
rect 6809 26581 6885 26638
rect 6809 26535 6824 26581
rect 6870 26535 6885 26581
rect 6809 26478 6885 26535
rect 6809 26432 6824 26478
rect 6870 26432 6885 26478
rect 6809 26375 6885 26432
rect 6809 26329 6824 26375
rect 6870 26329 6885 26375
rect 6809 26272 6885 26329
rect 6809 26226 6824 26272
rect 6870 26226 6885 26272
rect 6809 26169 6885 26226
rect 6809 26123 6824 26169
rect 6870 26123 6885 26169
rect 6809 26065 6885 26123
rect 6809 26019 6824 26065
rect 6870 26019 6885 26065
rect 2264 25780 6759 25791
rect 2264 25734 2275 25780
rect 6739 25734 6759 25780
rect 2264 25723 6759 25734
rect 6809 25617 6885 26019
rect 7053 26993 7129 27006
rect 7053 26947 7068 26993
rect 7114 26947 7129 26993
rect 7053 26890 7129 26947
rect 7053 26844 7068 26890
rect 7114 26844 7129 26890
rect 7053 26787 7129 26844
rect 7053 26741 7068 26787
rect 7114 26741 7129 26787
rect 7053 26684 7129 26741
rect 7053 26638 7068 26684
rect 7114 26638 7129 26684
rect 7053 26581 7129 26638
rect 7053 26535 7068 26581
rect 7114 26535 7129 26581
rect 7053 26478 7129 26535
rect 7053 26432 7068 26478
rect 7114 26432 7129 26478
rect 7053 26375 7129 26432
rect 7053 26329 7068 26375
rect 7114 26329 7129 26375
rect 7053 26272 7129 26329
rect 7053 26226 7068 26272
rect 7114 26226 7129 26272
rect 7053 26169 7129 26226
rect 7053 26123 7068 26169
rect 7114 26123 7129 26169
rect 7053 26065 7129 26123
rect 7053 26019 7068 26065
rect 7114 26019 7129 26065
rect 7053 25791 7129 26019
rect 7297 26993 7373 27066
rect 7297 26947 7312 26993
rect 7358 26947 7373 26993
rect 7297 26890 7373 26947
rect 7297 26844 7312 26890
rect 7358 26844 7373 26890
rect 7297 26787 7373 26844
rect 7297 26741 7312 26787
rect 7358 26741 7373 26787
rect 7297 26684 7373 26741
rect 7297 26638 7312 26684
rect 7358 26638 7373 26684
rect 7297 26581 7373 26638
rect 7297 26535 7312 26581
rect 7358 26535 7373 26581
rect 7297 26478 7373 26535
rect 7297 26432 7312 26478
rect 7358 26432 7373 26478
rect 7297 26375 7373 26432
rect 7297 26329 7312 26375
rect 7358 26329 7373 26375
rect 7297 26272 7373 26329
rect 7297 26226 7312 26272
rect 7358 26226 7373 26272
rect 7297 26169 7373 26226
rect 7297 26123 7312 26169
rect 7358 26123 7373 26169
rect 7297 26065 7373 26123
rect 7297 26019 7312 26065
rect 7358 26019 7373 26065
rect 7297 25979 7373 26019
rect 7541 26993 7617 27006
rect 7541 26947 7556 26993
rect 7602 26947 7617 26993
rect 7541 26890 7617 26947
rect 7541 26844 7556 26890
rect 7602 26844 7617 26890
rect 7541 26787 7617 26844
rect 7541 26741 7556 26787
rect 7602 26741 7617 26787
rect 7541 26684 7617 26741
rect 7541 26638 7556 26684
rect 7602 26638 7617 26684
rect 7541 26581 7617 26638
rect 7541 26535 7556 26581
rect 7602 26535 7617 26581
rect 7541 26478 7617 26535
rect 7541 26432 7556 26478
rect 7602 26432 7617 26478
rect 7541 26375 7617 26432
rect 7541 26329 7556 26375
rect 7602 26329 7617 26375
rect 7541 26272 7617 26329
rect 7541 26226 7556 26272
rect 7602 26226 7617 26272
rect 7541 26169 7617 26226
rect 7541 26123 7556 26169
rect 7602 26123 7617 26169
rect 7541 26065 7617 26123
rect 7541 26019 7556 26065
rect 7602 26019 7617 26065
rect 7541 25791 7617 26019
rect 7785 26993 7861 27066
rect 7785 26947 7800 26993
rect 7846 26947 7861 26993
rect 7785 26890 7861 26947
rect 7785 26844 7800 26890
rect 7846 26844 7861 26890
rect 7785 26787 7861 26844
rect 7785 26741 7800 26787
rect 7846 26741 7861 26787
rect 7785 26684 7861 26741
rect 7785 26638 7800 26684
rect 7846 26638 7861 26684
rect 7785 26581 7861 26638
rect 7785 26535 7800 26581
rect 7846 26535 7861 26581
rect 7785 26478 7861 26535
rect 7785 26432 7800 26478
rect 7846 26432 7861 26478
rect 7785 26375 7861 26432
rect 7785 26329 7800 26375
rect 7846 26329 7861 26375
rect 7785 26272 7861 26329
rect 7785 26226 7800 26272
rect 7846 26226 7861 26272
rect 7785 26169 7861 26226
rect 7785 26123 7800 26169
rect 7846 26123 7861 26169
rect 7785 26065 7861 26123
rect 7785 26019 7800 26065
rect 7846 26019 7861 26065
rect 7785 25979 7861 26019
rect 8029 26993 8105 27006
rect 8029 26947 8044 26993
rect 8090 26947 8105 26993
rect 8029 26890 8105 26947
rect 8029 26844 8044 26890
rect 8090 26844 8105 26890
rect 8029 26787 8105 26844
rect 8029 26741 8044 26787
rect 8090 26741 8105 26787
rect 8029 26684 8105 26741
rect 8029 26638 8044 26684
rect 8090 26638 8105 26684
rect 8029 26581 8105 26638
rect 8029 26535 8044 26581
rect 8090 26535 8105 26581
rect 8029 26478 8105 26535
rect 8029 26432 8044 26478
rect 8090 26432 8105 26478
rect 8029 26375 8105 26432
rect 8029 26329 8044 26375
rect 8090 26329 8105 26375
rect 8029 26272 8105 26329
rect 8029 26226 8044 26272
rect 8090 26226 8105 26272
rect 8029 26169 8105 26226
rect 8029 26123 8044 26169
rect 8090 26123 8105 26169
rect 8029 26065 8105 26123
rect 8029 26019 8044 26065
rect 8090 26019 8105 26065
rect 8029 25791 8105 26019
rect 10630 25888 10641 27156
rect 10687 25888 10698 27156
rect 10630 25791 10698 25888
rect 6935 25780 7247 25791
rect 6935 25734 6975 25780
rect 7209 25734 7247 25780
rect 6935 25723 7247 25734
rect 7423 25780 7735 25791
rect 7423 25734 7445 25780
rect 7679 25734 7735 25780
rect 7423 25723 7735 25734
rect 7911 25780 10698 25791
rect 7911 25734 8009 25780
rect 10687 25734 10698 25780
rect 7911 25723 10698 25734
rect 1213 25597 11749 25617
rect 1213 25545 1233 25597
rect 1285 25545 1341 25597
rect 1393 25545 11569 25597
rect 11621 25545 11677 25597
rect 11729 25545 11749 25597
rect 1213 25489 11749 25545
rect 1213 25437 1233 25489
rect 1285 25437 1341 25489
rect 1393 25437 11569 25489
rect 11621 25437 11677 25489
rect 11729 25437 11749 25489
rect 1213 25417 11749 25437
<< via1 >>
rect 1233 25545 1285 25597
rect 1341 25545 1393 25597
rect 11569 25545 11621 25597
rect 11677 25545 11729 25597
rect 1233 25437 1285 25489
rect 1341 25437 1393 25489
rect 11569 25437 11621 25489
rect 11677 25437 11729 25489
<< metal2 >>
rect 1221 25597 1405 25609
rect 1221 25545 1233 25597
rect 1285 25545 1341 25597
rect 1393 25545 1405 25597
rect 1221 25489 1405 25545
rect 1221 25437 1233 25489
rect 1285 25437 1341 25489
rect 1393 25437 1405 25489
rect 1221 25425 1405 25437
rect 11557 25597 11741 25609
rect 11557 25545 11569 25597
rect 11621 25545 11677 25597
rect 11729 25545 11741 25597
rect 11557 25489 11741 25545
rect 11557 25437 11569 25489
rect 11621 25437 11677 25489
rect 11729 25437 11741 25489
rect 11557 25425 11741 25437
use comp018green_esd_rc_v5p0  comp018green_esd_rc_v5p0_0
timestamp 1758726819
transform 1 0 -356 0 -1 46507
box -51 491 13725 17038
use nmos_clamp_20_50_4  nmos_clamp_20_50_4_0
timestamp 1764277317
transform 1 0 0 0 1 0
box -51 -51 13013 25617
use top_route_1  top_route_1_0
timestamp 1758726819
transform 1 0 43 0 1 25617
box 0 0 12876 21798
<< end >>
