magic
tech gf180mcuD
magscale 1 10
timestamp 1764277680
<< nwell >>
rect 2167 27752 10795 29296
<< hvnmos >>
rect 4129 26006 4269 27006
rect 5191 26006 5331 27006
rect 5435 26006 5575 27006
rect 5679 26006 5819 27006
rect 5923 26006 6063 27006
rect 6167 26006 6307 27006
rect 6411 26006 6551 27006
rect 6655 26006 6795 27006
rect 6899 26006 7039 27006
rect 7143 26006 7283 27006
rect 7387 26006 7527 27006
rect 7631 26006 7771 27006
rect 7875 26006 8015 27006
<< hvpmos >>
rect 2665 27917 2805 28917
rect 2909 27917 3049 28917
rect 3153 27917 3293 28917
rect 3397 27917 3537 28917
rect 3641 27917 3781 28917
rect 3885 27917 4025 28917
rect 4129 27917 4269 28917
rect 4545 27917 4685 28917
rect 4789 27917 4929 28917
rect 5033 27917 5173 28917
rect 5277 27917 5417 28917
rect 5521 27917 5661 28917
rect 5765 27917 5905 28917
rect 6009 27917 6149 28917
rect 6253 27917 6393 28917
rect 6497 27917 6637 28917
rect 6741 27917 6881 28917
rect 6985 27917 7125 28917
rect 7229 27917 7369 28917
rect 7473 27917 7613 28917
rect 7717 27917 7857 28917
rect 7961 27917 8101 28917
rect 8205 27917 8345 28917
rect 8449 27917 8589 28917
rect 8693 27917 8833 28917
rect 8937 27917 9077 28917
rect 9181 27917 9321 28917
rect 9425 27917 9565 28917
rect 9669 27917 9809 28917
rect 9913 27917 10053 28917
rect 10157 27917 10297 28917
<< mvndiff >>
rect 4041 26993 4129 27006
rect 4041 26947 4054 26993
rect 4100 26947 4129 26993
rect 4041 26890 4129 26947
rect 4041 26844 4054 26890
rect 4100 26844 4129 26890
rect 4041 26787 4129 26844
rect 4041 26741 4054 26787
rect 4100 26741 4129 26787
rect 4041 26684 4129 26741
rect 4041 26638 4054 26684
rect 4100 26638 4129 26684
rect 4041 26581 4129 26638
rect 4041 26535 4054 26581
rect 4100 26535 4129 26581
rect 4041 26478 4129 26535
rect 4041 26432 4054 26478
rect 4100 26432 4129 26478
rect 4041 26375 4129 26432
rect 4041 26329 4054 26375
rect 4100 26329 4129 26375
rect 4041 26272 4129 26329
rect 4041 26226 4054 26272
rect 4100 26226 4129 26272
rect 4041 26169 4129 26226
rect 4041 26123 4054 26169
rect 4100 26123 4129 26169
rect 4041 26065 4129 26123
rect 4041 26019 4054 26065
rect 4100 26019 4129 26065
rect 4041 26006 4129 26019
rect 4269 26993 4357 27006
rect 4269 26947 4298 26993
rect 4344 26947 4357 26993
rect 4269 26890 4357 26947
rect 4269 26844 4298 26890
rect 4344 26844 4357 26890
rect 4269 26787 4357 26844
rect 4269 26741 4298 26787
rect 4344 26741 4357 26787
rect 4269 26684 4357 26741
rect 4269 26638 4298 26684
rect 4344 26638 4357 26684
rect 4269 26581 4357 26638
rect 4269 26535 4298 26581
rect 4344 26535 4357 26581
rect 4269 26478 4357 26535
rect 4269 26432 4298 26478
rect 4344 26432 4357 26478
rect 4269 26375 4357 26432
rect 4269 26329 4298 26375
rect 4344 26329 4357 26375
rect 4269 26272 4357 26329
rect 4269 26226 4298 26272
rect 4344 26226 4357 26272
rect 4269 26169 4357 26226
rect 4269 26123 4298 26169
rect 4344 26123 4357 26169
rect 4269 26065 4357 26123
rect 4269 26019 4298 26065
rect 4344 26019 4357 26065
rect 4269 26006 4357 26019
rect 5103 26993 5191 27006
rect 5103 26947 5116 26993
rect 5162 26947 5191 26993
rect 5103 26890 5191 26947
rect 5103 26844 5116 26890
rect 5162 26844 5191 26890
rect 5103 26787 5191 26844
rect 5103 26741 5116 26787
rect 5162 26741 5191 26787
rect 5103 26684 5191 26741
rect 5103 26638 5116 26684
rect 5162 26638 5191 26684
rect 5103 26581 5191 26638
rect 5103 26535 5116 26581
rect 5162 26535 5191 26581
rect 5103 26478 5191 26535
rect 5103 26432 5116 26478
rect 5162 26432 5191 26478
rect 5103 26375 5191 26432
rect 5103 26329 5116 26375
rect 5162 26329 5191 26375
rect 5103 26272 5191 26329
rect 5103 26226 5116 26272
rect 5162 26226 5191 26272
rect 5103 26169 5191 26226
rect 5103 26123 5116 26169
rect 5162 26123 5191 26169
rect 5103 26065 5191 26123
rect 5103 26019 5116 26065
rect 5162 26019 5191 26065
rect 5103 26006 5191 26019
rect 5331 26993 5435 27006
rect 5331 26947 5360 26993
rect 5406 26947 5435 26993
rect 5331 26890 5435 26947
rect 5331 26844 5360 26890
rect 5406 26844 5435 26890
rect 5331 26787 5435 26844
rect 5331 26741 5360 26787
rect 5406 26741 5435 26787
rect 5331 26684 5435 26741
rect 5331 26638 5360 26684
rect 5406 26638 5435 26684
rect 5331 26581 5435 26638
rect 5331 26535 5360 26581
rect 5406 26535 5435 26581
rect 5331 26478 5435 26535
rect 5331 26432 5360 26478
rect 5406 26432 5435 26478
rect 5331 26375 5435 26432
rect 5331 26329 5360 26375
rect 5406 26329 5435 26375
rect 5331 26272 5435 26329
rect 5331 26226 5360 26272
rect 5406 26226 5435 26272
rect 5331 26169 5435 26226
rect 5331 26123 5360 26169
rect 5406 26123 5435 26169
rect 5331 26065 5435 26123
rect 5331 26019 5360 26065
rect 5406 26019 5435 26065
rect 5331 26006 5435 26019
rect 5575 26993 5679 27006
rect 5575 26947 5604 26993
rect 5650 26947 5679 26993
rect 5575 26890 5679 26947
rect 5575 26844 5604 26890
rect 5650 26844 5679 26890
rect 5575 26787 5679 26844
rect 5575 26741 5604 26787
rect 5650 26741 5679 26787
rect 5575 26684 5679 26741
rect 5575 26638 5604 26684
rect 5650 26638 5679 26684
rect 5575 26581 5679 26638
rect 5575 26535 5604 26581
rect 5650 26535 5679 26581
rect 5575 26478 5679 26535
rect 5575 26432 5604 26478
rect 5650 26432 5679 26478
rect 5575 26375 5679 26432
rect 5575 26329 5604 26375
rect 5650 26329 5679 26375
rect 5575 26272 5679 26329
rect 5575 26226 5604 26272
rect 5650 26226 5679 26272
rect 5575 26169 5679 26226
rect 5575 26123 5604 26169
rect 5650 26123 5679 26169
rect 5575 26065 5679 26123
rect 5575 26019 5604 26065
rect 5650 26019 5679 26065
rect 5575 26006 5679 26019
rect 5819 26993 5923 27006
rect 5819 26947 5848 26993
rect 5894 26947 5923 26993
rect 5819 26890 5923 26947
rect 5819 26844 5848 26890
rect 5894 26844 5923 26890
rect 5819 26787 5923 26844
rect 5819 26741 5848 26787
rect 5894 26741 5923 26787
rect 5819 26684 5923 26741
rect 5819 26638 5848 26684
rect 5894 26638 5923 26684
rect 5819 26581 5923 26638
rect 5819 26535 5848 26581
rect 5894 26535 5923 26581
rect 5819 26478 5923 26535
rect 5819 26432 5848 26478
rect 5894 26432 5923 26478
rect 5819 26375 5923 26432
rect 5819 26329 5848 26375
rect 5894 26329 5923 26375
rect 5819 26272 5923 26329
rect 5819 26226 5848 26272
rect 5894 26226 5923 26272
rect 5819 26169 5923 26226
rect 5819 26123 5848 26169
rect 5894 26123 5923 26169
rect 5819 26065 5923 26123
rect 5819 26019 5848 26065
rect 5894 26019 5923 26065
rect 5819 26006 5923 26019
rect 6063 26993 6167 27006
rect 6063 26947 6092 26993
rect 6138 26947 6167 26993
rect 6063 26890 6167 26947
rect 6063 26844 6092 26890
rect 6138 26844 6167 26890
rect 6063 26787 6167 26844
rect 6063 26741 6092 26787
rect 6138 26741 6167 26787
rect 6063 26684 6167 26741
rect 6063 26638 6092 26684
rect 6138 26638 6167 26684
rect 6063 26581 6167 26638
rect 6063 26535 6092 26581
rect 6138 26535 6167 26581
rect 6063 26478 6167 26535
rect 6063 26432 6092 26478
rect 6138 26432 6167 26478
rect 6063 26375 6167 26432
rect 6063 26329 6092 26375
rect 6138 26329 6167 26375
rect 6063 26272 6167 26329
rect 6063 26226 6092 26272
rect 6138 26226 6167 26272
rect 6063 26169 6167 26226
rect 6063 26123 6092 26169
rect 6138 26123 6167 26169
rect 6063 26065 6167 26123
rect 6063 26019 6092 26065
rect 6138 26019 6167 26065
rect 6063 26006 6167 26019
rect 6307 26993 6411 27006
rect 6307 26947 6336 26993
rect 6382 26947 6411 26993
rect 6307 26890 6411 26947
rect 6307 26844 6336 26890
rect 6382 26844 6411 26890
rect 6307 26787 6411 26844
rect 6307 26741 6336 26787
rect 6382 26741 6411 26787
rect 6307 26684 6411 26741
rect 6307 26638 6336 26684
rect 6382 26638 6411 26684
rect 6307 26581 6411 26638
rect 6307 26535 6336 26581
rect 6382 26535 6411 26581
rect 6307 26478 6411 26535
rect 6307 26432 6336 26478
rect 6382 26432 6411 26478
rect 6307 26375 6411 26432
rect 6307 26329 6336 26375
rect 6382 26329 6411 26375
rect 6307 26272 6411 26329
rect 6307 26226 6336 26272
rect 6382 26226 6411 26272
rect 6307 26169 6411 26226
rect 6307 26123 6336 26169
rect 6382 26123 6411 26169
rect 6307 26065 6411 26123
rect 6307 26019 6336 26065
rect 6382 26019 6411 26065
rect 6307 26006 6411 26019
rect 6551 26993 6655 27006
rect 6551 26947 6580 26993
rect 6626 26947 6655 26993
rect 6551 26890 6655 26947
rect 6551 26844 6580 26890
rect 6626 26844 6655 26890
rect 6551 26787 6655 26844
rect 6551 26741 6580 26787
rect 6626 26741 6655 26787
rect 6551 26684 6655 26741
rect 6551 26638 6580 26684
rect 6626 26638 6655 26684
rect 6551 26581 6655 26638
rect 6551 26535 6580 26581
rect 6626 26535 6655 26581
rect 6551 26478 6655 26535
rect 6551 26432 6580 26478
rect 6626 26432 6655 26478
rect 6551 26375 6655 26432
rect 6551 26329 6580 26375
rect 6626 26329 6655 26375
rect 6551 26272 6655 26329
rect 6551 26226 6580 26272
rect 6626 26226 6655 26272
rect 6551 26169 6655 26226
rect 6551 26123 6580 26169
rect 6626 26123 6655 26169
rect 6551 26065 6655 26123
rect 6551 26019 6580 26065
rect 6626 26019 6655 26065
rect 6551 26006 6655 26019
rect 6795 26993 6899 27006
rect 6795 26947 6824 26993
rect 6870 26947 6899 26993
rect 6795 26890 6899 26947
rect 6795 26844 6824 26890
rect 6870 26844 6899 26890
rect 6795 26787 6899 26844
rect 6795 26741 6824 26787
rect 6870 26741 6899 26787
rect 6795 26684 6899 26741
rect 6795 26638 6824 26684
rect 6870 26638 6899 26684
rect 6795 26581 6899 26638
rect 6795 26535 6824 26581
rect 6870 26535 6899 26581
rect 6795 26478 6899 26535
rect 6795 26432 6824 26478
rect 6870 26432 6899 26478
rect 6795 26375 6899 26432
rect 6795 26329 6824 26375
rect 6870 26329 6899 26375
rect 6795 26272 6899 26329
rect 6795 26226 6824 26272
rect 6870 26226 6899 26272
rect 6795 26169 6899 26226
rect 6795 26123 6824 26169
rect 6870 26123 6899 26169
rect 6795 26065 6899 26123
rect 6795 26019 6824 26065
rect 6870 26019 6899 26065
rect 6795 26006 6899 26019
rect 7039 26993 7143 27006
rect 7039 26947 7068 26993
rect 7114 26947 7143 26993
rect 7039 26890 7143 26947
rect 7039 26844 7068 26890
rect 7114 26844 7143 26890
rect 7039 26787 7143 26844
rect 7039 26741 7068 26787
rect 7114 26741 7143 26787
rect 7039 26684 7143 26741
rect 7039 26638 7068 26684
rect 7114 26638 7143 26684
rect 7039 26581 7143 26638
rect 7039 26535 7068 26581
rect 7114 26535 7143 26581
rect 7039 26478 7143 26535
rect 7039 26432 7068 26478
rect 7114 26432 7143 26478
rect 7039 26375 7143 26432
rect 7039 26329 7068 26375
rect 7114 26329 7143 26375
rect 7039 26272 7143 26329
rect 7039 26226 7068 26272
rect 7114 26226 7143 26272
rect 7039 26169 7143 26226
rect 7039 26123 7068 26169
rect 7114 26123 7143 26169
rect 7039 26065 7143 26123
rect 7039 26019 7068 26065
rect 7114 26019 7143 26065
rect 7039 26006 7143 26019
rect 7283 26993 7387 27006
rect 7283 26947 7312 26993
rect 7358 26947 7387 26993
rect 7283 26890 7387 26947
rect 7283 26844 7312 26890
rect 7358 26844 7387 26890
rect 7283 26787 7387 26844
rect 7283 26741 7312 26787
rect 7358 26741 7387 26787
rect 7283 26684 7387 26741
rect 7283 26638 7312 26684
rect 7358 26638 7387 26684
rect 7283 26581 7387 26638
rect 7283 26535 7312 26581
rect 7358 26535 7387 26581
rect 7283 26478 7387 26535
rect 7283 26432 7312 26478
rect 7358 26432 7387 26478
rect 7283 26375 7387 26432
rect 7283 26329 7312 26375
rect 7358 26329 7387 26375
rect 7283 26272 7387 26329
rect 7283 26226 7312 26272
rect 7358 26226 7387 26272
rect 7283 26169 7387 26226
rect 7283 26123 7312 26169
rect 7358 26123 7387 26169
rect 7283 26065 7387 26123
rect 7283 26019 7312 26065
rect 7358 26019 7387 26065
rect 7283 26006 7387 26019
rect 7527 26993 7631 27006
rect 7527 26947 7556 26993
rect 7602 26947 7631 26993
rect 7527 26890 7631 26947
rect 7527 26844 7556 26890
rect 7602 26844 7631 26890
rect 7527 26787 7631 26844
rect 7527 26741 7556 26787
rect 7602 26741 7631 26787
rect 7527 26684 7631 26741
rect 7527 26638 7556 26684
rect 7602 26638 7631 26684
rect 7527 26581 7631 26638
rect 7527 26535 7556 26581
rect 7602 26535 7631 26581
rect 7527 26478 7631 26535
rect 7527 26432 7556 26478
rect 7602 26432 7631 26478
rect 7527 26375 7631 26432
rect 7527 26329 7556 26375
rect 7602 26329 7631 26375
rect 7527 26272 7631 26329
rect 7527 26226 7556 26272
rect 7602 26226 7631 26272
rect 7527 26169 7631 26226
rect 7527 26123 7556 26169
rect 7602 26123 7631 26169
rect 7527 26065 7631 26123
rect 7527 26019 7556 26065
rect 7602 26019 7631 26065
rect 7527 26006 7631 26019
rect 7771 26993 7875 27006
rect 7771 26947 7800 26993
rect 7846 26947 7875 26993
rect 7771 26890 7875 26947
rect 7771 26844 7800 26890
rect 7846 26844 7875 26890
rect 7771 26787 7875 26844
rect 7771 26741 7800 26787
rect 7846 26741 7875 26787
rect 7771 26684 7875 26741
rect 7771 26638 7800 26684
rect 7846 26638 7875 26684
rect 7771 26581 7875 26638
rect 7771 26535 7800 26581
rect 7846 26535 7875 26581
rect 7771 26478 7875 26535
rect 7771 26432 7800 26478
rect 7846 26432 7875 26478
rect 7771 26375 7875 26432
rect 7771 26329 7800 26375
rect 7846 26329 7875 26375
rect 7771 26272 7875 26329
rect 7771 26226 7800 26272
rect 7846 26226 7875 26272
rect 7771 26169 7875 26226
rect 7771 26123 7800 26169
rect 7846 26123 7875 26169
rect 7771 26065 7875 26123
rect 7771 26019 7800 26065
rect 7846 26019 7875 26065
rect 7771 26006 7875 26019
rect 8015 26993 8103 27006
rect 8015 26947 8044 26993
rect 8090 26947 8103 26993
rect 8015 26890 8103 26947
rect 8015 26844 8044 26890
rect 8090 26844 8103 26890
rect 8015 26787 8103 26844
rect 8015 26741 8044 26787
rect 8090 26741 8103 26787
rect 8015 26684 8103 26741
rect 8015 26638 8044 26684
rect 8090 26638 8103 26684
rect 8015 26581 8103 26638
rect 8015 26535 8044 26581
rect 8090 26535 8103 26581
rect 8015 26478 8103 26535
rect 8015 26432 8044 26478
rect 8090 26432 8103 26478
rect 8015 26375 8103 26432
rect 8015 26329 8044 26375
rect 8090 26329 8103 26375
rect 8015 26272 8103 26329
rect 8015 26226 8044 26272
rect 8090 26226 8103 26272
rect 8015 26169 8103 26226
rect 8015 26123 8044 26169
rect 8090 26123 8103 26169
rect 8015 26065 8103 26123
rect 8015 26019 8044 26065
rect 8090 26019 8103 26065
rect 8015 26006 8103 26019
<< mvpdiff >>
rect 2577 28904 2665 28917
rect 2577 28858 2590 28904
rect 2636 28858 2665 28904
rect 2577 28801 2665 28858
rect 2577 28755 2590 28801
rect 2636 28755 2665 28801
rect 2577 28698 2665 28755
rect 2577 28652 2590 28698
rect 2636 28652 2665 28698
rect 2577 28595 2665 28652
rect 2577 28549 2590 28595
rect 2636 28549 2665 28595
rect 2577 28492 2665 28549
rect 2577 28446 2590 28492
rect 2636 28446 2665 28492
rect 2577 28389 2665 28446
rect 2577 28343 2590 28389
rect 2636 28343 2665 28389
rect 2577 28286 2665 28343
rect 2577 28240 2590 28286
rect 2636 28240 2665 28286
rect 2577 28183 2665 28240
rect 2577 28137 2590 28183
rect 2636 28137 2665 28183
rect 2577 28080 2665 28137
rect 2577 28034 2590 28080
rect 2636 28034 2665 28080
rect 2577 27976 2665 28034
rect 2577 27930 2590 27976
rect 2636 27930 2665 27976
rect 2577 27917 2665 27930
rect 2805 28904 2909 28917
rect 2805 28858 2834 28904
rect 2880 28858 2909 28904
rect 2805 28801 2909 28858
rect 2805 28755 2834 28801
rect 2880 28755 2909 28801
rect 2805 28698 2909 28755
rect 2805 28652 2834 28698
rect 2880 28652 2909 28698
rect 2805 28595 2909 28652
rect 2805 28549 2834 28595
rect 2880 28549 2909 28595
rect 2805 28492 2909 28549
rect 2805 28446 2834 28492
rect 2880 28446 2909 28492
rect 2805 28389 2909 28446
rect 2805 28343 2834 28389
rect 2880 28343 2909 28389
rect 2805 28286 2909 28343
rect 2805 28240 2834 28286
rect 2880 28240 2909 28286
rect 2805 28183 2909 28240
rect 2805 28137 2834 28183
rect 2880 28137 2909 28183
rect 2805 28080 2909 28137
rect 2805 28034 2834 28080
rect 2880 28034 2909 28080
rect 2805 27976 2909 28034
rect 2805 27930 2834 27976
rect 2880 27930 2909 27976
rect 2805 27917 2909 27930
rect 3049 28904 3153 28917
rect 3049 28858 3078 28904
rect 3124 28858 3153 28904
rect 3049 28801 3153 28858
rect 3049 28755 3078 28801
rect 3124 28755 3153 28801
rect 3049 28698 3153 28755
rect 3049 28652 3078 28698
rect 3124 28652 3153 28698
rect 3049 28595 3153 28652
rect 3049 28549 3078 28595
rect 3124 28549 3153 28595
rect 3049 28492 3153 28549
rect 3049 28446 3078 28492
rect 3124 28446 3153 28492
rect 3049 28389 3153 28446
rect 3049 28343 3078 28389
rect 3124 28343 3153 28389
rect 3049 28286 3153 28343
rect 3049 28240 3078 28286
rect 3124 28240 3153 28286
rect 3049 28183 3153 28240
rect 3049 28137 3078 28183
rect 3124 28137 3153 28183
rect 3049 28080 3153 28137
rect 3049 28034 3078 28080
rect 3124 28034 3153 28080
rect 3049 27976 3153 28034
rect 3049 27930 3078 27976
rect 3124 27930 3153 27976
rect 3049 27917 3153 27930
rect 3293 28904 3397 28917
rect 3293 28858 3322 28904
rect 3368 28858 3397 28904
rect 3293 28801 3397 28858
rect 3293 28755 3322 28801
rect 3368 28755 3397 28801
rect 3293 28698 3397 28755
rect 3293 28652 3322 28698
rect 3368 28652 3397 28698
rect 3293 28595 3397 28652
rect 3293 28549 3322 28595
rect 3368 28549 3397 28595
rect 3293 28492 3397 28549
rect 3293 28446 3322 28492
rect 3368 28446 3397 28492
rect 3293 28389 3397 28446
rect 3293 28343 3322 28389
rect 3368 28343 3397 28389
rect 3293 28286 3397 28343
rect 3293 28240 3322 28286
rect 3368 28240 3397 28286
rect 3293 28183 3397 28240
rect 3293 28137 3322 28183
rect 3368 28137 3397 28183
rect 3293 28080 3397 28137
rect 3293 28034 3322 28080
rect 3368 28034 3397 28080
rect 3293 27976 3397 28034
rect 3293 27930 3322 27976
rect 3368 27930 3397 27976
rect 3293 27917 3397 27930
rect 3537 28904 3641 28917
rect 3537 28858 3566 28904
rect 3612 28858 3641 28904
rect 3537 28801 3641 28858
rect 3537 28755 3566 28801
rect 3612 28755 3641 28801
rect 3537 28698 3641 28755
rect 3537 28652 3566 28698
rect 3612 28652 3641 28698
rect 3537 28595 3641 28652
rect 3537 28549 3566 28595
rect 3612 28549 3641 28595
rect 3537 28492 3641 28549
rect 3537 28446 3566 28492
rect 3612 28446 3641 28492
rect 3537 28389 3641 28446
rect 3537 28343 3566 28389
rect 3612 28343 3641 28389
rect 3537 28286 3641 28343
rect 3537 28240 3566 28286
rect 3612 28240 3641 28286
rect 3537 28183 3641 28240
rect 3537 28137 3566 28183
rect 3612 28137 3641 28183
rect 3537 28080 3641 28137
rect 3537 28034 3566 28080
rect 3612 28034 3641 28080
rect 3537 27976 3641 28034
rect 3537 27930 3566 27976
rect 3612 27930 3641 27976
rect 3537 27917 3641 27930
rect 3781 28904 3885 28917
rect 3781 28858 3810 28904
rect 3856 28858 3885 28904
rect 3781 28801 3885 28858
rect 3781 28755 3810 28801
rect 3856 28755 3885 28801
rect 3781 28698 3885 28755
rect 3781 28652 3810 28698
rect 3856 28652 3885 28698
rect 3781 28595 3885 28652
rect 3781 28549 3810 28595
rect 3856 28549 3885 28595
rect 3781 28492 3885 28549
rect 3781 28446 3810 28492
rect 3856 28446 3885 28492
rect 3781 28389 3885 28446
rect 3781 28343 3810 28389
rect 3856 28343 3885 28389
rect 3781 28286 3885 28343
rect 3781 28240 3810 28286
rect 3856 28240 3885 28286
rect 3781 28183 3885 28240
rect 3781 28137 3810 28183
rect 3856 28137 3885 28183
rect 3781 28080 3885 28137
rect 3781 28034 3810 28080
rect 3856 28034 3885 28080
rect 3781 27976 3885 28034
rect 3781 27930 3810 27976
rect 3856 27930 3885 27976
rect 3781 27917 3885 27930
rect 4025 28904 4129 28917
rect 4025 28858 4054 28904
rect 4100 28858 4129 28904
rect 4025 28801 4129 28858
rect 4025 28755 4054 28801
rect 4100 28755 4129 28801
rect 4025 28698 4129 28755
rect 4025 28652 4054 28698
rect 4100 28652 4129 28698
rect 4025 28595 4129 28652
rect 4025 28549 4054 28595
rect 4100 28549 4129 28595
rect 4025 28492 4129 28549
rect 4025 28446 4054 28492
rect 4100 28446 4129 28492
rect 4025 28389 4129 28446
rect 4025 28343 4054 28389
rect 4100 28343 4129 28389
rect 4025 28286 4129 28343
rect 4025 28240 4054 28286
rect 4100 28240 4129 28286
rect 4025 28183 4129 28240
rect 4025 28137 4054 28183
rect 4100 28137 4129 28183
rect 4025 28080 4129 28137
rect 4025 28034 4054 28080
rect 4100 28034 4129 28080
rect 4025 27976 4129 28034
rect 4025 27930 4054 27976
rect 4100 27930 4129 27976
rect 4025 27917 4129 27930
rect 4269 28904 4357 28917
rect 4269 28858 4298 28904
rect 4344 28858 4357 28904
rect 4269 28801 4357 28858
rect 4269 28755 4298 28801
rect 4344 28755 4357 28801
rect 4269 28698 4357 28755
rect 4269 28652 4298 28698
rect 4344 28652 4357 28698
rect 4269 28595 4357 28652
rect 4269 28549 4298 28595
rect 4344 28549 4357 28595
rect 4269 28492 4357 28549
rect 4269 28446 4298 28492
rect 4344 28446 4357 28492
rect 4269 28389 4357 28446
rect 4269 28343 4298 28389
rect 4344 28343 4357 28389
rect 4269 28286 4357 28343
rect 4269 28240 4298 28286
rect 4344 28240 4357 28286
rect 4269 28183 4357 28240
rect 4269 28137 4298 28183
rect 4344 28137 4357 28183
rect 4269 28080 4357 28137
rect 4269 28034 4298 28080
rect 4344 28034 4357 28080
rect 4269 27976 4357 28034
rect 4269 27930 4298 27976
rect 4344 27930 4357 27976
rect 4269 27917 4357 27930
rect 4457 28904 4545 28917
rect 4457 28858 4470 28904
rect 4516 28858 4545 28904
rect 4457 28801 4545 28858
rect 4457 28755 4470 28801
rect 4516 28755 4545 28801
rect 4457 28698 4545 28755
rect 4457 28652 4470 28698
rect 4516 28652 4545 28698
rect 4457 28595 4545 28652
rect 4457 28549 4470 28595
rect 4516 28549 4545 28595
rect 4457 28492 4545 28549
rect 4457 28446 4470 28492
rect 4516 28446 4545 28492
rect 4457 28389 4545 28446
rect 4457 28343 4470 28389
rect 4516 28343 4545 28389
rect 4457 28286 4545 28343
rect 4457 28240 4470 28286
rect 4516 28240 4545 28286
rect 4457 28183 4545 28240
rect 4457 28137 4470 28183
rect 4516 28137 4545 28183
rect 4457 28080 4545 28137
rect 4457 28034 4470 28080
rect 4516 28034 4545 28080
rect 4457 27976 4545 28034
rect 4457 27930 4470 27976
rect 4516 27930 4545 27976
rect 4457 27917 4545 27930
rect 4685 28904 4789 28917
rect 4685 28858 4714 28904
rect 4760 28858 4789 28904
rect 4685 28801 4789 28858
rect 4685 28755 4714 28801
rect 4760 28755 4789 28801
rect 4685 28698 4789 28755
rect 4685 28652 4714 28698
rect 4760 28652 4789 28698
rect 4685 28595 4789 28652
rect 4685 28549 4714 28595
rect 4760 28549 4789 28595
rect 4685 28492 4789 28549
rect 4685 28446 4714 28492
rect 4760 28446 4789 28492
rect 4685 28389 4789 28446
rect 4685 28343 4714 28389
rect 4760 28343 4789 28389
rect 4685 28286 4789 28343
rect 4685 28240 4714 28286
rect 4760 28240 4789 28286
rect 4685 28183 4789 28240
rect 4685 28137 4714 28183
rect 4760 28137 4789 28183
rect 4685 28080 4789 28137
rect 4685 28034 4714 28080
rect 4760 28034 4789 28080
rect 4685 27976 4789 28034
rect 4685 27930 4714 27976
rect 4760 27930 4789 27976
rect 4685 27917 4789 27930
rect 4929 28904 5033 28917
rect 4929 28858 4958 28904
rect 5004 28858 5033 28904
rect 4929 28801 5033 28858
rect 4929 28755 4958 28801
rect 5004 28755 5033 28801
rect 4929 28698 5033 28755
rect 4929 28652 4958 28698
rect 5004 28652 5033 28698
rect 4929 28595 5033 28652
rect 4929 28549 4958 28595
rect 5004 28549 5033 28595
rect 4929 28492 5033 28549
rect 4929 28446 4958 28492
rect 5004 28446 5033 28492
rect 4929 28389 5033 28446
rect 4929 28343 4958 28389
rect 5004 28343 5033 28389
rect 4929 28286 5033 28343
rect 4929 28240 4958 28286
rect 5004 28240 5033 28286
rect 4929 28183 5033 28240
rect 4929 28137 4958 28183
rect 5004 28137 5033 28183
rect 4929 28080 5033 28137
rect 4929 28034 4958 28080
rect 5004 28034 5033 28080
rect 4929 27976 5033 28034
rect 4929 27930 4958 27976
rect 5004 27930 5033 27976
rect 4929 27917 5033 27930
rect 5173 28904 5277 28917
rect 5173 28858 5202 28904
rect 5248 28858 5277 28904
rect 5173 28801 5277 28858
rect 5173 28755 5202 28801
rect 5248 28755 5277 28801
rect 5173 28698 5277 28755
rect 5173 28652 5202 28698
rect 5248 28652 5277 28698
rect 5173 28595 5277 28652
rect 5173 28549 5202 28595
rect 5248 28549 5277 28595
rect 5173 28492 5277 28549
rect 5173 28446 5202 28492
rect 5248 28446 5277 28492
rect 5173 28389 5277 28446
rect 5173 28343 5202 28389
rect 5248 28343 5277 28389
rect 5173 28286 5277 28343
rect 5173 28240 5202 28286
rect 5248 28240 5277 28286
rect 5173 28183 5277 28240
rect 5173 28137 5202 28183
rect 5248 28137 5277 28183
rect 5173 28080 5277 28137
rect 5173 28034 5202 28080
rect 5248 28034 5277 28080
rect 5173 27976 5277 28034
rect 5173 27930 5202 27976
rect 5248 27930 5277 27976
rect 5173 27917 5277 27930
rect 5417 28904 5521 28917
rect 5417 28858 5446 28904
rect 5492 28858 5521 28904
rect 5417 28801 5521 28858
rect 5417 28755 5446 28801
rect 5492 28755 5521 28801
rect 5417 28698 5521 28755
rect 5417 28652 5446 28698
rect 5492 28652 5521 28698
rect 5417 28595 5521 28652
rect 5417 28549 5446 28595
rect 5492 28549 5521 28595
rect 5417 28492 5521 28549
rect 5417 28446 5446 28492
rect 5492 28446 5521 28492
rect 5417 28389 5521 28446
rect 5417 28343 5446 28389
rect 5492 28343 5521 28389
rect 5417 28286 5521 28343
rect 5417 28240 5446 28286
rect 5492 28240 5521 28286
rect 5417 28183 5521 28240
rect 5417 28137 5446 28183
rect 5492 28137 5521 28183
rect 5417 28080 5521 28137
rect 5417 28034 5446 28080
rect 5492 28034 5521 28080
rect 5417 27976 5521 28034
rect 5417 27930 5446 27976
rect 5492 27930 5521 27976
rect 5417 27917 5521 27930
rect 5661 28904 5765 28917
rect 5661 28858 5690 28904
rect 5736 28858 5765 28904
rect 5661 28801 5765 28858
rect 5661 28755 5690 28801
rect 5736 28755 5765 28801
rect 5661 28698 5765 28755
rect 5661 28652 5690 28698
rect 5736 28652 5765 28698
rect 5661 28595 5765 28652
rect 5661 28549 5690 28595
rect 5736 28549 5765 28595
rect 5661 28492 5765 28549
rect 5661 28446 5690 28492
rect 5736 28446 5765 28492
rect 5661 28389 5765 28446
rect 5661 28343 5690 28389
rect 5736 28343 5765 28389
rect 5661 28286 5765 28343
rect 5661 28240 5690 28286
rect 5736 28240 5765 28286
rect 5661 28183 5765 28240
rect 5661 28137 5690 28183
rect 5736 28137 5765 28183
rect 5661 28080 5765 28137
rect 5661 28034 5690 28080
rect 5736 28034 5765 28080
rect 5661 27976 5765 28034
rect 5661 27930 5690 27976
rect 5736 27930 5765 27976
rect 5661 27917 5765 27930
rect 5905 28904 6009 28917
rect 5905 28858 5934 28904
rect 5980 28858 6009 28904
rect 5905 28801 6009 28858
rect 5905 28755 5934 28801
rect 5980 28755 6009 28801
rect 5905 28698 6009 28755
rect 5905 28652 5934 28698
rect 5980 28652 6009 28698
rect 5905 28595 6009 28652
rect 5905 28549 5934 28595
rect 5980 28549 6009 28595
rect 5905 28492 6009 28549
rect 5905 28446 5934 28492
rect 5980 28446 6009 28492
rect 5905 28389 6009 28446
rect 5905 28343 5934 28389
rect 5980 28343 6009 28389
rect 5905 28286 6009 28343
rect 5905 28240 5934 28286
rect 5980 28240 6009 28286
rect 5905 28183 6009 28240
rect 5905 28137 5934 28183
rect 5980 28137 6009 28183
rect 5905 28080 6009 28137
rect 5905 28034 5934 28080
rect 5980 28034 6009 28080
rect 5905 27976 6009 28034
rect 5905 27930 5934 27976
rect 5980 27930 6009 27976
rect 5905 27917 6009 27930
rect 6149 28904 6253 28917
rect 6149 28858 6178 28904
rect 6224 28858 6253 28904
rect 6149 28801 6253 28858
rect 6149 28755 6178 28801
rect 6224 28755 6253 28801
rect 6149 28698 6253 28755
rect 6149 28652 6178 28698
rect 6224 28652 6253 28698
rect 6149 28595 6253 28652
rect 6149 28549 6178 28595
rect 6224 28549 6253 28595
rect 6149 28492 6253 28549
rect 6149 28446 6178 28492
rect 6224 28446 6253 28492
rect 6149 28389 6253 28446
rect 6149 28343 6178 28389
rect 6224 28343 6253 28389
rect 6149 28286 6253 28343
rect 6149 28240 6178 28286
rect 6224 28240 6253 28286
rect 6149 28183 6253 28240
rect 6149 28137 6178 28183
rect 6224 28137 6253 28183
rect 6149 28080 6253 28137
rect 6149 28034 6178 28080
rect 6224 28034 6253 28080
rect 6149 27976 6253 28034
rect 6149 27930 6178 27976
rect 6224 27930 6253 27976
rect 6149 27917 6253 27930
rect 6393 28904 6497 28917
rect 6393 28858 6422 28904
rect 6468 28858 6497 28904
rect 6393 28801 6497 28858
rect 6393 28755 6422 28801
rect 6468 28755 6497 28801
rect 6393 28698 6497 28755
rect 6393 28652 6422 28698
rect 6468 28652 6497 28698
rect 6393 28595 6497 28652
rect 6393 28549 6422 28595
rect 6468 28549 6497 28595
rect 6393 28492 6497 28549
rect 6393 28446 6422 28492
rect 6468 28446 6497 28492
rect 6393 28389 6497 28446
rect 6393 28343 6422 28389
rect 6468 28343 6497 28389
rect 6393 28286 6497 28343
rect 6393 28240 6422 28286
rect 6468 28240 6497 28286
rect 6393 28183 6497 28240
rect 6393 28137 6422 28183
rect 6468 28137 6497 28183
rect 6393 28080 6497 28137
rect 6393 28034 6422 28080
rect 6468 28034 6497 28080
rect 6393 27976 6497 28034
rect 6393 27930 6422 27976
rect 6468 27930 6497 27976
rect 6393 27917 6497 27930
rect 6637 28904 6741 28917
rect 6637 28858 6666 28904
rect 6712 28858 6741 28904
rect 6637 28801 6741 28858
rect 6637 28755 6666 28801
rect 6712 28755 6741 28801
rect 6637 28698 6741 28755
rect 6637 28652 6666 28698
rect 6712 28652 6741 28698
rect 6637 28595 6741 28652
rect 6637 28549 6666 28595
rect 6712 28549 6741 28595
rect 6637 28492 6741 28549
rect 6637 28446 6666 28492
rect 6712 28446 6741 28492
rect 6637 28389 6741 28446
rect 6637 28343 6666 28389
rect 6712 28343 6741 28389
rect 6637 28286 6741 28343
rect 6637 28240 6666 28286
rect 6712 28240 6741 28286
rect 6637 28183 6741 28240
rect 6637 28137 6666 28183
rect 6712 28137 6741 28183
rect 6637 28080 6741 28137
rect 6637 28034 6666 28080
rect 6712 28034 6741 28080
rect 6637 27976 6741 28034
rect 6637 27930 6666 27976
rect 6712 27930 6741 27976
rect 6637 27917 6741 27930
rect 6881 28904 6985 28917
rect 6881 28858 6910 28904
rect 6956 28858 6985 28904
rect 6881 28801 6985 28858
rect 6881 28755 6910 28801
rect 6956 28755 6985 28801
rect 6881 28698 6985 28755
rect 6881 28652 6910 28698
rect 6956 28652 6985 28698
rect 6881 28595 6985 28652
rect 6881 28549 6910 28595
rect 6956 28549 6985 28595
rect 6881 28492 6985 28549
rect 6881 28446 6910 28492
rect 6956 28446 6985 28492
rect 6881 28389 6985 28446
rect 6881 28343 6910 28389
rect 6956 28343 6985 28389
rect 6881 28286 6985 28343
rect 6881 28240 6910 28286
rect 6956 28240 6985 28286
rect 6881 28183 6985 28240
rect 6881 28137 6910 28183
rect 6956 28137 6985 28183
rect 6881 28080 6985 28137
rect 6881 28034 6910 28080
rect 6956 28034 6985 28080
rect 6881 27976 6985 28034
rect 6881 27930 6910 27976
rect 6956 27930 6985 27976
rect 6881 27917 6985 27930
rect 7125 28904 7229 28917
rect 7125 28858 7154 28904
rect 7200 28858 7229 28904
rect 7125 28801 7229 28858
rect 7125 28755 7154 28801
rect 7200 28755 7229 28801
rect 7125 28698 7229 28755
rect 7125 28652 7154 28698
rect 7200 28652 7229 28698
rect 7125 28595 7229 28652
rect 7125 28549 7154 28595
rect 7200 28549 7229 28595
rect 7125 28492 7229 28549
rect 7125 28446 7154 28492
rect 7200 28446 7229 28492
rect 7125 28389 7229 28446
rect 7125 28343 7154 28389
rect 7200 28343 7229 28389
rect 7125 28286 7229 28343
rect 7125 28240 7154 28286
rect 7200 28240 7229 28286
rect 7125 28183 7229 28240
rect 7125 28137 7154 28183
rect 7200 28137 7229 28183
rect 7125 28080 7229 28137
rect 7125 28034 7154 28080
rect 7200 28034 7229 28080
rect 7125 27976 7229 28034
rect 7125 27930 7154 27976
rect 7200 27930 7229 27976
rect 7125 27917 7229 27930
rect 7369 28904 7473 28917
rect 7369 28858 7398 28904
rect 7444 28858 7473 28904
rect 7369 28801 7473 28858
rect 7369 28755 7398 28801
rect 7444 28755 7473 28801
rect 7369 28698 7473 28755
rect 7369 28652 7398 28698
rect 7444 28652 7473 28698
rect 7369 28595 7473 28652
rect 7369 28549 7398 28595
rect 7444 28549 7473 28595
rect 7369 28492 7473 28549
rect 7369 28446 7398 28492
rect 7444 28446 7473 28492
rect 7369 28389 7473 28446
rect 7369 28343 7398 28389
rect 7444 28343 7473 28389
rect 7369 28286 7473 28343
rect 7369 28240 7398 28286
rect 7444 28240 7473 28286
rect 7369 28183 7473 28240
rect 7369 28137 7398 28183
rect 7444 28137 7473 28183
rect 7369 28080 7473 28137
rect 7369 28034 7398 28080
rect 7444 28034 7473 28080
rect 7369 27976 7473 28034
rect 7369 27930 7398 27976
rect 7444 27930 7473 27976
rect 7369 27917 7473 27930
rect 7613 28904 7717 28917
rect 7613 28858 7642 28904
rect 7688 28858 7717 28904
rect 7613 28801 7717 28858
rect 7613 28755 7642 28801
rect 7688 28755 7717 28801
rect 7613 28698 7717 28755
rect 7613 28652 7642 28698
rect 7688 28652 7717 28698
rect 7613 28595 7717 28652
rect 7613 28549 7642 28595
rect 7688 28549 7717 28595
rect 7613 28492 7717 28549
rect 7613 28446 7642 28492
rect 7688 28446 7717 28492
rect 7613 28389 7717 28446
rect 7613 28343 7642 28389
rect 7688 28343 7717 28389
rect 7613 28286 7717 28343
rect 7613 28240 7642 28286
rect 7688 28240 7717 28286
rect 7613 28183 7717 28240
rect 7613 28137 7642 28183
rect 7688 28137 7717 28183
rect 7613 28080 7717 28137
rect 7613 28034 7642 28080
rect 7688 28034 7717 28080
rect 7613 27976 7717 28034
rect 7613 27930 7642 27976
rect 7688 27930 7717 27976
rect 7613 27917 7717 27930
rect 7857 28904 7961 28917
rect 7857 28858 7886 28904
rect 7932 28858 7961 28904
rect 7857 28801 7961 28858
rect 7857 28755 7886 28801
rect 7932 28755 7961 28801
rect 7857 28698 7961 28755
rect 7857 28652 7886 28698
rect 7932 28652 7961 28698
rect 7857 28595 7961 28652
rect 7857 28549 7886 28595
rect 7932 28549 7961 28595
rect 7857 28492 7961 28549
rect 7857 28446 7886 28492
rect 7932 28446 7961 28492
rect 7857 28389 7961 28446
rect 7857 28343 7886 28389
rect 7932 28343 7961 28389
rect 7857 28286 7961 28343
rect 7857 28240 7886 28286
rect 7932 28240 7961 28286
rect 7857 28183 7961 28240
rect 7857 28137 7886 28183
rect 7932 28137 7961 28183
rect 7857 28080 7961 28137
rect 7857 28034 7886 28080
rect 7932 28034 7961 28080
rect 7857 27976 7961 28034
rect 7857 27930 7886 27976
rect 7932 27930 7961 27976
rect 7857 27917 7961 27930
rect 8101 28904 8205 28917
rect 8101 28858 8130 28904
rect 8176 28858 8205 28904
rect 8101 28801 8205 28858
rect 8101 28755 8130 28801
rect 8176 28755 8205 28801
rect 8101 28698 8205 28755
rect 8101 28652 8130 28698
rect 8176 28652 8205 28698
rect 8101 28595 8205 28652
rect 8101 28549 8130 28595
rect 8176 28549 8205 28595
rect 8101 28492 8205 28549
rect 8101 28446 8130 28492
rect 8176 28446 8205 28492
rect 8101 28389 8205 28446
rect 8101 28343 8130 28389
rect 8176 28343 8205 28389
rect 8101 28286 8205 28343
rect 8101 28240 8130 28286
rect 8176 28240 8205 28286
rect 8101 28183 8205 28240
rect 8101 28137 8130 28183
rect 8176 28137 8205 28183
rect 8101 28080 8205 28137
rect 8101 28034 8130 28080
rect 8176 28034 8205 28080
rect 8101 27976 8205 28034
rect 8101 27930 8130 27976
rect 8176 27930 8205 27976
rect 8101 27917 8205 27930
rect 8345 28904 8449 28917
rect 8345 28858 8374 28904
rect 8420 28858 8449 28904
rect 8345 28801 8449 28858
rect 8345 28755 8374 28801
rect 8420 28755 8449 28801
rect 8345 28698 8449 28755
rect 8345 28652 8374 28698
rect 8420 28652 8449 28698
rect 8345 28595 8449 28652
rect 8345 28549 8374 28595
rect 8420 28549 8449 28595
rect 8345 28492 8449 28549
rect 8345 28446 8374 28492
rect 8420 28446 8449 28492
rect 8345 28389 8449 28446
rect 8345 28343 8374 28389
rect 8420 28343 8449 28389
rect 8345 28286 8449 28343
rect 8345 28240 8374 28286
rect 8420 28240 8449 28286
rect 8345 28183 8449 28240
rect 8345 28137 8374 28183
rect 8420 28137 8449 28183
rect 8345 28080 8449 28137
rect 8345 28034 8374 28080
rect 8420 28034 8449 28080
rect 8345 27976 8449 28034
rect 8345 27930 8374 27976
rect 8420 27930 8449 27976
rect 8345 27917 8449 27930
rect 8589 28904 8693 28917
rect 8589 28858 8618 28904
rect 8664 28858 8693 28904
rect 8589 28801 8693 28858
rect 8589 28755 8618 28801
rect 8664 28755 8693 28801
rect 8589 28698 8693 28755
rect 8589 28652 8618 28698
rect 8664 28652 8693 28698
rect 8589 28595 8693 28652
rect 8589 28549 8618 28595
rect 8664 28549 8693 28595
rect 8589 28492 8693 28549
rect 8589 28446 8618 28492
rect 8664 28446 8693 28492
rect 8589 28389 8693 28446
rect 8589 28343 8618 28389
rect 8664 28343 8693 28389
rect 8589 28286 8693 28343
rect 8589 28240 8618 28286
rect 8664 28240 8693 28286
rect 8589 28183 8693 28240
rect 8589 28137 8618 28183
rect 8664 28137 8693 28183
rect 8589 28080 8693 28137
rect 8589 28034 8618 28080
rect 8664 28034 8693 28080
rect 8589 27976 8693 28034
rect 8589 27930 8618 27976
rect 8664 27930 8693 27976
rect 8589 27917 8693 27930
rect 8833 28904 8937 28917
rect 8833 28858 8862 28904
rect 8908 28858 8937 28904
rect 8833 28801 8937 28858
rect 8833 28755 8862 28801
rect 8908 28755 8937 28801
rect 8833 28698 8937 28755
rect 8833 28652 8862 28698
rect 8908 28652 8937 28698
rect 8833 28595 8937 28652
rect 8833 28549 8862 28595
rect 8908 28549 8937 28595
rect 8833 28492 8937 28549
rect 8833 28446 8862 28492
rect 8908 28446 8937 28492
rect 8833 28389 8937 28446
rect 8833 28343 8862 28389
rect 8908 28343 8937 28389
rect 8833 28286 8937 28343
rect 8833 28240 8862 28286
rect 8908 28240 8937 28286
rect 8833 28183 8937 28240
rect 8833 28137 8862 28183
rect 8908 28137 8937 28183
rect 8833 28080 8937 28137
rect 8833 28034 8862 28080
rect 8908 28034 8937 28080
rect 8833 27976 8937 28034
rect 8833 27930 8862 27976
rect 8908 27930 8937 27976
rect 8833 27917 8937 27930
rect 9077 28904 9181 28917
rect 9077 28858 9106 28904
rect 9152 28858 9181 28904
rect 9077 28801 9181 28858
rect 9077 28755 9106 28801
rect 9152 28755 9181 28801
rect 9077 28698 9181 28755
rect 9077 28652 9106 28698
rect 9152 28652 9181 28698
rect 9077 28595 9181 28652
rect 9077 28549 9106 28595
rect 9152 28549 9181 28595
rect 9077 28492 9181 28549
rect 9077 28446 9106 28492
rect 9152 28446 9181 28492
rect 9077 28389 9181 28446
rect 9077 28343 9106 28389
rect 9152 28343 9181 28389
rect 9077 28286 9181 28343
rect 9077 28240 9106 28286
rect 9152 28240 9181 28286
rect 9077 28183 9181 28240
rect 9077 28137 9106 28183
rect 9152 28137 9181 28183
rect 9077 28080 9181 28137
rect 9077 28034 9106 28080
rect 9152 28034 9181 28080
rect 9077 27976 9181 28034
rect 9077 27930 9106 27976
rect 9152 27930 9181 27976
rect 9077 27917 9181 27930
rect 9321 28904 9425 28917
rect 9321 28858 9350 28904
rect 9396 28858 9425 28904
rect 9321 28801 9425 28858
rect 9321 28755 9350 28801
rect 9396 28755 9425 28801
rect 9321 28698 9425 28755
rect 9321 28652 9350 28698
rect 9396 28652 9425 28698
rect 9321 28595 9425 28652
rect 9321 28549 9350 28595
rect 9396 28549 9425 28595
rect 9321 28492 9425 28549
rect 9321 28446 9350 28492
rect 9396 28446 9425 28492
rect 9321 28389 9425 28446
rect 9321 28343 9350 28389
rect 9396 28343 9425 28389
rect 9321 28286 9425 28343
rect 9321 28240 9350 28286
rect 9396 28240 9425 28286
rect 9321 28183 9425 28240
rect 9321 28137 9350 28183
rect 9396 28137 9425 28183
rect 9321 28080 9425 28137
rect 9321 28034 9350 28080
rect 9396 28034 9425 28080
rect 9321 27976 9425 28034
rect 9321 27930 9350 27976
rect 9396 27930 9425 27976
rect 9321 27917 9425 27930
rect 9565 28904 9669 28917
rect 9565 28858 9594 28904
rect 9640 28858 9669 28904
rect 9565 28801 9669 28858
rect 9565 28755 9594 28801
rect 9640 28755 9669 28801
rect 9565 28698 9669 28755
rect 9565 28652 9594 28698
rect 9640 28652 9669 28698
rect 9565 28595 9669 28652
rect 9565 28549 9594 28595
rect 9640 28549 9669 28595
rect 9565 28492 9669 28549
rect 9565 28446 9594 28492
rect 9640 28446 9669 28492
rect 9565 28389 9669 28446
rect 9565 28343 9594 28389
rect 9640 28343 9669 28389
rect 9565 28286 9669 28343
rect 9565 28240 9594 28286
rect 9640 28240 9669 28286
rect 9565 28183 9669 28240
rect 9565 28137 9594 28183
rect 9640 28137 9669 28183
rect 9565 28080 9669 28137
rect 9565 28034 9594 28080
rect 9640 28034 9669 28080
rect 9565 27976 9669 28034
rect 9565 27930 9594 27976
rect 9640 27930 9669 27976
rect 9565 27917 9669 27930
rect 9809 28904 9913 28917
rect 9809 28858 9838 28904
rect 9884 28858 9913 28904
rect 9809 28801 9913 28858
rect 9809 28755 9838 28801
rect 9884 28755 9913 28801
rect 9809 28698 9913 28755
rect 9809 28652 9838 28698
rect 9884 28652 9913 28698
rect 9809 28595 9913 28652
rect 9809 28549 9838 28595
rect 9884 28549 9913 28595
rect 9809 28492 9913 28549
rect 9809 28446 9838 28492
rect 9884 28446 9913 28492
rect 9809 28389 9913 28446
rect 9809 28343 9838 28389
rect 9884 28343 9913 28389
rect 9809 28286 9913 28343
rect 9809 28240 9838 28286
rect 9884 28240 9913 28286
rect 9809 28183 9913 28240
rect 9809 28137 9838 28183
rect 9884 28137 9913 28183
rect 9809 28080 9913 28137
rect 9809 28034 9838 28080
rect 9884 28034 9913 28080
rect 9809 27976 9913 28034
rect 9809 27930 9838 27976
rect 9884 27930 9913 27976
rect 9809 27917 9913 27930
rect 10053 28904 10157 28917
rect 10053 28858 10082 28904
rect 10128 28858 10157 28904
rect 10053 28801 10157 28858
rect 10053 28755 10082 28801
rect 10128 28755 10157 28801
rect 10053 28698 10157 28755
rect 10053 28652 10082 28698
rect 10128 28652 10157 28698
rect 10053 28595 10157 28652
rect 10053 28549 10082 28595
rect 10128 28549 10157 28595
rect 10053 28492 10157 28549
rect 10053 28446 10082 28492
rect 10128 28446 10157 28492
rect 10053 28389 10157 28446
rect 10053 28343 10082 28389
rect 10128 28343 10157 28389
rect 10053 28286 10157 28343
rect 10053 28240 10082 28286
rect 10128 28240 10157 28286
rect 10053 28183 10157 28240
rect 10053 28137 10082 28183
rect 10128 28137 10157 28183
rect 10053 28080 10157 28137
rect 10053 28034 10082 28080
rect 10128 28034 10157 28080
rect 10053 27976 10157 28034
rect 10053 27930 10082 27976
rect 10128 27930 10157 27976
rect 10053 27917 10157 27930
rect 10297 28904 10385 28917
rect 10297 28858 10326 28904
rect 10372 28858 10385 28904
rect 10297 28801 10385 28858
rect 10297 28755 10326 28801
rect 10372 28755 10385 28801
rect 10297 28698 10385 28755
rect 10297 28652 10326 28698
rect 10372 28652 10385 28698
rect 10297 28595 10385 28652
rect 10297 28549 10326 28595
rect 10372 28549 10385 28595
rect 10297 28492 10385 28549
rect 10297 28446 10326 28492
rect 10372 28446 10385 28492
rect 10297 28389 10385 28446
rect 10297 28343 10326 28389
rect 10372 28343 10385 28389
rect 10297 28286 10385 28343
rect 10297 28240 10326 28286
rect 10372 28240 10385 28286
rect 10297 28183 10385 28240
rect 10297 28137 10326 28183
rect 10372 28137 10385 28183
rect 10297 28080 10385 28137
rect 10297 28034 10326 28080
rect 10372 28034 10385 28080
rect 10297 27976 10385 28034
rect 10297 27930 10326 27976
rect 10372 27930 10385 27976
rect 10297 27917 10385 27930
<< mvndiffc >>
rect 4054 26947 4100 26993
rect 4054 26844 4100 26890
rect 4054 26741 4100 26787
rect 4054 26638 4100 26684
rect 4054 26535 4100 26581
rect 4054 26432 4100 26478
rect 4054 26329 4100 26375
rect 4054 26226 4100 26272
rect 4054 26123 4100 26169
rect 4054 26019 4100 26065
rect 4298 26947 4344 26993
rect 4298 26844 4344 26890
rect 4298 26741 4344 26787
rect 4298 26638 4344 26684
rect 4298 26535 4344 26581
rect 4298 26432 4344 26478
rect 4298 26329 4344 26375
rect 4298 26226 4344 26272
rect 4298 26123 4344 26169
rect 4298 26019 4344 26065
rect 5116 26947 5162 26993
rect 5116 26844 5162 26890
rect 5116 26741 5162 26787
rect 5116 26638 5162 26684
rect 5116 26535 5162 26581
rect 5116 26432 5162 26478
rect 5116 26329 5162 26375
rect 5116 26226 5162 26272
rect 5116 26123 5162 26169
rect 5116 26019 5162 26065
rect 5360 26947 5406 26993
rect 5360 26844 5406 26890
rect 5360 26741 5406 26787
rect 5360 26638 5406 26684
rect 5360 26535 5406 26581
rect 5360 26432 5406 26478
rect 5360 26329 5406 26375
rect 5360 26226 5406 26272
rect 5360 26123 5406 26169
rect 5360 26019 5406 26065
rect 5604 26947 5650 26993
rect 5604 26844 5650 26890
rect 5604 26741 5650 26787
rect 5604 26638 5650 26684
rect 5604 26535 5650 26581
rect 5604 26432 5650 26478
rect 5604 26329 5650 26375
rect 5604 26226 5650 26272
rect 5604 26123 5650 26169
rect 5604 26019 5650 26065
rect 5848 26947 5894 26993
rect 5848 26844 5894 26890
rect 5848 26741 5894 26787
rect 5848 26638 5894 26684
rect 5848 26535 5894 26581
rect 5848 26432 5894 26478
rect 5848 26329 5894 26375
rect 5848 26226 5894 26272
rect 5848 26123 5894 26169
rect 5848 26019 5894 26065
rect 6092 26947 6138 26993
rect 6092 26844 6138 26890
rect 6092 26741 6138 26787
rect 6092 26638 6138 26684
rect 6092 26535 6138 26581
rect 6092 26432 6138 26478
rect 6092 26329 6138 26375
rect 6092 26226 6138 26272
rect 6092 26123 6138 26169
rect 6092 26019 6138 26065
rect 6336 26947 6382 26993
rect 6336 26844 6382 26890
rect 6336 26741 6382 26787
rect 6336 26638 6382 26684
rect 6336 26535 6382 26581
rect 6336 26432 6382 26478
rect 6336 26329 6382 26375
rect 6336 26226 6382 26272
rect 6336 26123 6382 26169
rect 6336 26019 6382 26065
rect 6580 26947 6626 26993
rect 6580 26844 6626 26890
rect 6580 26741 6626 26787
rect 6580 26638 6626 26684
rect 6580 26535 6626 26581
rect 6580 26432 6626 26478
rect 6580 26329 6626 26375
rect 6580 26226 6626 26272
rect 6580 26123 6626 26169
rect 6580 26019 6626 26065
rect 6824 26947 6870 26993
rect 6824 26844 6870 26890
rect 6824 26741 6870 26787
rect 6824 26638 6870 26684
rect 6824 26535 6870 26581
rect 6824 26432 6870 26478
rect 6824 26329 6870 26375
rect 6824 26226 6870 26272
rect 6824 26123 6870 26169
rect 6824 26019 6870 26065
rect 7068 26947 7114 26993
rect 7068 26844 7114 26890
rect 7068 26741 7114 26787
rect 7068 26638 7114 26684
rect 7068 26535 7114 26581
rect 7068 26432 7114 26478
rect 7068 26329 7114 26375
rect 7068 26226 7114 26272
rect 7068 26123 7114 26169
rect 7068 26019 7114 26065
rect 7312 26947 7358 26993
rect 7312 26844 7358 26890
rect 7312 26741 7358 26787
rect 7312 26638 7358 26684
rect 7312 26535 7358 26581
rect 7312 26432 7358 26478
rect 7312 26329 7358 26375
rect 7312 26226 7358 26272
rect 7312 26123 7358 26169
rect 7312 26019 7358 26065
rect 7556 26947 7602 26993
rect 7556 26844 7602 26890
rect 7556 26741 7602 26787
rect 7556 26638 7602 26684
rect 7556 26535 7602 26581
rect 7556 26432 7602 26478
rect 7556 26329 7602 26375
rect 7556 26226 7602 26272
rect 7556 26123 7602 26169
rect 7556 26019 7602 26065
rect 7800 26947 7846 26993
rect 7800 26844 7846 26890
rect 7800 26741 7846 26787
rect 7800 26638 7846 26684
rect 7800 26535 7846 26581
rect 7800 26432 7846 26478
rect 7800 26329 7846 26375
rect 7800 26226 7846 26272
rect 7800 26123 7846 26169
rect 7800 26019 7846 26065
rect 8044 26947 8090 26993
rect 8044 26844 8090 26890
rect 8044 26741 8090 26787
rect 8044 26638 8090 26684
rect 8044 26535 8090 26581
rect 8044 26432 8090 26478
rect 8044 26329 8090 26375
rect 8044 26226 8090 26272
rect 8044 26123 8090 26169
rect 8044 26019 8090 26065
<< mvpdiffc >>
rect 2590 28858 2636 28904
rect 2590 28755 2636 28801
rect 2590 28652 2636 28698
rect 2590 28549 2636 28595
rect 2590 28446 2636 28492
rect 2590 28343 2636 28389
rect 2590 28240 2636 28286
rect 2590 28137 2636 28183
rect 2590 28034 2636 28080
rect 2590 27930 2636 27976
rect 2834 28858 2880 28904
rect 2834 28755 2880 28801
rect 2834 28652 2880 28698
rect 2834 28549 2880 28595
rect 2834 28446 2880 28492
rect 2834 28343 2880 28389
rect 2834 28240 2880 28286
rect 2834 28137 2880 28183
rect 2834 28034 2880 28080
rect 2834 27930 2880 27976
rect 3078 28858 3124 28904
rect 3078 28755 3124 28801
rect 3078 28652 3124 28698
rect 3078 28549 3124 28595
rect 3078 28446 3124 28492
rect 3078 28343 3124 28389
rect 3078 28240 3124 28286
rect 3078 28137 3124 28183
rect 3078 28034 3124 28080
rect 3078 27930 3124 27976
rect 3322 28858 3368 28904
rect 3322 28755 3368 28801
rect 3322 28652 3368 28698
rect 3322 28549 3368 28595
rect 3322 28446 3368 28492
rect 3322 28343 3368 28389
rect 3322 28240 3368 28286
rect 3322 28137 3368 28183
rect 3322 28034 3368 28080
rect 3322 27930 3368 27976
rect 3566 28858 3612 28904
rect 3566 28755 3612 28801
rect 3566 28652 3612 28698
rect 3566 28549 3612 28595
rect 3566 28446 3612 28492
rect 3566 28343 3612 28389
rect 3566 28240 3612 28286
rect 3566 28137 3612 28183
rect 3566 28034 3612 28080
rect 3566 27930 3612 27976
rect 3810 28858 3856 28904
rect 3810 28755 3856 28801
rect 3810 28652 3856 28698
rect 3810 28549 3856 28595
rect 3810 28446 3856 28492
rect 3810 28343 3856 28389
rect 3810 28240 3856 28286
rect 3810 28137 3856 28183
rect 3810 28034 3856 28080
rect 3810 27930 3856 27976
rect 4054 28858 4100 28904
rect 4054 28755 4100 28801
rect 4054 28652 4100 28698
rect 4054 28549 4100 28595
rect 4054 28446 4100 28492
rect 4054 28343 4100 28389
rect 4054 28240 4100 28286
rect 4054 28137 4100 28183
rect 4054 28034 4100 28080
rect 4054 27930 4100 27976
rect 4298 28858 4344 28904
rect 4298 28755 4344 28801
rect 4298 28652 4344 28698
rect 4298 28549 4344 28595
rect 4298 28446 4344 28492
rect 4298 28343 4344 28389
rect 4298 28240 4344 28286
rect 4298 28137 4344 28183
rect 4298 28034 4344 28080
rect 4298 27930 4344 27976
rect 4470 28858 4516 28904
rect 4470 28755 4516 28801
rect 4470 28652 4516 28698
rect 4470 28549 4516 28595
rect 4470 28446 4516 28492
rect 4470 28343 4516 28389
rect 4470 28240 4516 28286
rect 4470 28137 4516 28183
rect 4470 28034 4516 28080
rect 4470 27930 4516 27976
rect 4714 28858 4760 28904
rect 4714 28755 4760 28801
rect 4714 28652 4760 28698
rect 4714 28549 4760 28595
rect 4714 28446 4760 28492
rect 4714 28343 4760 28389
rect 4714 28240 4760 28286
rect 4714 28137 4760 28183
rect 4714 28034 4760 28080
rect 4714 27930 4760 27976
rect 4958 28858 5004 28904
rect 4958 28755 5004 28801
rect 4958 28652 5004 28698
rect 4958 28549 5004 28595
rect 4958 28446 5004 28492
rect 4958 28343 5004 28389
rect 4958 28240 5004 28286
rect 4958 28137 5004 28183
rect 4958 28034 5004 28080
rect 4958 27930 5004 27976
rect 5202 28858 5248 28904
rect 5202 28755 5248 28801
rect 5202 28652 5248 28698
rect 5202 28549 5248 28595
rect 5202 28446 5248 28492
rect 5202 28343 5248 28389
rect 5202 28240 5248 28286
rect 5202 28137 5248 28183
rect 5202 28034 5248 28080
rect 5202 27930 5248 27976
rect 5446 28858 5492 28904
rect 5446 28755 5492 28801
rect 5446 28652 5492 28698
rect 5446 28549 5492 28595
rect 5446 28446 5492 28492
rect 5446 28343 5492 28389
rect 5446 28240 5492 28286
rect 5446 28137 5492 28183
rect 5446 28034 5492 28080
rect 5446 27930 5492 27976
rect 5690 28858 5736 28904
rect 5690 28755 5736 28801
rect 5690 28652 5736 28698
rect 5690 28549 5736 28595
rect 5690 28446 5736 28492
rect 5690 28343 5736 28389
rect 5690 28240 5736 28286
rect 5690 28137 5736 28183
rect 5690 28034 5736 28080
rect 5690 27930 5736 27976
rect 5934 28858 5980 28904
rect 5934 28755 5980 28801
rect 5934 28652 5980 28698
rect 5934 28549 5980 28595
rect 5934 28446 5980 28492
rect 5934 28343 5980 28389
rect 5934 28240 5980 28286
rect 5934 28137 5980 28183
rect 5934 28034 5980 28080
rect 5934 27930 5980 27976
rect 6178 28858 6224 28904
rect 6178 28755 6224 28801
rect 6178 28652 6224 28698
rect 6178 28549 6224 28595
rect 6178 28446 6224 28492
rect 6178 28343 6224 28389
rect 6178 28240 6224 28286
rect 6178 28137 6224 28183
rect 6178 28034 6224 28080
rect 6178 27930 6224 27976
rect 6422 28858 6468 28904
rect 6422 28755 6468 28801
rect 6422 28652 6468 28698
rect 6422 28549 6468 28595
rect 6422 28446 6468 28492
rect 6422 28343 6468 28389
rect 6422 28240 6468 28286
rect 6422 28137 6468 28183
rect 6422 28034 6468 28080
rect 6422 27930 6468 27976
rect 6666 28858 6712 28904
rect 6666 28755 6712 28801
rect 6666 28652 6712 28698
rect 6666 28549 6712 28595
rect 6666 28446 6712 28492
rect 6666 28343 6712 28389
rect 6666 28240 6712 28286
rect 6666 28137 6712 28183
rect 6666 28034 6712 28080
rect 6666 27930 6712 27976
rect 6910 28858 6956 28904
rect 6910 28755 6956 28801
rect 6910 28652 6956 28698
rect 6910 28549 6956 28595
rect 6910 28446 6956 28492
rect 6910 28343 6956 28389
rect 6910 28240 6956 28286
rect 6910 28137 6956 28183
rect 6910 28034 6956 28080
rect 6910 27930 6956 27976
rect 7154 28858 7200 28904
rect 7154 28755 7200 28801
rect 7154 28652 7200 28698
rect 7154 28549 7200 28595
rect 7154 28446 7200 28492
rect 7154 28343 7200 28389
rect 7154 28240 7200 28286
rect 7154 28137 7200 28183
rect 7154 28034 7200 28080
rect 7154 27930 7200 27976
rect 7398 28858 7444 28904
rect 7398 28755 7444 28801
rect 7398 28652 7444 28698
rect 7398 28549 7444 28595
rect 7398 28446 7444 28492
rect 7398 28343 7444 28389
rect 7398 28240 7444 28286
rect 7398 28137 7444 28183
rect 7398 28034 7444 28080
rect 7398 27930 7444 27976
rect 7642 28858 7688 28904
rect 7642 28755 7688 28801
rect 7642 28652 7688 28698
rect 7642 28549 7688 28595
rect 7642 28446 7688 28492
rect 7642 28343 7688 28389
rect 7642 28240 7688 28286
rect 7642 28137 7688 28183
rect 7642 28034 7688 28080
rect 7642 27930 7688 27976
rect 7886 28858 7932 28904
rect 7886 28755 7932 28801
rect 7886 28652 7932 28698
rect 7886 28549 7932 28595
rect 7886 28446 7932 28492
rect 7886 28343 7932 28389
rect 7886 28240 7932 28286
rect 7886 28137 7932 28183
rect 7886 28034 7932 28080
rect 7886 27930 7932 27976
rect 8130 28858 8176 28904
rect 8130 28755 8176 28801
rect 8130 28652 8176 28698
rect 8130 28549 8176 28595
rect 8130 28446 8176 28492
rect 8130 28343 8176 28389
rect 8130 28240 8176 28286
rect 8130 28137 8176 28183
rect 8130 28034 8176 28080
rect 8130 27930 8176 27976
rect 8374 28858 8420 28904
rect 8374 28755 8420 28801
rect 8374 28652 8420 28698
rect 8374 28549 8420 28595
rect 8374 28446 8420 28492
rect 8374 28343 8420 28389
rect 8374 28240 8420 28286
rect 8374 28137 8420 28183
rect 8374 28034 8420 28080
rect 8374 27930 8420 27976
rect 8618 28858 8664 28904
rect 8618 28755 8664 28801
rect 8618 28652 8664 28698
rect 8618 28549 8664 28595
rect 8618 28446 8664 28492
rect 8618 28343 8664 28389
rect 8618 28240 8664 28286
rect 8618 28137 8664 28183
rect 8618 28034 8664 28080
rect 8618 27930 8664 27976
rect 8862 28858 8908 28904
rect 8862 28755 8908 28801
rect 8862 28652 8908 28698
rect 8862 28549 8908 28595
rect 8862 28446 8908 28492
rect 8862 28343 8908 28389
rect 8862 28240 8908 28286
rect 8862 28137 8908 28183
rect 8862 28034 8908 28080
rect 8862 27930 8908 27976
rect 9106 28858 9152 28904
rect 9106 28755 9152 28801
rect 9106 28652 9152 28698
rect 9106 28549 9152 28595
rect 9106 28446 9152 28492
rect 9106 28343 9152 28389
rect 9106 28240 9152 28286
rect 9106 28137 9152 28183
rect 9106 28034 9152 28080
rect 9106 27930 9152 27976
rect 9350 28858 9396 28904
rect 9350 28755 9396 28801
rect 9350 28652 9396 28698
rect 9350 28549 9396 28595
rect 9350 28446 9396 28492
rect 9350 28343 9396 28389
rect 9350 28240 9396 28286
rect 9350 28137 9396 28183
rect 9350 28034 9396 28080
rect 9350 27930 9396 27976
rect 9594 28858 9640 28904
rect 9594 28755 9640 28801
rect 9594 28652 9640 28698
rect 9594 28549 9640 28595
rect 9594 28446 9640 28492
rect 9594 28343 9640 28389
rect 9594 28240 9640 28286
rect 9594 28137 9640 28183
rect 9594 28034 9640 28080
rect 9594 27930 9640 27976
rect 9838 28858 9884 28904
rect 9838 28755 9884 28801
rect 9838 28652 9884 28698
rect 9838 28549 9884 28595
rect 9838 28446 9884 28492
rect 9838 28343 9884 28389
rect 9838 28240 9884 28286
rect 9838 28137 9884 28183
rect 9838 28034 9884 28080
rect 9838 27930 9884 27976
rect 10082 28858 10128 28904
rect 10082 28755 10128 28801
rect 10082 28652 10128 28698
rect 10082 28549 10128 28595
rect 10082 28446 10128 28492
rect 10082 28343 10128 28389
rect 10082 28240 10128 28286
rect 10082 28137 10128 28183
rect 10082 28034 10128 28080
rect 10082 27930 10128 27976
rect 10326 28858 10372 28904
rect 10326 28755 10372 28801
rect 10326 28652 10372 28698
rect 10326 28549 10372 28595
rect 10326 28446 10372 28492
rect 10326 28343 10372 28389
rect 10326 28240 10372 28286
rect 10326 28137 10372 28183
rect 10326 28034 10372 28080
rect 10326 27930 10372 27976
<< psubdiff >>
rect 2253 27485 10709 27507
rect 2253 27439 3748 27485
rect 6520 27439 6889 27485
rect 10225 27439 10709 27485
rect 2253 27417 10709 27439
rect 2253 27156 2343 27417
rect 2253 25888 2275 27156
rect 2321 25888 2343 27156
rect 10619 27156 10709 27417
rect 2253 25802 2343 25888
rect 10619 25888 10641 27156
rect 10687 25888 10709 27156
rect 10619 25802 10709 25888
rect 2253 25780 10709 25802
rect 2253 25734 2275 25780
rect 6739 25734 6975 25780
rect 7209 25734 7445 25780
rect 7679 25734 8009 25780
rect 10687 25734 10709 25780
rect 2253 25712 10709 25734
<< nsubdiff >>
rect 2253 29188 10709 29210
rect 2253 29142 2275 29188
rect 10687 29142 10709 29188
rect 2253 29120 10709 29142
rect 2253 29034 2343 29120
rect 2253 27860 2275 29034
rect 2321 27860 2343 29034
rect 10619 29034 10709 29120
rect 2253 27838 2343 27860
rect 10619 27860 10641 29034
rect 10687 27860 10709 29034
rect 10619 27838 10709 27860
<< psubdiffcont >>
rect 3748 27439 6520 27485
rect 6889 27439 10225 27485
rect 2275 25888 2321 27156
rect 10641 25888 10687 27156
rect 2275 25734 6739 25780
rect 6975 25734 7209 25780
rect 7445 25734 7679 25780
rect 8009 25734 10687 25780
<< nsubdiffcont >>
rect 2275 29142 10687 29188
rect 2275 27860 2321 29034
rect 10641 27860 10687 29034
<< polysilicon >>
rect 2665 28917 2805 28961
rect 2909 28917 3049 28961
rect 3153 28917 3293 28961
rect 3397 28917 3537 28961
rect 3641 28917 3781 28961
rect 3885 28917 4025 28961
rect 4129 28917 4269 28961
rect 4545 28917 4685 28961
rect 4789 28917 4929 28961
rect 5033 28917 5173 28961
rect 5277 28917 5417 28961
rect 5521 28917 5661 28961
rect 5765 28917 5905 28961
rect 6009 28917 6149 28961
rect 6253 28917 6393 28961
rect 6497 28917 6637 28961
rect 6741 28917 6881 28961
rect 6985 28917 7125 28961
rect 7229 28917 7369 28961
rect 7473 28917 7613 28961
rect 7717 28917 7857 28961
rect 7961 28917 8101 28961
rect 8205 28917 8345 28961
rect 8449 28917 8589 28961
rect 8693 28917 8833 28961
rect 8937 28917 9077 28961
rect 9181 28917 9321 28961
rect 9425 28917 9565 28961
rect 9669 28917 9809 28961
rect 9913 28917 10053 28961
rect 10157 28917 10297 28961
rect 2665 27729 2805 27917
rect 2909 27729 3049 27917
rect 3153 27729 3293 27917
rect 3397 27729 3537 27917
rect 2665 27710 3537 27729
rect 2665 27664 2749 27710
rect 3453 27664 3537 27710
rect 2665 27645 3537 27664
rect 3641 27729 3781 27917
rect 3885 27729 4025 27917
rect 4129 27729 4269 27917
rect 3641 27710 4269 27729
rect 3641 27664 3697 27710
rect 4213 27664 4269 27710
rect 3641 27645 4269 27664
rect 4545 27729 4685 27917
rect 4789 27729 4929 27917
rect 5033 27729 5173 27917
rect 5277 27729 5417 27917
rect 5521 27729 5661 27917
rect 5765 27729 5905 27917
rect 6009 27729 6149 27917
rect 6253 27729 6393 27917
rect 6497 27729 6637 27917
rect 6741 27729 6881 27917
rect 6985 27729 7125 27917
rect 7229 27729 7369 27917
rect 7473 27729 7613 27917
rect 7717 27729 7857 27917
rect 7961 27729 8101 27917
rect 8205 27729 8345 27917
rect 8449 27729 8589 27917
rect 8693 27729 8833 27917
rect 8937 27729 9077 27917
rect 9181 27729 9321 27917
rect 9425 27729 9565 27917
rect 9669 27729 9809 27917
rect 9913 27729 10053 27917
rect 10157 27729 10297 27917
rect 4545 27710 10297 27729
rect 4545 27664 4578 27710
rect 10264 27664 10297 27710
rect 4545 27645 10297 27664
rect 5191 27259 6551 27278
rect 5191 27213 5237 27259
rect 6505 27213 6551 27259
rect 5191 27194 6551 27213
rect 4053 27131 4269 27150
rect 4053 27085 4072 27131
rect 4212 27085 4269 27131
rect 4053 27066 4269 27085
rect 4129 27006 4269 27066
rect 5191 27006 5331 27194
rect 5435 27006 5575 27194
rect 5679 27006 5819 27194
rect 5923 27006 6063 27194
rect 6167 27006 6307 27194
rect 6411 27006 6551 27194
rect 6655 27259 8015 27278
rect 6655 27213 6701 27259
rect 7969 27213 8015 27259
rect 6655 27194 8015 27213
rect 6655 27006 6795 27194
rect 6899 27006 7039 27194
rect 7143 27006 7283 27194
rect 7387 27006 7527 27194
rect 7631 27006 7771 27194
rect 7875 27006 8015 27194
rect 4129 25962 4269 26006
rect 5191 25962 5331 26006
rect 5435 25962 5575 26006
rect 5679 25962 5819 26006
rect 5923 25962 6063 26006
rect 6167 25962 6307 26006
rect 6411 25962 6551 26006
rect 6655 25962 6795 26006
rect 6899 25962 7039 26006
rect 7143 25962 7283 26006
rect 7387 25962 7527 26006
rect 7631 25962 7771 26006
rect 7875 25962 8015 26006
<< polycontact >>
rect 2749 27664 3453 27710
rect 3697 27664 4213 27710
rect 4578 27664 10264 27710
rect 5237 27213 6505 27259
rect 4072 27085 4212 27131
rect 6701 27213 7969 27259
<< metal1 >>
rect 1481 45914 1665 45926
rect 1481 45862 1493 45914
rect 1545 45862 1601 45914
rect 1653 45862 1665 45914
rect 1481 45850 1665 45862
rect 3851 45914 4035 45926
rect 3851 45862 3863 45914
rect 3915 45862 3971 45914
rect 4023 45862 4035 45914
rect 3851 45850 4035 45862
rect 6227 45914 6735 45926
rect 6227 45862 6239 45914
rect 6291 45862 6347 45914
rect 6399 45862 6455 45914
rect 6507 45862 6563 45914
rect 6615 45862 6671 45914
rect 6723 45862 6735 45914
rect 6227 45850 6735 45862
rect 8927 45914 9111 45926
rect 8927 45862 8939 45914
rect 8991 45862 9047 45914
rect 9099 45862 9111 45914
rect 8927 45850 9111 45862
rect 11297 45914 11481 45926
rect 11297 45862 11309 45914
rect 11361 45862 11417 45914
rect 11469 45862 11481 45914
rect 11297 45850 11481 45862
rect 1481 42174 1665 42186
rect 1481 42122 1493 42174
rect 1545 42122 1601 42174
rect 1653 42122 1665 42174
rect 1481 42110 1665 42122
rect 3851 42174 4035 42186
rect 3851 42122 3863 42174
rect 3915 42122 3971 42174
rect 4023 42122 4035 42174
rect 3851 42110 4035 42122
rect 6227 42174 6735 42186
rect 6227 42122 6239 42174
rect 6291 42122 6347 42174
rect 6399 42122 6455 42174
rect 6507 42122 6563 42174
rect 6615 42122 6671 42174
rect 6723 42122 6735 42174
rect 6227 42110 6735 42122
rect 8927 42174 9111 42186
rect 8927 42122 8939 42174
rect 8991 42122 9047 42174
rect 9099 42122 9111 42174
rect 8927 42110 9111 42122
rect 11297 42174 11481 42186
rect 11297 42122 11309 42174
rect 11361 42122 11417 42174
rect 11469 42122 11481 42174
rect 11297 42110 11481 42122
rect 1748 41735 3768 41747
rect 1748 41683 1760 41735
rect 1812 41683 1868 41735
rect 1920 41683 1976 41735
rect 2028 41683 2084 41735
rect 2136 41683 2192 41735
rect 2244 41683 2300 41735
rect 2352 41683 2408 41735
rect 2460 41683 2516 41735
rect 2568 41683 2624 41735
rect 2676 41683 2732 41735
rect 2784 41683 2840 41735
rect 2892 41683 2948 41735
rect 3000 41683 3056 41735
rect 3108 41683 3164 41735
rect 3216 41683 3272 41735
rect 3324 41683 3380 41735
rect 3432 41683 3488 41735
rect 3540 41683 3596 41735
rect 3648 41683 3704 41735
rect 3756 41683 3768 41735
rect 1748 41627 3768 41683
rect 1748 41575 1760 41627
rect 1812 41575 1868 41627
rect 1920 41575 1976 41627
rect 2028 41575 2084 41627
rect 2136 41575 2192 41627
rect 2244 41575 2300 41627
rect 2352 41575 2408 41627
rect 2460 41575 2516 41627
rect 2568 41575 2624 41627
rect 2676 41575 2732 41627
rect 2784 41575 2840 41627
rect 2892 41575 2948 41627
rect 3000 41575 3056 41627
rect 3108 41575 3164 41627
rect 3216 41575 3272 41627
rect 3324 41575 3380 41627
rect 3432 41575 3488 41627
rect 3540 41575 3596 41627
rect 3648 41575 3704 41627
rect 3756 41575 3768 41627
rect 1748 41563 3768 41575
rect 4118 41735 6138 41747
rect 4118 41683 4130 41735
rect 4182 41683 4238 41735
rect 4290 41683 4346 41735
rect 4398 41683 4454 41735
rect 4506 41683 4562 41735
rect 4614 41683 4670 41735
rect 4722 41683 4778 41735
rect 4830 41683 4886 41735
rect 4938 41683 4994 41735
rect 5046 41683 5102 41735
rect 5154 41683 5210 41735
rect 5262 41683 5318 41735
rect 5370 41683 5426 41735
rect 5478 41683 5534 41735
rect 5586 41683 5642 41735
rect 5694 41683 5750 41735
rect 5802 41683 5858 41735
rect 5910 41683 5966 41735
rect 6018 41683 6074 41735
rect 6126 41683 6138 41735
rect 4118 41627 6138 41683
rect 4118 41575 4130 41627
rect 4182 41575 4238 41627
rect 4290 41575 4346 41627
rect 4398 41575 4454 41627
rect 4506 41575 4562 41627
rect 4614 41575 4670 41627
rect 4722 41575 4778 41627
rect 4830 41575 4886 41627
rect 4938 41575 4994 41627
rect 5046 41575 5102 41627
rect 5154 41575 5210 41627
rect 5262 41575 5318 41627
rect 5370 41575 5426 41627
rect 5478 41575 5534 41627
rect 5586 41575 5642 41627
rect 5694 41575 5750 41627
rect 5802 41575 5858 41627
rect 5910 41575 5966 41627
rect 6018 41575 6074 41627
rect 6126 41575 6138 41627
rect 4118 41563 6138 41575
rect 6824 41735 8844 41747
rect 6824 41683 6836 41735
rect 6888 41683 6944 41735
rect 6996 41683 7052 41735
rect 7104 41683 7160 41735
rect 7212 41683 7268 41735
rect 7320 41683 7376 41735
rect 7428 41683 7484 41735
rect 7536 41683 7592 41735
rect 7644 41683 7700 41735
rect 7752 41683 7808 41735
rect 7860 41683 7916 41735
rect 7968 41683 8024 41735
rect 8076 41683 8132 41735
rect 8184 41683 8240 41735
rect 8292 41683 8348 41735
rect 8400 41683 8456 41735
rect 8508 41683 8564 41735
rect 8616 41683 8672 41735
rect 8724 41683 8780 41735
rect 8832 41683 8844 41735
rect 6824 41627 8844 41683
rect 6824 41575 6836 41627
rect 6888 41575 6944 41627
rect 6996 41575 7052 41627
rect 7104 41575 7160 41627
rect 7212 41575 7268 41627
rect 7320 41575 7376 41627
rect 7428 41575 7484 41627
rect 7536 41575 7592 41627
rect 7644 41575 7700 41627
rect 7752 41575 7808 41627
rect 7860 41575 7916 41627
rect 7968 41575 8024 41627
rect 8076 41575 8132 41627
rect 8184 41575 8240 41627
rect 8292 41575 8348 41627
rect 8400 41575 8456 41627
rect 8508 41575 8564 41627
rect 8616 41575 8672 41627
rect 8724 41575 8780 41627
rect 8832 41575 8844 41627
rect 6824 41563 8844 41575
rect 9194 41735 11214 41747
rect 9194 41683 9206 41735
rect 9258 41683 9314 41735
rect 9366 41683 9422 41735
rect 9474 41683 9530 41735
rect 9582 41683 9638 41735
rect 9690 41683 9746 41735
rect 9798 41683 9854 41735
rect 9906 41683 9962 41735
rect 10014 41683 10070 41735
rect 10122 41683 10178 41735
rect 10230 41683 10286 41735
rect 10338 41683 10394 41735
rect 10446 41683 10502 41735
rect 10554 41683 10610 41735
rect 10662 41683 10718 41735
rect 10770 41683 10826 41735
rect 10878 41683 10934 41735
rect 10986 41683 11042 41735
rect 11094 41683 11150 41735
rect 11202 41683 11214 41735
rect 9194 41627 11214 41683
rect 9194 41575 9206 41627
rect 9258 41575 9314 41627
rect 9366 41575 9422 41627
rect 9474 41575 9530 41627
rect 9582 41575 9638 41627
rect 9690 41575 9746 41627
rect 9798 41575 9854 41627
rect 9906 41575 9962 41627
rect 10014 41575 10070 41627
rect 10122 41575 10178 41627
rect 10230 41575 10286 41627
rect 10338 41575 10394 41627
rect 10446 41575 10502 41627
rect 10554 41575 10610 41627
rect 10662 41575 10718 41627
rect 10770 41575 10826 41627
rect 10878 41575 10934 41627
rect 10986 41575 11042 41627
rect 11094 41575 11150 41627
rect 11202 41575 11214 41627
rect 9194 41563 11214 41575
rect 1790 35998 3726 36010
rect 1790 35946 1802 35998
rect 1854 35946 1926 35998
rect 1978 35946 2050 35998
rect 2102 35946 2174 35998
rect 2226 35946 2298 35998
rect 2350 35946 2422 35998
rect 2474 35946 2546 35998
rect 2598 35946 2670 35998
rect 2722 35946 2794 35998
rect 2846 35946 2918 35998
rect 2970 35946 3042 35998
rect 3094 35946 3166 35998
rect 3218 35946 3290 35998
rect 3342 35946 3414 35998
rect 3466 35946 3538 35998
rect 3590 35946 3662 35998
rect 3714 35946 3726 35998
rect 1790 35874 3726 35946
rect 1790 35822 1802 35874
rect 1854 35822 1926 35874
rect 1978 35822 2050 35874
rect 2102 35822 2174 35874
rect 2226 35822 2298 35874
rect 2350 35822 2422 35874
rect 2474 35822 2546 35874
rect 2598 35822 2670 35874
rect 2722 35822 2794 35874
rect 2846 35822 2918 35874
rect 2970 35822 3042 35874
rect 3094 35822 3166 35874
rect 3218 35822 3290 35874
rect 3342 35822 3414 35874
rect 3466 35822 3538 35874
rect 3590 35822 3662 35874
rect 3714 35822 3726 35874
rect 1790 35750 3726 35822
rect 1790 35698 1802 35750
rect 1854 35698 1926 35750
rect 1978 35698 2050 35750
rect 2102 35698 2174 35750
rect 2226 35698 2298 35750
rect 2350 35698 2422 35750
rect 2474 35698 2546 35750
rect 2598 35698 2670 35750
rect 2722 35698 2794 35750
rect 2846 35698 2918 35750
rect 2970 35698 3042 35750
rect 3094 35698 3166 35750
rect 3218 35698 3290 35750
rect 3342 35698 3414 35750
rect 3466 35698 3538 35750
rect 3590 35698 3662 35750
rect 3714 35698 3726 35750
rect 1790 35626 3726 35698
rect 1790 35574 1802 35626
rect 1854 35574 1926 35626
rect 1978 35574 2050 35626
rect 2102 35574 2174 35626
rect 2226 35574 2298 35626
rect 2350 35574 2422 35626
rect 2474 35574 2546 35626
rect 2598 35574 2670 35626
rect 2722 35574 2794 35626
rect 2846 35574 2918 35626
rect 2970 35574 3042 35626
rect 3094 35574 3166 35626
rect 3218 35574 3290 35626
rect 3342 35574 3414 35626
rect 3466 35574 3538 35626
rect 3590 35574 3662 35626
rect 3714 35574 3726 35626
rect 1790 35502 3726 35574
rect 1790 35450 1802 35502
rect 1854 35450 1926 35502
rect 1978 35450 2050 35502
rect 2102 35450 2174 35502
rect 2226 35450 2298 35502
rect 2350 35450 2422 35502
rect 2474 35450 2546 35502
rect 2598 35450 2670 35502
rect 2722 35450 2794 35502
rect 2846 35450 2918 35502
rect 2970 35450 3042 35502
rect 3094 35450 3166 35502
rect 3218 35450 3290 35502
rect 3342 35450 3414 35502
rect 3466 35450 3538 35502
rect 3590 35450 3662 35502
rect 3714 35450 3726 35502
rect 1790 35378 3726 35450
rect 1790 35326 1802 35378
rect 1854 35326 1926 35378
rect 1978 35326 2050 35378
rect 2102 35326 2174 35378
rect 2226 35326 2298 35378
rect 2350 35326 2422 35378
rect 2474 35326 2546 35378
rect 2598 35326 2670 35378
rect 2722 35326 2794 35378
rect 2846 35326 2918 35378
rect 2970 35326 3042 35378
rect 3094 35326 3166 35378
rect 3218 35326 3290 35378
rect 3342 35326 3414 35378
rect 3466 35326 3538 35378
rect 3590 35326 3662 35378
rect 3714 35326 3726 35378
rect 1790 35314 3726 35326
rect 4160 35998 6096 36010
rect 4160 35946 4172 35998
rect 4224 35946 4296 35998
rect 4348 35946 4420 35998
rect 4472 35946 4544 35998
rect 4596 35946 4668 35998
rect 4720 35946 4792 35998
rect 4844 35946 4916 35998
rect 4968 35946 5040 35998
rect 5092 35946 5164 35998
rect 5216 35946 5288 35998
rect 5340 35946 5412 35998
rect 5464 35946 5536 35998
rect 5588 35946 5660 35998
rect 5712 35946 5784 35998
rect 5836 35946 5908 35998
rect 5960 35946 6032 35998
rect 6084 35946 6096 35998
rect 4160 35874 6096 35946
rect 4160 35822 4172 35874
rect 4224 35822 4296 35874
rect 4348 35822 4420 35874
rect 4472 35822 4544 35874
rect 4596 35822 4668 35874
rect 4720 35822 4792 35874
rect 4844 35822 4916 35874
rect 4968 35822 5040 35874
rect 5092 35822 5164 35874
rect 5216 35822 5288 35874
rect 5340 35822 5412 35874
rect 5464 35822 5536 35874
rect 5588 35822 5660 35874
rect 5712 35822 5784 35874
rect 5836 35822 5908 35874
rect 5960 35822 6032 35874
rect 6084 35822 6096 35874
rect 4160 35750 6096 35822
rect 4160 35698 4172 35750
rect 4224 35698 4296 35750
rect 4348 35698 4420 35750
rect 4472 35698 4544 35750
rect 4596 35698 4668 35750
rect 4720 35698 4792 35750
rect 4844 35698 4916 35750
rect 4968 35698 5040 35750
rect 5092 35698 5164 35750
rect 5216 35698 5288 35750
rect 5340 35698 5412 35750
rect 5464 35698 5536 35750
rect 5588 35698 5660 35750
rect 5712 35698 5784 35750
rect 5836 35698 5908 35750
rect 5960 35698 6032 35750
rect 6084 35698 6096 35750
rect 4160 35626 6096 35698
rect 4160 35574 4172 35626
rect 4224 35574 4296 35626
rect 4348 35574 4420 35626
rect 4472 35574 4544 35626
rect 4596 35574 4668 35626
rect 4720 35574 4792 35626
rect 4844 35574 4916 35626
rect 4968 35574 5040 35626
rect 5092 35574 5164 35626
rect 5216 35574 5288 35626
rect 5340 35574 5412 35626
rect 5464 35574 5536 35626
rect 5588 35574 5660 35626
rect 5712 35574 5784 35626
rect 5836 35574 5908 35626
rect 5960 35574 6032 35626
rect 6084 35574 6096 35626
rect 4160 35502 6096 35574
rect 4160 35450 4172 35502
rect 4224 35450 4296 35502
rect 4348 35450 4420 35502
rect 4472 35450 4544 35502
rect 4596 35450 4668 35502
rect 4720 35450 4792 35502
rect 4844 35450 4916 35502
rect 4968 35450 5040 35502
rect 5092 35450 5164 35502
rect 5216 35450 5288 35502
rect 5340 35450 5412 35502
rect 5464 35450 5536 35502
rect 5588 35450 5660 35502
rect 5712 35450 5784 35502
rect 5836 35450 5908 35502
rect 5960 35450 6032 35502
rect 6084 35450 6096 35502
rect 4160 35378 6096 35450
rect 4160 35326 4172 35378
rect 4224 35326 4296 35378
rect 4348 35326 4420 35378
rect 4472 35326 4544 35378
rect 4596 35326 4668 35378
rect 4720 35326 4792 35378
rect 4844 35326 4916 35378
rect 4968 35326 5040 35378
rect 5092 35326 5164 35378
rect 5216 35326 5288 35378
rect 5340 35326 5412 35378
rect 5464 35326 5536 35378
rect 5588 35326 5660 35378
rect 5712 35326 5784 35378
rect 5836 35326 5908 35378
rect 5960 35326 6032 35378
rect 6084 35326 6096 35378
rect 4160 35314 6096 35326
rect 6866 35998 8802 36010
rect 6866 35946 6878 35998
rect 6930 35946 7002 35998
rect 7054 35946 7126 35998
rect 7178 35946 7250 35998
rect 7302 35946 7374 35998
rect 7426 35946 7498 35998
rect 7550 35946 7622 35998
rect 7674 35946 7746 35998
rect 7798 35946 7870 35998
rect 7922 35946 7994 35998
rect 8046 35946 8118 35998
rect 8170 35946 8242 35998
rect 8294 35946 8366 35998
rect 8418 35946 8490 35998
rect 8542 35946 8614 35998
rect 8666 35946 8738 35998
rect 8790 35946 8802 35998
rect 6866 35874 8802 35946
rect 6866 35822 6878 35874
rect 6930 35822 7002 35874
rect 7054 35822 7126 35874
rect 7178 35822 7250 35874
rect 7302 35822 7374 35874
rect 7426 35822 7498 35874
rect 7550 35822 7622 35874
rect 7674 35822 7746 35874
rect 7798 35822 7870 35874
rect 7922 35822 7994 35874
rect 8046 35822 8118 35874
rect 8170 35822 8242 35874
rect 8294 35822 8366 35874
rect 8418 35822 8490 35874
rect 8542 35822 8614 35874
rect 8666 35822 8738 35874
rect 8790 35822 8802 35874
rect 6866 35750 8802 35822
rect 6866 35698 6878 35750
rect 6930 35698 7002 35750
rect 7054 35698 7126 35750
rect 7178 35698 7250 35750
rect 7302 35698 7374 35750
rect 7426 35698 7498 35750
rect 7550 35698 7622 35750
rect 7674 35698 7746 35750
rect 7798 35698 7870 35750
rect 7922 35698 7994 35750
rect 8046 35698 8118 35750
rect 8170 35698 8242 35750
rect 8294 35698 8366 35750
rect 8418 35698 8490 35750
rect 8542 35698 8614 35750
rect 8666 35698 8738 35750
rect 8790 35698 8802 35750
rect 6866 35626 8802 35698
rect 6866 35574 6878 35626
rect 6930 35574 7002 35626
rect 7054 35574 7126 35626
rect 7178 35574 7250 35626
rect 7302 35574 7374 35626
rect 7426 35574 7498 35626
rect 7550 35574 7622 35626
rect 7674 35574 7746 35626
rect 7798 35574 7870 35626
rect 7922 35574 7994 35626
rect 8046 35574 8118 35626
rect 8170 35574 8242 35626
rect 8294 35574 8366 35626
rect 8418 35574 8490 35626
rect 8542 35574 8614 35626
rect 8666 35574 8738 35626
rect 8790 35574 8802 35626
rect 6866 35502 8802 35574
rect 6866 35450 6878 35502
rect 6930 35450 7002 35502
rect 7054 35450 7126 35502
rect 7178 35450 7250 35502
rect 7302 35450 7374 35502
rect 7426 35450 7498 35502
rect 7550 35450 7622 35502
rect 7674 35450 7746 35502
rect 7798 35450 7870 35502
rect 7922 35450 7994 35502
rect 8046 35450 8118 35502
rect 8170 35450 8242 35502
rect 8294 35450 8366 35502
rect 8418 35450 8490 35502
rect 8542 35450 8614 35502
rect 8666 35450 8738 35502
rect 8790 35450 8802 35502
rect 6866 35378 8802 35450
rect 6866 35326 6878 35378
rect 6930 35326 7002 35378
rect 7054 35326 7126 35378
rect 7178 35326 7250 35378
rect 7302 35326 7374 35378
rect 7426 35326 7498 35378
rect 7550 35326 7622 35378
rect 7674 35326 7746 35378
rect 7798 35326 7870 35378
rect 7922 35326 7994 35378
rect 8046 35326 8118 35378
rect 8170 35326 8242 35378
rect 8294 35326 8366 35378
rect 8418 35326 8490 35378
rect 8542 35326 8614 35378
rect 8666 35326 8738 35378
rect 8790 35326 8802 35378
rect 6866 35314 8802 35326
rect 9236 35998 11172 36010
rect 9236 35946 9248 35998
rect 9300 35946 9372 35998
rect 9424 35946 9496 35998
rect 9548 35946 9620 35998
rect 9672 35946 9744 35998
rect 9796 35946 9868 35998
rect 9920 35946 9992 35998
rect 10044 35946 10116 35998
rect 10168 35946 10240 35998
rect 10292 35946 10364 35998
rect 10416 35946 10488 35998
rect 10540 35946 10612 35998
rect 10664 35946 10736 35998
rect 10788 35946 10860 35998
rect 10912 35946 10984 35998
rect 11036 35946 11108 35998
rect 11160 35946 11172 35998
rect 9236 35874 11172 35946
rect 9236 35822 9248 35874
rect 9300 35822 9372 35874
rect 9424 35822 9496 35874
rect 9548 35822 9620 35874
rect 9672 35822 9744 35874
rect 9796 35822 9868 35874
rect 9920 35822 9992 35874
rect 10044 35822 10116 35874
rect 10168 35822 10240 35874
rect 10292 35822 10364 35874
rect 10416 35822 10488 35874
rect 10540 35822 10612 35874
rect 10664 35822 10736 35874
rect 10788 35822 10860 35874
rect 10912 35822 10984 35874
rect 11036 35822 11108 35874
rect 11160 35822 11172 35874
rect 9236 35750 11172 35822
rect 9236 35698 9248 35750
rect 9300 35698 9372 35750
rect 9424 35698 9496 35750
rect 9548 35698 9620 35750
rect 9672 35698 9744 35750
rect 9796 35698 9868 35750
rect 9920 35698 9992 35750
rect 10044 35698 10116 35750
rect 10168 35698 10240 35750
rect 10292 35698 10364 35750
rect 10416 35698 10488 35750
rect 10540 35698 10612 35750
rect 10664 35698 10736 35750
rect 10788 35698 10860 35750
rect 10912 35698 10984 35750
rect 11036 35698 11108 35750
rect 11160 35698 11172 35750
rect 9236 35626 11172 35698
rect 9236 35574 9248 35626
rect 9300 35574 9372 35626
rect 9424 35574 9496 35626
rect 9548 35574 9620 35626
rect 9672 35574 9744 35626
rect 9796 35574 9868 35626
rect 9920 35574 9992 35626
rect 10044 35574 10116 35626
rect 10168 35574 10240 35626
rect 10292 35574 10364 35626
rect 10416 35574 10488 35626
rect 10540 35574 10612 35626
rect 10664 35574 10736 35626
rect 10788 35574 10860 35626
rect 10912 35574 10984 35626
rect 11036 35574 11108 35626
rect 11160 35574 11172 35626
rect 9236 35502 11172 35574
rect 9236 35450 9248 35502
rect 9300 35450 9372 35502
rect 9424 35450 9496 35502
rect 9548 35450 9620 35502
rect 9672 35450 9744 35502
rect 9796 35450 9868 35502
rect 9920 35450 9992 35502
rect 10044 35450 10116 35502
rect 10168 35450 10240 35502
rect 10292 35450 10364 35502
rect 10416 35450 10488 35502
rect 10540 35450 10612 35502
rect 10664 35450 10736 35502
rect 10788 35450 10860 35502
rect 10912 35450 10984 35502
rect 11036 35450 11108 35502
rect 11160 35450 11172 35502
rect 9236 35378 11172 35450
rect 9236 35326 9248 35378
rect 9300 35326 9372 35378
rect 9424 35326 9496 35378
rect 9548 35326 9620 35378
rect 9672 35326 9744 35378
rect 9796 35326 9868 35378
rect 9920 35326 9992 35378
rect 10044 35326 10116 35378
rect 10168 35326 10240 35378
rect 10292 35326 10364 35378
rect 10416 35326 10488 35378
rect 10540 35326 10612 35378
rect 10664 35326 10736 35378
rect 10788 35326 10860 35378
rect 10912 35326 10984 35378
rect 11036 35326 11108 35378
rect 11160 35326 11172 35378
rect 9236 35314 11172 35326
rect -50 27721 110 30038
rect 1748 29651 3768 29663
rect 1748 29599 1760 29651
rect 1812 29599 1868 29651
rect 1920 29599 1976 29651
rect 2028 29599 2084 29651
rect 2136 29599 2192 29651
rect 2244 29599 2300 29651
rect 2352 29599 2408 29651
rect 2460 29599 2516 29651
rect 2568 29599 2624 29651
rect 2676 29599 2732 29651
rect 2784 29599 2840 29651
rect 2892 29599 2948 29651
rect 3000 29599 3056 29651
rect 3108 29599 3164 29651
rect 3216 29599 3272 29651
rect 3324 29599 3380 29651
rect 3432 29599 3488 29651
rect 3540 29599 3596 29651
rect 3648 29599 3704 29651
rect 3756 29599 3768 29651
rect 1748 29543 3768 29599
rect 1748 29491 1760 29543
rect 1812 29491 1868 29543
rect 1920 29491 1976 29543
rect 2028 29491 2084 29543
rect 2136 29491 2192 29543
rect 2244 29491 2300 29543
rect 2352 29491 2408 29543
rect 2460 29491 2516 29543
rect 2568 29491 2624 29543
rect 2676 29491 2732 29543
rect 2784 29491 2840 29543
rect 2892 29491 2948 29543
rect 3000 29491 3056 29543
rect 3108 29491 3164 29543
rect 3216 29491 3272 29543
rect 3324 29491 3380 29543
rect 3432 29491 3488 29543
rect 3540 29491 3596 29543
rect 3648 29491 3704 29543
rect 3756 29491 3768 29543
rect 1748 29479 3768 29491
rect 4118 29651 6138 29663
rect 4118 29599 4130 29651
rect 4182 29599 4238 29651
rect 4290 29599 4346 29651
rect 4398 29599 4454 29651
rect 4506 29599 4562 29651
rect 4614 29599 4670 29651
rect 4722 29599 4778 29651
rect 4830 29599 4886 29651
rect 4938 29599 4994 29651
rect 5046 29599 5102 29651
rect 5154 29599 5210 29651
rect 5262 29599 5318 29651
rect 5370 29599 5426 29651
rect 5478 29599 5534 29651
rect 5586 29599 5642 29651
rect 5694 29599 5750 29651
rect 5802 29599 5858 29651
rect 5910 29599 5966 29651
rect 6018 29599 6074 29651
rect 6126 29599 6138 29651
rect 4118 29543 6138 29599
rect 4118 29491 4130 29543
rect 4182 29491 4238 29543
rect 4290 29491 4346 29543
rect 4398 29491 4454 29543
rect 4506 29491 4562 29543
rect 4614 29491 4670 29543
rect 4722 29491 4778 29543
rect 4830 29491 4886 29543
rect 4938 29491 4994 29543
rect 5046 29491 5102 29543
rect 5154 29491 5210 29543
rect 5262 29491 5318 29543
rect 5370 29491 5426 29543
rect 5478 29491 5534 29543
rect 5586 29491 5642 29543
rect 5694 29491 5750 29543
rect 5802 29491 5858 29543
rect 5910 29491 5966 29543
rect 6018 29491 6074 29543
rect 6126 29491 6138 29543
rect 4118 29479 6138 29491
rect 6824 29651 8844 29663
rect 6824 29599 6836 29651
rect 6888 29599 6944 29651
rect 6996 29599 7052 29651
rect 7104 29599 7160 29651
rect 7212 29599 7268 29651
rect 7320 29599 7376 29651
rect 7428 29599 7484 29651
rect 7536 29599 7592 29651
rect 7644 29599 7700 29651
rect 7752 29599 7808 29651
rect 7860 29599 7916 29651
rect 7968 29599 8024 29651
rect 8076 29599 8132 29651
rect 8184 29599 8240 29651
rect 8292 29599 8348 29651
rect 8400 29599 8456 29651
rect 8508 29599 8564 29651
rect 8616 29599 8672 29651
rect 8724 29599 8780 29651
rect 8832 29599 8844 29651
rect 6824 29543 8844 29599
rect 6824 29491 6836 29543
rect 6888 29491 6944 29543
rect 6996 29491 7052 29543
rect 7104 29491 7160 29543
rect 7212 29491 7268 29543
rect 7320 29491 7376 29543
rect 7428 29491 7484 29543
rect 7536 29491 7592 29543
rect 7644 29491 7700 29543
rect 7752 29491 7808 29543
rect 7860 29491 7916 29543
rect 7968 29491 8024 29543
rect 8076 29491 8132 29543
rect 8184 29491 8240 29543
rect 8292 29491 8348 29543
rect 8400 29491 8456 29543
rect 8508 29491 8564 29543
rect 8616 29491 8672 29543
rect 8724 29491 8780 29543
rect 8832 29491 8844 29543
rect 6824 29479 8844 29491
rect 9194 29651 11214 29663
rect 9194 29599 9206 29651
rect 9258 29599 9314 29651
rect 9366 29599 9422 29651
rect 9474 29599 9530 29651
rect 9582 29599 9638 29651
rect 9690 29599 9746 29651
rect 9798 29599 9854 29651
rect 9906 29599 9962 29651
rect 10014 29599 10070 29651
rect 10122 29599 10178 29651
rect 10230 29599 10286 29651
rect 10338 29599 10394 29651
rect 10446 29599 10502 29651
rect 10554 29599 10610 29651
rect 10662 29599 10718 29651
rect 10770 29599 10826 29651
rect 10878 29599 10934 29651
rect 10986 29599 11042 29651
rect 11094 29599 11150 29651
rect 11202 29599 11214 29651
rect 9194 29543 11214 29599
rect 9194 29491 9206 29543
rect 9258 29491 9314 29543
rect 9366 29491 9422 29543
rect 9474 29491 9530 29543
rect 9582 29491 9638 29543
rect 9690 29491 9746 29543
rect 9798 29491 9854 29543
rect 9906 29491 9962 29543
rect 10014 29491 10070 29543
rect 10122 29491 10178 29543
rect 10230 29491 10286 29543
rect 10338 29491 10394 29543
rect 10446 29491 10502 29543
rect 10554 29491 10610 29543
rect 10662 29491 10718 29543
rect 10770 29491 10826 29543
rect 10878 29491 10934 29543
rect 10986 29491 11042 29543
rect 11094 29491 11150 29543
rect 11202 29491 11214 29543
rect 9194 29479 11214 29491
rect 1473 29188 11489 29199
rect 1473 29187 2275 29188
rect 10687 29187 11489 29188
rect 1473 29135 1495 29187
rect 1651 29142 2275 29187
rect 10687 29142 11311 29187
rect 1651 29135 3865 29142
rect 4021 29135 6247 29142
rect 6715 29135 8941 29142
rect 9097 29135 11311 29142
rect 11467 29135 11489 29187
rect 1473 29131 11489 29135
rect 1473 29123 2332 29131
rect 2264 29034 2332 29123
rect 2264 27860 2275 29034
rect 2321 27860 2332 29034
rect 2575 28904 2651 29131
rect 2575 28858 2590 28904
rect 2636 28858 2651 28904
rect 2575 28801 2651 28858
rect 2575 28755 2590 28801
rect 2636 28755 2651 28801
rect 2575 28698 2651 28755
rect 2575 28652 2590 28698
rect 2636 28652 2651 28698
rect 2575 28595 2651 28652
rect 2575 28549 2590 28595
rect 2636 28549 2651 28595
rect 2575 28492 2651 28549
rect 2575 28446 2590 28492
rect 2636 28446 2651 28492
rect 2575 28389 2651 28446
rect 2575 28343 2590 28389
rect 2636 28343 2651 28389
rect 2575 28286 2651 28343
rect 2575 28240 2590 28286
rect 2636 28240 2651 28286
rect 2575 28183 2651 28240
rect 2575 28137 2590 28183
rect 2636 28137 2651 28183
rect 2575 28080 2651 28137
rect 2575 28034 2590 28080
rect 2636 28034 2651 28080
rect 2575 27976 2651 28034
rect 2575 27930 2590 27976
rect 2636 27930 2651 27976
rect 2575 27917 2651 27930
rect 2819 28904 2895 28917
rect 2819 28858 2834 28904
rect 2880 28858 2895 28904
rect 2819 28801 2895 28858
rect 2819 28755 2834 28801
rect 2880 28755 2895 28801
rect 2819 28698 2895 28755
rect 2819 28652 2834 28698
rect 2880 28652 2895 28698
rect 2819 28595 2895 28652
rect 2819 28549 2834 28595
rect 2880 28549 2895 28595
rect 2819 28492 2895 28549
rect 2819 28446 2834 28492
rect 2880 28446 2895 28492
rect 2819 28389 2895 28446
rect 2819 28343 2834 28389
rect 2880 28343 2895 28389
rect 2819 28286 2895 28343
rect 2819 28240 2834 28286
rect 2880 28240 2895 28286
rect 2819 28183 2895 28240
rect 2819 28137 2834 28183
rect 2880 28137 2895 28183
rect 2819 28080 2895 28137
rect 2819 28034 2834 28080
rect 2880 28034 2895 28080
rect 2819 27976 2895 28034
rect 2819 27930 2834 27976
rect 2880 27930 2895 27976
rect 2264 27849 2332 27860
rect 2819 27857 2895 27930
rect 3063 28904 3139 29131
rect 3063 28858 3078 28904
rect 3124 28858 3139 28904
rect 3063 28801 3139 28858
rect 3063 28755 3078 28801
rect 3124 28755 3139 28801
rect 3063 28698 3139 28755
rect 3063 28652 3078 28698
rect 3124 28652 3139 28698
rect 3063 28595 3139 28652
rect 3063 28549 3078 28595
rect 3124 28549 3139 28595
rect 3063 28492 3139 28549
rect 3063 28446 3078 28492
rect 3124 28446 3139 28492
rect 3063 28389 3139 28446
rect 3063 28343 3078 28389
rect 3124 28343 3139 28389
rect 3063 28286 3139 28343
rect 3063 28240 3078 28286
rect 3124 28240 3139 28286
rect 3063 28183 3139 28240
rect 3063 28137 3078 28183
rect 3124 28137 3139 28183
rect 3063 28080 3139 28137
rect 3063 28034 3078 28080
rect 3124 28034 3139 28080
rect 3063 27976 3139 28034
rect 3063 27930 3078 27976
rect 3124 27930 3139 27976
rect 3063 27917 3139 27930
rect 3307 28904 3383 28917
rect 3307 28858 3322 28904
rect 3368 28858 3383 28904
rect 3307 28801 3383 28858
rect 3307 28755 3322 28801
rect 3368 28755 3383 28801
rect 3307 28698 3383 28755
rect 3307 28652 3322 28698
rect 3368 28652 3383 28698
rect 3307 28595 3383 28652
rect 3307 28549 3322 28595
rect 3368 28549 3383 28595
rect 3307 28492 3383 28549
rect 3307 28446 3322 28492
rect 3368 28446 3383 28492
rect 3307 28389 3383 28446
rect 3307 28343 3322 28389
rect 3368 28343 3383 28389
rect 3307 28286 3383 28343
rect 3307 28240 3322 28286
rect 3368 28240 3383 28286
rect 3307 28183 3383 28240
rect 3307 28137 3322 28183
rect 3368 28137 3383 28183
rect 3307 28080 3383 28137
rect 3307 28034 3322 28080
rect 3368 28034 3383 28080
rect 3307 27976 3383 28034
rect 3307 27930 3322 27976
rect 3368 27930 3383 27976
rect 3307 27857 3383 27930
rect 3551 28904 3627 29131
rect 3853 29123 4115 29131
rect 3551 28858 3566 28904
rect 3612 28858 3627 28904
rect 3551 28801 3627 28858
rect 3551 28755 3566 28801
rect 3612 28755 3627 28801
rect 3551 28698 3627 28755
rect 3551 28652 3566 28698
rect 3612 28652 3627 28698
rect 3551 28595 3627 28652
rect 3551 28549 3566 28595
rect 3612 28549 3627 28595
rect 3551 28492 3627 28549
rect 3551 28446 3566 28492
rect 3612 28446 3627 28492
rect 3551 28389 3627 28446
rect 3551 28343 3566 28389
rect 3612 28343 3627 28389
rect 3551 28286 3627 28343
rect 3551 28240 3566 28286
rect 3612 28240 3627 28286
rect 3551 28183 3627 28240
rect 3551 28137 3566 28183
rect 3612 28137 3627 28183
rect 3551 28080 3627 28137
rect 3551 28034 3566 28080
rect 3612 28034 3627 28080
rect 3551 27976 3627 28034
rect 3551 27930 3566 27976
rect 3612 27930 3627 27976
rect 3551 27917 3627 27930
rect 3795 28904 3871 28917
rect 3795 28858 3810 28904
rect 3856 28858 3871 28904
rect 3795 28801 3871 28858
rect 3795 28755 3810 28801
rect 3856 28755 3871 28801
rect 3795 28698 3871 28755
rect 3795 28652 3810 28698
rect 3856 28652 3871 28698
rect 3795 28595 3871 28652
rect 3795 28549 3810 28595
rect 3856 28549 3871 28595
rect 3795 28492 3871 28549
rect 3795 28446 3810 28492
rect 3856 28446 3871 28492
rect 3795 28389 3871 28446
rect 3795 28343 3810 28389
rect 3856 28343 3871 28389
rect 3795 28286 3871 28343
rect 3795 28240 3810 28286
rect 3856 28240 3871 28286
rect 3795 28183 3871 28240
rect 3795 28137 3810 28183
rect 3856 28137 3871 28183
rect 3795 28080 3871 28137
rect 3795 28034 3810 28080
rect 3856 28034 3871 28080
rect 3795 27976 3871 28034
rect 3795 27930 3810 27976
rect 3856 27930 3871 27976
rect 3795 27857 3871 27930
rect 4039 28904 4115 29123
rect 4039 28858 4054 28904
rect 4100 28858 4115 28904
rect 4039 28801 4115 28858
rect 4039 28755 4054 28801
rect 4100 28755 4115 28801
rect 4039 28698 4115 28755
rect 4039 28652 4054 28698
rect 4100 28652 4115 28698
rect 4039 28595 4115 28652
rect 4039 28549 4054 28595
rect 4100 28549 4115 28595
rect 4039 28492 4115 28549
rect 4039 28446 4054 28492
rect 4100 28446 4115 28492
rect 4039 28389 4115 28446
rect 4039 28343 4054 28389
rect 4100 28343 4115 28389
rect 4039 28286 4115 28343
rect 4039 28240 4054 28286
rect 4100 28240 4115 28286
rect 4039 28183 4115 28240
rect 4039 28137 4054 28183
rect 4100 28137 4115 28183
rect 4039 28080 4115 28137
rect 4039 28034 4054 28080
rect 4100 28034 4115 28080
rect 4039 27976 4115 28034
rect 4039 27930 4054 27976
rect 4100 27930 4115 27976
rect 4039 27917 4115 27930
rect 4283 28904 4359 28917
rect 4283 28858 4298 28904
rect 4344 28858 4359 28904
rect 4283 28801 4359 28858
rect 4283 28755 4298 28801
rect 4344 28755 4359 28801
rect 4283 28698 4359 28755
rect 4283 28652 4298 28698
rect 4344 28652 4359 28698
rect 4283 28595 4359 28652
rect 4283 28549 4298 28595
rect 4344 28549 4359 28595
rect 4283 28492 4359 28549
rect 4283 28446 4298 28492
rect 4344 28446 4359 28492
rect 4283 28389 4359 28446
rect 4283 28343 4298 28389
rect 4344 28343 4359 28389
rect 4283 28286 4359 28343
rect 4283 28240 4298 28286
rect 4344 28240 4359 28286
rect 4283 28183 4359 28240
rect 4283 28137 4298 28183
rect 4344 28137 4359 28183
rect 4283 28080 4359 28137
rect 4283 28034 4298 28080
rect 4344 28034 4359 28080
rect 4283 27976 4359 28034
rect 4283 27930 4298 27976
rect 4344 27930 4359 27976
rect 4283 27857 4359 27930
rect 4455 28904 4531 29131
rect 4455 28858 4470 28904
rect 4516 28858 4531 28904
rect 4455 28801 4531 28858
rect 4455 28755 4470 28801
rect 4516 28755 4531 28801
rect 4455 28698 4531 28755
rect 4455 28652 4470 28698
rect 4516 28652 4531 28698
rect 4455 28595 4531 28652
rect 4455 28549 4470 28595
rect 4516 28549 4531 28595
rect 4455 28492 4531 28549
rect 4455 28446 4470 28492
rect 4516 28446 4531 28492
rect 4455 28389 4531 28446
rect 4455 28343 4470 28389
rect 4516 28343 4531 28389
rect 4455 28286 4531 28343
rect 4455 28240 4470 28286
rect 4516 28240 4531 28286
rect 4455 28183 4531 28240
rect 4455 28137 4470 28183
rect 4516 28137 4531 28183
rect 4455 28080 4531 28137
rect 4455 28034 4470 28080
rect 4516 28034 4531 28080
rect 4455 27976 4531 28034
rect 4455 27930 4470 27976
rect 4516 27930 4531 27976
rect 4455 27917 4531 27930
rect 4699 28904 4775 28917
rect 4699 28858 4714 28904
rect 4760 28858 4775 28904
rect 4699 28801 4775 28858
rect 4699 28755 4714 28801
rect 4760 28755 4775 28801
rect 4699 28698 4775 28755
rect 4699 28652 4714 28698
rect 4760 28652 4775 28698
rect 4699 28595 4775 28652
rect 4699 28549 4714 28595
rect 4760 28549 4775 28595
rect 4699 28492 4775 28549
rect 4699 28446 4714 28492
rect 4760 28446 4775 28492
rect 4699 28389 4775 28446
rect 4699 28343 4714 28389
rect 4760 28343 4775 28389
rect 4699 28286 4775 28343
rect 4699 28240 4714 28286
rect 4760 28240 4775 28286
rect 4699 28183 4775 28240
rect 4699 28137 4714 28183
rect 4760 28137 4775 28183
rect 4699 28080 4775 28137
rect 4699 28034 4714 28080
rect 4760 28034 4775 28080
rect 4699 27976 4775 28034
rect 4699 27930 4714 27976
rect 4760 27930 4775 27976
rect 2819 27781 3627 27857
rect 3795 27781 4359 27857
rect 4699 27857 4775 27930
rect 4943 28904 5019 29131
rect 4943 28858 4958 28904
rect 5004 28858 5019 28904
rect 4943 28801 5019 28858
rect 4943 28755 4958 28801
rect 5004 28755 5019 28801
rect 4943 28698 5019 28755
rect 4943 28652 4958 28698
rect 5004 28652 5019 28698
rect 4943 28595 5019 28652
rect 4943 28549 4958 28595
rect 5004 28549 5019 28595
rect 4943 28492 5019 28549
rect 4943 28446 4958 28492
rect 5004 28446 5019 28492
rect 4943 28389 5019 28446
rect 4943 28343 4958 28389
rect 5004 28343 5019 28389
rect 4943 28286 5019 28343
rect 4943 28240 4958 28286
rect 5004 28240 5019 28286
rect 4943 28183 5019 28240
rect 4943 28137 4958 28183
rect 5004 28137 5019 28183
rect 4943 28080 5019 28137
rect 4943 28034 4958 28080
rect 5004 28034 5019 28080
rect 4943 27976 5019 28034
rect 4943 27930 4958 27976
rect 5004 27930 5019 27976
rect 4943 27917 5019 27930
rect 5187 28904 5263 28917
rect 5187 28858 5202 28904
rect 5248 28858 5263 28904
rect 5187 28801 5263 28858
rect 5187 28755 5202 28801
rect 5248 28755 5263 28801
rect 5187 28698 5263 28755
rect 5187 28652 5202 28698
rect 5248 28652 5263 28698
rect 5187 28595 5263 28652
rect 5187 28549 5202 28595
rect 5248 28549 5263 28595
rect 5187 28492 5263 28549
rect 5187 28446 5202 28492
rect 5248 28446 5263 28492
rect 5187 28389 5263 28446
rect 5187 28343 5202 28389
rect 5248 28343 5263 28389
rect 5187 28286 5263 28343
rect 5187 28240 5202 28286
rect 5248 28240 5263 28286
rect 5187 28183 5263 28240
rect 5187 28137 5202 28183
rect 5248 28137 5263 28183
rect 5187 28080 5263 28137
rect 5187 28034 5202 28080
rect 5248 28034 5263 28080
rect 5187 27976 5263 28034
rect 5187 27930 5202 27976
rect 5248 27930 5263 27976
rect 5187 27857 5263 27930
rect 5431 28904 5507 29131
rect 5431 28858 5446 28904
rect 5492 28858 5507 28904
rect 5431 28801 5507 28858
rect 5431 28755 5446 28801
rect 5492 28755 5507 28801
rect 5431 28698 5507 28755
rect 5431 28652 5446 28698
rect 5492 28652 5507 28698
rect 5431 28595 5507 28652
rect 5431 28549 5446 28595
rect 5492 28549 5507 28595
rect 5431 28492 5507 28549
rect 5431 28446 5446 28492
rect 5492 28446 5507 28492
rect 5431 28389 5507 28446
rect 5431 28343 5446 28389
rect 5492 28343 5507 28389
rect 5431 28286 5507 28343
rect 5431 28240 5446 28286
rect 5492 28240 5507 28286
rect 5431 28183 5507 28240
rect 5431 28137 5446 28183
rect 5492 28137 5507 28183
rect 5431 28080 5507 28137
rect 5431 28034 5446 28080
rect 5492 28034 5507 28080
rect 5431 27976 5507 28034
rect 5431 27930 5446 27976
rect 5492 27930 5507 27976
rect 5431 27917 5507 27930
rect 5675 28904 5751 28917
rect 5675 28858 5690 28904
rect 5736 28858 5751 28904
rect 5675 28801 5751 28858
rect 5675 28755 5690 28801
rect 5736 28755 5751 28801
rect 5675 28698 5751 28755
rect 5675 28652 5690 28698
rect 5736 28652 5751 28698
rect 5675 28595 5751 28652
rect 5675 28549 5690 28595
rect 5736 28549 5751 28595
rect 5675 28492 5751 28549
rect 5675 28446 5690 28492
rect 5736 28446 5751 28492
rect 5675 28389 5751 28446
rect 5675 28343 5690 28389
rect 5736 28343 5751 28389
rect 5675 28286 5751 28343
rect 5675 28240 5690 28286
rect 5736 28240 5751 28286
rect 5675 28183 5751 28240
rect 5675 28137 5690 28183
rect 5736 28137 5751 28183
rect 5675 28080 5751 28137
rect 5675 28034 5690 28080
rect 5736 28034 5751 28080
rect 5675 27976 5751 28034
rect 5675 27930 5690 27976
rect 5736 27930 5751 27976
rect 5675 27857 5751 27930
rect 5919 28904 5995 29131
rect 6235 29123 6727 29131
rect 5919 28858 5934 28904
rect 5980 28858 5995 28904
rect 5919 28801 5995 28858
rect 5919 28755 5934 28801
rect 5980 28755 5995 28801
rect 5919 28698 5995 28755
rect 5919 28652 5934 28698
rect 5980 28652 5995 28698
rect 5919 28595 5995 28652
rect 5919 28549 5934 28595
rect 5980 28549 5995 28595
rect 5919 28492 5995 28549
rect 5919 28446 5934 28492
rect 5980 28446 5995 28492
rect 5919 28389 5995 28446
rect 5919 28343 5934 28389
rect 5980 28343 5995 28389
rect 5919 28286 5995 28343
rect 5919 28240 5934 28286
rect 5980 28240 5995 28286
rect 5919 28183 5995 28240
rect 5919 28137 5934 28183
rect 5980 28137 5995 28183
rect 5919 28080 5995 28137
rect 5919 28034 5934 28080
rect 5980 28034 5995 28080
rect 5919 27976 5995 28034
rect 5919 27930 5934 27976
rect 5980 27930 5995 27976
rect 5919 27917 5995 27930
rect 6163 28904 6239 28917
rect 6163 28858 6178 28904
rect 6224 28858 6239 28904
rect 6163 28801 6239 28858
rect 6163 28755 6178 28801
rect 6224 28755 6239 28801
rect 6163 28698 6239 28755
rect 6163 28652 6178 28698
rect 6224 28652 6239 28698
rect 6163 28595 6239 28652
rect 6163 28549 6178 28595
rect 6224 28549 6239 28595
rect 6163 28492 6239 28549
rect 6163 28446 6178 28492
rect 6224 28446 6239 28492
rect 6163 28389 6239 28446
rect 6163 28343 6178 28389
rect 6224 28343 6239 28389
rect 6163 28286 6239 28343
rect 6163 28240 6178 28286
rect 6224 28240 6239 28286
rect 6163 28183 6239 28240
rect 6163 28137 6178 28183
rect 6224 28137 6239 28183
rect 6163 28080 6239 28137
rect 6163 28034 6178 28080
rect 6224 28034 6239 28080
rect 6163 27976 6239 28034
rect 6163 27930 6178 27976
rect 6224 27930 6239 27976
rect 6163 27857 6239 27930
rect 6407 28904 6483 29123
rect 6407 28858 6422 28904
rect 6468 28858 6483 28904
rect 6407 28801 6483 28858
rect 6407 28755 6422 28801
rect 6468 28755 6483 28801
rect 6407 28698 6483 28755
rect 6407 28652 6422 28698
rect 6468 28652 6483 28698
rect 6407 28595 6483 28652
rect 6407 28549 6422 28595
rect 6468 28549 6483 28595
rect 6407 28492 6483 28549
rect 6407 28446 6422 28492
rect 6468 28446 6483 28492
rect 6407 28389 6483 28446
rect 6407 28343 6422 28389
rect 6468 28343 6483 28389
rect 6407 28286 6483 28343
rect 6407 28240 6422 28286
rect 6468 28240 6483 28286
rect 6407 28183 6483 28240
rect 6407 28137 6422 28183
rect 6468 28137 6483 28183
rect 6407 28080 6483 28137
rect 6407 28034 6422 28080
rect 6468 28034 6483 28080
rect 6407 27976 6483 28034
rect 6407 27930 6422 27976
rect 6468 27930 6483 27976
rect 6407 27917 6483 27930
rect 6651 28904 6727 28917
rect 6651 28858 6666 28904
rect 6712 28858 6727 28904
rect 6651 28801 6727 28858
rect 6651 28755 6666 28801
rect 6712 28755 6727 28801
rect 6651 28698 6727 28755
rect 6651 28652 6666 28698
rect 6712 28652 6727 28698
rect 6651 28595 6727 28652
rect 6651 28549 6666 28595
rect 6712 28549 6727 28595
rect 6651 28492 6727 28549
rect 6651 28446 6666 28492
rect 6712 28446 6727 28492
rect 6651 28389 6727 28446
rect 6651 28343 6666 28389
rect 6712 28343 6727 28389
rect 6651 28286 6727 28343
rect 6651 28240 6666 28286
rect 6712 28240 6727 28286
rect 6651 28183 6727 28240
rect 6651 28137 6666 28183
rect 6712 28137 6727 28183
rect 6651 28080 6727 28137
rect 6651 28034 6666 28080
rect 6712 28034 6727 28080
rect 6651 27976 6727 28034
rect 6651 27930 6666 27976
rect 6712 27930 6727 27976
rect 6651 27857 6727 27930
rect 6895 28904 6971 29131
rect 6895 28858 6910 28904
rect 6956 28858 6971 28904
rect 6895 28801 6971 28858
rect 6895 28755 6910 28801
rect 6956 28755 6971 28801
rect 6895 28698 6971 28755
rect 6895 28652 6910 28698
rect 6956 28652 6971 28698
rect 6895 28595 6971 28652
rect 6895 28549 6910 28595
rect 6956 28549 6971 28595
rect 6895 28492 6971 28549
rect 6895 28446 6910 28492
rect 6956 28446 6971 28492
rect 6895 28389 6971 28446
rect 6895 28343 6910 28389
rect 6956 28343 6971 28389
rect 6895 28286 6971 28343
rect 6895 28240 6910 28286
rect 6956 28240 6971 28286
rect 6895 28183 6971 28240
rect 6895 28137 6910 28183
rect 6956 28137 6971 28183
rect 6895 28080 6971 28137
rect 6895 28034 6910 28080
rect 6956 28034 6971 28080
rect 6895 27976 6971 28034
rect 6895 27930 6910 27976
rect 6956 27930 6971 27976
rect 6895 27917 6971 27930
rect 7139 28904 7215 28917
rect 7139 28858 7154 28904
rect 7200 28858 7215 28904
rect 7139 28801 7215 28858
rect 7139 28755 7154 28801
rect 7200 28755 7215 28801
rect 7139 28698 7215 28755
rect 7139 28652 7154 28698
rect 7200 28652 7215 28698
rect 7139 28595 7215 28652
rect 7139 28549 7154 28595
rect 7200 28549 7215 28595
rect 7139 28492 7215 28549
rect 7139 28446 7154 28492
rect 7200 28446 7215 28492
rect 7139 28389 7215 28446
rect 7139 28343 7154 28389
rect 7200 28343 7215 28389
rect 7139 28286 7215 28343
rect 7139 28240 7154 28286
rect 7200 28240 7215 28286
rect 7139 28183 7215 28240
rect 7139 28137 7154 28183
rect 7200 28137 7215 28183
rect 7139 28080 7215 28137
rect 7139 28034 7154 28080
rect 7200 28034 7215 28080
rect 7139 27976 7215 28034
rect 7139 27930 7154 27976
rect 7200 27930 7215 27976
rect 7139 27857 7215 27930
rect 7383 28904 7459 29131
rect 7383 28858 7398 28904
rect 7444 28858 7459 28904
rect 7383 28801 7459 28858
rect 7383 28755 7398 28801
rect 7444 28755 7459 28801
rect 7383 28698 7459 28755
rect 7383 28652 7398 28698
rect 7444 28652 7459 28698
rect 7383 28595 7459 28652
rect 7383 28549 7398 28595
rect 7444 28549 7459 28595
rect 7383 28492 7459 28549
rect 7383 28446 7398 28492
rect 7444 28446 7459 28492
rect 7383 28389 7459 28446
rect 7383 28343 7398 28389
rect 7444 28343 7459 28389
rect 7383 28286 7459 28343
rect 7383 28240 7398 28286
rect 7444 28240 7459 28286
rect 7383 28183 7459 28240
rect 7383 28137 7398 28183
rect 7444 28137 7459 28183
rect 7383 28080 7459 28137
rect 7383 28034 7398 28080
rect 7444 28034 7459 28080
rect 7383 27976 7459 28034
rect 7383 27930 7398 27976
rect 7444 27930 7459 27976
rect 7383 27917 7459 27930
rect 7627 28904 7703 28917
rect 7627 28858 7642 28904
rect 7688 28858 7703 28904
rect 7627 28801 7703 28858
rect 7627 28755 7642 28801
rect 7688 28755 7703 28801
rect 7627 28698 7703 28755
rect 7627 28652 7642 28698
rect 7688 28652 7703 28698
rect 7627 28595 7703 28652
rect 7627 28549 7642 28595
rect 7688 28549 7703 28595
rect 7627 28492 7703 28549
rect 7627 28446 7642 28492
rect 7688 28446 7703 28492
rect 7627 28389 7703 28446
rect 7627 28343 7642 28389
rect 7688 28343 7703 28389
rect 7627 28286 7703 28343
rect 7627 28240 7642 28286
rect 7688 28240 7703 28286
rect 7627 28183 7703 28240
rect 7627 28137 7642 28183
rect 7688 28137 7703 28183
rect 7627 28080 7703 28137
rect 7627 28034 7642 28080
rect 7688 28034 7703 28080
rect 7627 27976 7703 28034
rect 7627 27930 7642 27976
rect 7688 27930 7703 27976
rect 7627 27857 7703 27930
rect 7871 28904 7947 29131
rect 7871 28858 7886 28904
rect 7932 28858 7947 28904
rect 7871 28801 7947 28858
rect 7871 28755 7886 28801
rect 7932 28755 7947 28801
rect 7871 28698 7947 28755
rect 7871 28652 7886 28698
rect 7932 28652 7947 28698
rect 7871 28595 7947 28652
rect 7871 28549 7886 28595
rect 7932 28549 7947 28595
rect 7871 28492 7947 28549
rect 7871 28446 7886 28492
rect 7932 28446 7947 28492
rect 7871 28389 7947 28446
rect 7871 28343 7886 28389
rect 7932 28343 7947 28389
rect 7871 28286 7947 28343
rect 7871 28240 7886 28286
rect 7932 28240 7947 28286
rect 7871 28183 7947 28240
rect 7871 28137 7886 28183
rect 7932 28137 7947 28183
rect 7871 28080 7947 28137
rect 7871 28034 7886 28080
rect 7932 28034 7947 28080
rect 7871 27976 7947 28034
rect 7871 27930 7886 27976
rect 7932 27930 7947 27976
rect 7871 27917 7947 27930
rect 8115 28904 8191 28917
rect 8115 28858 8130 28904
rect 8176 28858 8191 28904
rect 8115 28801 8191 28858
rect 8115 28755 8130 28801
rect 8176 28755 8191 28801
rect 8115 28698 8191 28755
rect 8115 28652 8130 28698
rect 8176 28652 8191 28698
rect 8115 28595 8191 28652
rect 8115 28549 8130 28595
rect 8176 28549 8191 28595
rect 8115 28492 8191 28549
rect 8115 28446 8130 28492
rect 8176 28446 8191 28492
rect 8115 28389 8191 28446
rect 8115 28343 8130 28389
rect 8176 28343 8191 28389
rect 8115 28286 8191 28343
rect 8115 28240 8130 28286
rect 8176 28240 8191 28286
rect 8115 28183 8191 28240
rect 8115 28137 8130 28183
rect 8176 28137 8191 28183
rect 8115 28080 8191 28137
rect 8115 28034 8130 28080
rect 8176 28034 8191 28080
rect 8115 27976 8191 28034
rect 8115 27930 8130 27976
rect 8176 27930 8191 27976
rect 8115 27857 8191 27930
rect 8359 28904 8435 29131
rect 8847 29123 9109 29131
rect 8359 28858 8374 28904
rect 8420 28858 8435 28904
rect 8359 28801 8435 28858
rect 8359 28755 8374 28801
rect 8420 28755 8435 28801
rect 8359 28698 8435 28755
rect 8359 28652 8374 28698
rect 8420 28652 8435 28698
rect 8359 28595 8435 28652
rect 8359 28549 8374 28595
rect 8420 28549 8435 28595
rect 8359 28492 8435 28549
rect 8359 28446 8374 28492
rect 8420 28446 8435 28492
rect 8359 28389 8435 28446
rect 8359 28343 8374 28389
rect 8420 28343 8435 28389
rect 8359 28286 8435 28343
rect 8359 28240 8374 28286
rect 8420 28240 8435 28286
rect 8359 28183 8435 28240
rect 8359 28137 8374 28183
rect 8420 28137 8435 28183
rect 8359 28080 8435 28137
rect 8359 28034 8374 28080
rect 8420 28034 8435 28080
rect 8359 27976 8435 28034
rect 8359 27930 8374 27976
rect 8420 27930 8435 27976
rect 8359 27917 8435 27930
rect 8603 28904 8679 28917
rect 8603 28858 8618 28904
rect 8664 28858 8679 28904
rect 8603 28801 8679 28858
rect 8603 28755 8618 28801
rect 8664 28755 8679 28801
rect 8603 28698 8679 28755
rect 8603 28652 8618 28698
rect 8664 28652 8679 28698
rect 8603 28595 8679 28652
rect 8603 28549 8618 28595
rect 8664 28549 8679 28595
rect 8603 28492 8679 28549
rect 8603 28446 8618 28492
rect 8664 28446 8679 28492
rect 8603 28389 8679 28446
rect 8603 28343 8618 28389
rect 8664 28343 8679 28389
rect 8603 28286 8679 28343
rect 8603 28240 8618 28286
rect 8664 28240 8679 28286
rect 8603 28183 8679 28240
rect 8603 28137 8618 28183
rect 8664 28137 8679 28183
rect 8603 28080 8679 28137
rect 8603 28034 8618 28080
rect 8664 28034 8679 28080
rect 8603 27976 8679 28034
rect 8603 27930 8618 27976
rect 8664 27930 8679 27976
rect 8603 27857 8679 27930
rect 8847 28904 8923 29123
rect 8847 28858 8862 28904
rect 8908 28858 8923 28904
rect 8847 28801 8923 28858
rect 8847 28755 8862 28801
rect 8908 28755 8923 28801
rect 8847 28698 8923 28755
rect 8847 28652 8862 28698
rect 8908 28652 8923 28698
rect 8847 28595 8923 28652
rect 8847 28549 8862 28595
rect 8908 28549 8923 28595
rect 8847 28492 8923 28549
rect 8847 28446 8862 28492
rect 8908 28446 8923 28492
rect 8847 28389 8923 28446
rect 8847 28343 8862 28389
rect 8908 28343 8923 28389
rect 8847 28286 8923 28343
rect 8847 28240 8862 28286
rect 8908 28240 8923 28286
rect 8847 28183 8923 28240
rect 8847 28137 8862 28183
rect 8908 28137 8923 28183
rect 8847 28080 8923 28137
rect 8847 28034 8862 28080
rect 8908 28034 8923 28080
rect 8847 27976 8923 28034
rect 8847 27930 8862 27976
rect 8908 27930 8923 27976
rect 8847 27917 8923 27930
rect 9091 28904 9167 28917
rect 9091 28858 9106 28904
rect 9152 28858 9167 28904
rect 9091 28801 9167 28858
rect 9091 28755 9106 28801
rect 9152 28755 9167 28801
rect 9091 28698 9167 28755
rect 9091 28652 9106 28698
rect 9152 28652 9167 28698
rect 9091 28595 9167 28652
rect 9091 28549 9106 28595
rect 9152 28549 9167 28595
rect 9091 28492 9167 28549
rect 9091 28446 9106 28492
rect 9152 28446 9167 28492
rect 9091 28389 9167 28446
rect 9091 28343 9106 28389
rect 9152 28343 9167 28389
rect 9091 28286 9167 28343
rect 9091 28240 9106 28286
rect 9152 28240 9167 28286
rect 9091 28183 9167 28240
rect 9091 28137 9106 28183
rect 9152 28137 9167 28183
rect 9091 28080 9167 28137
rect 9091 28034 9106 28080
rect 9152 28034 9167 28080
rect 9091 27976 9167 28034
rect 9091 27930 9106 27976
rect 9152 27930 9167 27976
rect 9091 27857 9167 27930
rect 9335 28904 9411 29131
rect 9335 28858 9350 28904
rect 9396 28858 9411 28904
rect 9335 28801 9411 28858
rect 9335 28755 9350 28801
rect 9396 28755 9411 28801
rect 9335 28698 9411 28755
rect 9335 28652 9350 28698
rect 9396 28652 9411 28698
rect 9335 28595 9411 28652
rect 9335 28549 9350 28595
rect 9396 28549 9411 28595
rect 9335 28492 9411 28549
rect 9335 28446 9350 28492
rect 9396 28446 9411 28492
rect 9335 28389 9411 28446
rect 9335 28343 9350 28389
rect 9396 28343 9411 28389
rect 9335 28286 9411 28343
rect 9335 28240 9350 28286
rect 9396 28240 9411 28286
rect 9335 28183 9411 28240
rect 9335 28137 9350 28183
rect 9396 28137 9411 28183
rect 9335 28080 9411 28137
rect 9335 28034 9350 28080
rect 9396 28034 9411 28080
rect 9335 27976 9411 28034
rect 9335 27930 9350 27976
rect 9396 27930 9411 27976
rect 9335 27917 9411 27930
rect 9579 28904 9655 28917
rect 9579 28858 9594 28904
rect 9640 28858 9655 28904
rect 9579 28801 9655 28858
rect 9579 28755 9594 28801
rect 9640 28755 9655 28801
rect 9579 28698 9655 28755
rect 9579 28652 9594 28698
rect 9640 28652 9655 28698
rect 9579 28595 9655 28652
rect 9579 28549 9594 28595
rect 9640 28549 9655 28595
rect 9579 28492 9655 28549
rect 9579 28446 9594 28492
rect 9640 28446 9655 28492
rect 9579 28389 9655 28446
rect 9579 28343 9594 28389
rect 9640 28343 9655 28389
rect 9579 28286 9655 28343
rect 9579 28240 9594 28286
rect 9640 28240 9655 28286
rect 9579 28183 9655 28240
rect 9579 28137 9594 28183
rect 9640 28137 9655 28183
rect 9579 28080 9655 28137
rect 9579 28034 9594 28080
rect 9640 28034 9655 28080
rect 9579 27976 9655 28034
rect 9579 27930 9594 27976
rect 9640 27930 9655 27976
rect 9579 27857 9655 27930
rect 9823 28904 9899 29131
rect 9823 28858 9838 28904
rect 9884 28858 9899 28904
rect 9823 28801 9899 28858
rect 9823 28755 9838 28801
rect 9884 28755 9899 28801
rect 9823 28698 9899 28755
rect 9823 28652 9838 28698
rect 9884 28652 9899 28698
rect 9823 28595 9899 28652
rect 9823 28549 9838 28595
rect 9884 28549 9899 28595
rect 9823 28492 9899 28549
rect 9823 28446 9838 28492
rect 9884 28446 9899 28492
rect 9823 28389 9899 28446
rect 9823 28343 9838 28389
rect 9884 28343 9899 28389
rect 9823 28286 9899 28343
rect 9823 28240 9838 28286
rect 9884 28240 9899 28286
rect 9823 28183 9899 28240
rect 9823 28137 9838 28183
rect 9884 28137 9899 28183
rect 9823 28080 9899 28137
rect 9823 28034 9838 28080
rect 9884 28034 9899 28080
rect 9823 27976 9899 28034
rect 9823 27930 9838 27976
rect 9884 27930 9899 27976
rect 9823 27917 9899 27930
rect 10067 28904 10143 28917
rect 10067 28858 10082 28904
rect 10128 28858 10143 28904
rect 10067 28801 10143 28858
rect 10067 28755 10082 28801
rect 10128 28755 10143 28801
rect 10067 28698 10143 28755
rect 10067 28652 10082 28698
rect 10128 28652 10143 28698
rect 10067 28595 10143 28652
rect 10067 28549 10082 28595
rect 10128 28549 10143 28595
rect 10067 28492 10143 28549
rect 10067 28446 10082 28492
rect 10128 28446 10143 28492
rect 10067 28389 10143 28446
rect 10067 28343 10082 28389
rect 10128 28343 10143 28389
rect 10067 28286 10143 28343
rect 10067 28240 10082 28286
rect 10128 28240 10143 28286
rect 10067 28183 10143 28240
rect 10067 28137 10082 28183
rect 10128 28137 10143 28183
rect 10067 28080 10143 28137
rect 10067 28034 10082 28080
rect 10128 28034 10143 28080
rect 10067 27976 10143 28034
rect 10067 27930 10082 27976
rect 10128 27930 10143 27976
rect 10067 27857 10143 27930
rect 10311 28904 10387 29131
rect 10311 28858 10326 28904
rect 10372 28858 10387 28904
rect 10311 28801 10387 28858
rect 10311 28755 10326 28801
rect 10372 28755 10387 28801
rect 10311 28698 10387 28755
rect 10311 28652 10326 28698
rect 10372 28652 10387 28698
rect 10311 28595 10387 28652
rect 10311 28549 10326 28595
rect 10372 28549 10387 28595
rect 10311 28492 10387 28549
rect 10311 28446 10326 28492
rect 10372 28446 10387 28492
rect 10311 28389 10387 28446
rect 10311 28343 10326 28389
rect 10372 28343 10387 28389
rect 10311 28286 10387 28343
rect 10311 28240 10326 28286
rect 10372 28240 10387 28286
rect 10311 28183 10387 28240
rect 10311 28137 10326 28183
rect 10372 28137 10387 28183
rect 10311 28080 10387 28137
rect 10311 28034 10326 28080
rect 10372 28034 10387 28080
rect 10311 27976 10387 28034
rect 10311 27930 10326 27976
rect 10372 27930 10387 27976
rect 10311 27917 10387 27930
rect 10630 29123 11489 29131
rect 10630 29034 10698 29123
rect 10630 27860 10641 29034
rect 10687 27860 10698 29034
rect 4699 27781 10433 27857
rect 10630 27849 10698 27860
rect 3551 27725 3627 27781
rect -50 27710 3464 27721
rect -50 27664 2749 27710
rect 3453 27664 3464 27710
rect -50 27521 3464 27664
rect 2264 27156 2340 27167
rect 2264 25888 2275 27156
rect 2321 27155 2340 27156
rect 2328 25959 2340 27155
rect 3388 27146 3464 27521
rect 3551 27710 4224 27725
rect 3551 27664 3697 27710
rect 4213 27664 4224 27710
rect 3551 27649 4224 27664
rect 4283 27721 4359 27781
rect 4283 27710 10275 27721
rect 4283 27664 4578 27710
rect 10264 27664 10275 27710
rect 3551 27274 3627 27649
rect 4283 27645 10275 27664
rect 3737 27485 6531 27496
rect 3737 27439 3748 27485
rect 6520 27439 6531 27485
rect 3737 27432 4166 27439
rect 6090 27432 6531 27439
rect 3737 27428 6531 27432
rect 4154 27420 6102 27428
rect 3551 27259 6516 27274
rect 3551 27213 5237 27259
rect 6505 27213 6516 27259
rect 3551 27198 6516 27213
rect 6652 27270 6728 27645
rect 6860 27485 10236 27496
rect 6860 27484 6889 27485
rect 6860 27432 6872 27484
rect 10225 27439 10236 27485
rect 8796 27432 9236 27439
rect 10224 27432 10236 27439
rect 6860 27428 10236 27432
rect 6860 27420 8808 27428
rect 9224 27420 10236 27428
rect 6652 27259 7980 27270
rect 6652 27213 6701 27259
rect 7969 27213 7980 27259
rect 6652 27202 7980 27213
rect 3388 27131 4223 27146
rect 3388 27085 4072 27131
rect 4212 27085 4223 27131
rect 3388 27070 4223 27085
rect 2321 25947 2340 25959
rect 4039 26993 4115 27006
rect 4039 26947 4054 26993
rect 4100 26947 4115 26993
rect 4039 26890 4115 26947
rect 4039 26844 4054 26890
rect 4100 26844 4115 26890
rect 4039 26787 4115 26844
rect 4039 26741 4054 26787
rect 4100 26741 4115 26787
rect 4039 26684 4115 26741
rect 4039 26638 4054 26684
rect 4100 26638 4115 26684
rect 4039 26581 4115 26638
rect 4039 26535 4054 26581
rect 4100 26535 4115 26581
rect 4039 26478 4115 26535
rect 4039 26432 4054 26478
rect 4100 26432 4115 26478
rect 4039 26375 4115 26432
rect 4039 26329 4054 26375
rect 4100 26329 4115 26375
rect 4039 26272 4115 26329
rect 4039 26226 4054 26272
rect 4100 26226 4115 26272
rect 4039 26169 4115 26226
rect 4039 26123 4054 26169
rect 4100 26123 4115 26169
rect 4039 26065 4115 26123
rect 4039 26019 4054 26065
rect 4100 26019 4115 26065
rect 2321 25888 2332 25947
rect 2264 25791 2332 25888
rect 4039 25799 4115 26019
rect 4283 26993 4359 27198
rect 6652 27142 6728 27202
rect 10357 27142 10433 27781
rect 5345 27066 6728 27142
rect 6809 27066 10433 27142
rect 10622 27156 10698 27167
rect 10622 27155 10641 27156
rect 4283 26947 4298 26993
rect 4344 26947 4359 26993
rect 4283 26890 4359 26947
rect 4283 26844 4298 26890
rect 4344 26844 4359 26890
rect 4283 26787 4359 26844
rect 4283 26741 4298 26787
rect 4344 26741 4359 26787
rect 4283 26684 4359 26741
rect 4283 26638 4298 26684
rect 4344 26638 4359 26684
rect 4283 26581 4359 26638
rect 4283 26535 4298 26581
rect 4344 26535 4359 26581
rect 4283 26478 4359 26535
rect 4283 26432 4298 26478
rect 4344 26432 4359 26478
rect 4283 26375 4359 26432
rect 4283 26329 4298 26375
rect 4344 26329 4359 26375
rect 4283 26272 4359 26329
rect 4283 26226 4298 26272
rect 4344 26226 4359 26272
rect 4283 26169 4359 26226
rect 4283 26123 4298 26169
rect 4344 26123 4359 26169
rect 4283 26065 4359 26123
rect 4283 26019 4298 26065
rect 4344 26019 4359 26065
rect 4283 26006 4359 26019
rect 5101 26993 5177 27006
rect 5101 26947 5116 26993
rect 5162 26947 5177 26993
rect 5101 26890 5177 26947
rect 5101 26844 5116 26890
rect 5162 26844 5177 26890
rect 5101 26787 5177 26844
rect 5101 26741 5116 26787
rect 5162 26741 5177 26787
rect 5101 26684 5177 26741
rect 5101 26638 5116 26684
rect 5162 26638 5177 26684
rect 5101 26581 5177 26638
rect 5101 26535 5116 26581
rect 5162 26535 5177 26581
rect 5101 26478 5177 26535
rect 5101 26432 5116 26478
rect 5162 26432 5177 26478
rect 5101 26375 5177 26432
rect 5101 26329 5116 26375
rect 5162 26329 5177 26375
rect 5101 26272 5177 26329
rect 5101 26226 5116 26272
rect 5162 26226 5177 26272
rect 5101 26169 5177 26226
rect 5101 26123 5116 26169
rect 5162 26123 5177 26169
rect 5101 26065 5177 26123
rect 5101 26019 5116 26065
rect 5162 26019 5177 26065
rect 4033 25791 4115 25799
rect 5101 25791 5177 26019
rect 5345 26993 5421 27066
rect 5345 26947 5360 26993
rect 5406 26947 5421 26993
rect 5345 26890 5421 26947
rect 5345 26844 5360 26890
rect 5406 26844 5421 26890
rect 5345 26787 5421 26844
rect 5345 26741 5360 26787
rect 5406 26741 5421 26787
rect 5345 26684 5421 26741
rect 5345 26638 5360 26684
rect 5406 26638 5421 26684
rect 5345 26581 5421 26638
rect 5345 26535 5360 26581
rect 5406 26535 5421 26581
rect 5345 26478 5421 26535
rect 5345 26432 5360 26478
rect 5406 26432 5421 26478
rect 5345 26375 5421 26432
rect 5345 26329 5360 26375
rect 5406 26329 5421 26375
rect 5345 26272 5421 26329
rect 5345 26226 5360 26272
rect 5406 26226 5421 26272
rect 5345 26169 5421 26226
rect 5345 26123 5360 26169
rect 5406 26123 5421 26169
rect 5345 26065 5421 26123
rect 5345 26019 5360 26065
rect 5406 26019 5421 26065
rect 5345 26006 5421 26019
rect 5589 26993 5665 27006
rect 5589 26947 5604 26993
rect 5650 26947 5665 26993
rect 5589 26890 5665 26947
rect 5589 26844 5604 26890
rect 5650 26844 5665 26890
rect 5589 26787 5665 26844
rect 5589 26741 5604 26787
rect 5650 26741 5665 26787
rect 5589 26684 5665 26741
rect 5589 26638 5604 26684
rect 5650 26638 5665 26684
rect 5589 26581 5665 26638
rect 5589 26535 5604 26581
rect 5650 26535 5665 26581
rect 5589 26478 5665 26535
rect 5589 26432 5604 26478
rect 5650 26432 5665 26478
rect 5589 26375 5665 26432
rect 5589 26329 5604 26375
rect 5650 26329 5665 26375
rect 5589 26272 5665 26329
rect 5589 26226 5604 26272
rect 5650 26226 5665 26272
rect 5589 26169 5665 26226
rect 5589 26123 5604 26169
rect 5650 26123 5665 26169
rect 5589 26065 5665 26123
rect 5589 26019 5604 26065
rect 5650 26019 5665 26065
rect 5589 25791 5665 26019
rect 5833 26993 5909 27066
rect 5833 26947 5848 26993
rect 5894 26947 5909 26993
rect 5833 26890 5909 26947
rect 5833 26844 5848 26890
rect 5894 26844 5909 26890
rect 5833 26787 5909 26844
rect 5833 26741 5848 26787
rect 5894 26741 5909 26787
rect 5833 26684 5909 26741
rect 5833 26638 5848 26684
rect 5894 26638 5909 26684
rect 5833 26581 5909 26638
rect 5833 26535 5848 26581
rect 5894 26535 5909 26581
rect 5833 26478 5909 26535
rect 5833 26432 5848 26478
rect 5894 26432 5909 26478
rect 5833 26375 5909 26432
rect 5833 26329 5848 26375
rect 5894 26329 5909 26375
rect 5833 26272 5909 26329
rect 5833 26226 5848 26272
rect 5894 26226 5909 26272
rect 5833 26169 5909 26226
rect 5833 26123 5848 26169
rect 5894 26123 5909 26169
rect 5833 26065 5909 26123
rect 5833 26019 5848 26065
rect 5894 26019 5909 26065
rect 5833 26006 5909 26019
rect 6077 26993 6153 27006
rect 6077 26947 6092 26993
rect 6138 26947 6153 26993
rect 6077 26890 6153 26947
rect 6077 26844 6092 26890
rect 6138 26844 6153 26890
rect 6077 26787 6153 26844
rect 6077 26741 6092 26787
rect 6138 26741 6153 26787
rect 6077 26684 6153 26741
rect 6077 26638 6092 26684
rect 6138 26638 6153 26684
rect 6077 26581 6153 26638
rect 6077 26535 6092 26581
rect 6138 26535 6153 26581
rect 6077 26478 6153 26535
rect 6077 26432 6092 26478
rect 6138 26432 6153 26478
rect 6077 26375 6153 26432
rect 6077 26329 6092 26375
rect 6138 26329 6153 26375
rect 6077 26272 6153 26329
rect 6077 26226 6092 26272
rect 6138 26226 6153 26272
rect 6077 26169 6153 26226
rect 6077 26123 6092 26169
rect 6138 26123 6153 26169
rect 6077 26065 6153 26123
rect 6077 26019 6092 26065
rect 6138 26019 6153 26065
rect 6077 25791 6153 26019
rect 6321 26993 6397 27066
rect 6321 26947 6336 26993
rect 6382 26947 6397 26993
rect 6321 26890 6397 26947
rect 6321 26844 6336 26890
rect 6382 26844 6397 26890
rect 6321 26787 6397 26844
rect 6321 26741 6336 26787
rect 6382 26741 6397 26787
rect 6321 26684 6397 26741
rect 6321 26638 6336 26684
rect 6382 26638 6397 26684
rect 6321 26581 6397 26638
rect 6321 26535 6336 26581
rect 6382 26535 6397 26581
rect 6321 26478 6397 26535
rect 6321 26432 6336 26478
rect 6382 26432 6397 26478
rect 6321 26375 6397 26432
rect 6321 26329 6336 26375
rect 6382 26329 6397 26375
rect 6321 26272 6397 26329
rect 6321 26226 6336 26272
rect 6382 26226 6397 26272
rect 6321 26169 6397 26226
rect 6321 26123 6336 26169
rect 6382 26123 6397 26169
rect 6321 26065 6397 26123
rect 6321 26019 6336 26065
rect 6382 26019 6397 26065
rect 6321 26006 6397 26019
rect 6565 26993 6641 27006
rect 6565 26947 6580 26993
rect 6626 26947 6641 26993
rect 6565 26890 6641 26947
rect 6565 26844 6580 26890
rect 6626 26844 6641 26890
rect 6565 26787 6641 26844
rect 6565 26741 6580 26787
rect 6626 26741 6641 26787
rect 6565 26684 6641 26741
rect 6565 26638 6580 26684
rect 6626 26638 6641 26684
rect 6565 26581 6641 26638
rect 6565 26535 6580 26581
rect 6626 26535 6641 26581
rect 6565 26478 6641 26535
rect 6565 26432 6580 26478
rect 6626 26432 6641 26478
rect 6565 26375 6641 26432
rect 6565 26329 6580 26375
rect 6626 26329 6641 26375
rect 6565 26272 6641 26329
rect 6565 26226 6580 26272
rect 6626 26226 6641 26272
rect 6565 26169 6641 26226
rect 6565 26123 6580 26169
rect 6626 26123 6641 26169
rect 6565 26065 6641 26123
rect 6565 26019 6580 26065
rect 6626 26019 6641 26065
rect 6565 25791 6641 26019
rect 6809 26993 6885 27066
rect 6809 26947 6824 26993
rect 6870 26947 6885 26993
rect 6809 26890 6885 26947
rect 6809 26844 6824 26890
rect 6870 26844 6885 26890
rect 6809 26787 6885 26844
rect 6809 26741 6824 26787
rect 6870 26741 6885 26787
rect 6809 26684 6885 26741
rect 6809 26638 6824 26684
rect 6870 26638 6885 26684
rect 6809 26581 6885 26638
rect 6809 26535 6824 26581
rect 6870 26535 6885 26581
rect 6809 26478 6885 26535
rect 6809 26432 6824 26478
rect 6870 26432 6885 26478
rect 6809 26375 6885 26432
rect 6809 26329 6824 26375
rect 6870 26329 6885 26375
rect 6809 26272 6885 26329
rect 6809 26226 6824 26272
rect 6870 26226 6885 26272
rect 6809 26169 6885 26226
rect 6809 26123 6824 26169
rect 6870 26123 6885 26169
rect 6809 26065 6885 26123
rect 6809 26019 6824 26065
rect 6870 26019 6885 26065
rect 2264 25780 6759 25791
rect 2264 25734 2275 25780
rect 6739 25734 6759 25780
rect 2264 25727 2276 25734
rect 3680 25727 4166 25734
rect 6090 25727 6759 25734
rect 2264 25723 6759 25727
rect 2264 25715 3692 25723
rect 4154 25715 6102 25723
rect 6809 25617 6885 26019
rect 7053 26993 7129 27006
rect 7053 26947 7068 26993
rect 7114 26947 7129 26993
rect 7053 26890 7129 26947
rect 7053 26844 7068 26890
rect 7114 26844 7129 26890
rect 7053 26787 7129 26844
rect 7053 26741 7068 26787
rect 7114 26741 7129 26787
rect 7053 26684 7129 26741
rect 7053 26638 7068 26684
rect 7114 26638 7129 26684
rect 7053 26581 7129 26638
rect 7053 26535 7068 26581
rect 7114 26535 7129 26581
rect 7053 26478 7129 26535
rect 7053 26432 7068 26478
rect 7114 26432 7129 26478
rect 7053 26375 7129 26432
rect 7053 26329 7068 26375
rect 7114 26329 7129 26375
rect 7053 26272 7129 26329
rect 7053 26226 7068 26272
rect 7114 26226 7129 26272
rect 7053 26169 7129 26226
rect 7053 26123 7068 26169
rect 7114 26123 7129 26169
rect 7053 26065 7129 26123
rect 7053 26019 7068 26065
rect 7114 26019 7129 26065
rect 7053 25791 7129 26019
rect 7297 26993 7373 27066
rect 7297 26947 7312 26993
rect 7358 26947 7373 26993
rect 7297 26890 7373 26947
rect 7297 26844 7312 26890
rect 7358 26844 7373 26890
rect 7297 26787 7373 26844
rect 7297 26741 7312 26787
rect 7358 26741 7373 26787
rect 7297 26684 7373 26741
rect 7297 26638 7312 26684
rect 7358 26638 7373 26684
rect 7297 26581 7373 26638
rect 7297 26535 7312 26581
rect 7358 26535 7373 26581
rect 7297 26478 7373 26535
rect 7297 26432 7312 26478
rect 7358 26432 7373 26478
rect 7297 26375 7373 26432
rect 7297 26329 7312 26375
rect 7358 26329 7373 26375
rect 7297 26272 7373 26329
rect 7297 26226 7312 26272
rect 7358 26226 7373 26272
rect 7297 26169 7373 26226
rect 7297 26123 7312 26169
rect 7358 26123 7373 26169
rect 7297 26065 7373 26123
rect 7297 26019 7312 26065
rect 7358 26019 7373 26065
rect 7297 25916 7373 26019
rect 7541 26993 7617 27006
rect 7541 26947 7556 26993
rect 7602 26947 7617 26993
rect 7541 26890 7617 26947
rect 7541 26844 7556 26890
rect 7602 26844 7617 26890
rect 7541 26787 7617 26844
rect 7541 26741 7556 26787
rect 7602 26741 7617 26787
rect 7541 26684 7617 26741
rect 7541 26638 7556 26684
rect 7602 26638 7617 26684
rect 7541 26581 7617 26638
rect 7541 26535 7556 26581
rect 7602 26535 7617 26581
rect 7541 26478 7617 26535
rect 7541 26432 7556 26478
rect 7602 26432 7617 26478
rect 7541 26375 7617 26432
rect 7541 26329 7556 26375
rect 7602 26329 7617 26375
rect 7541 26272 7617 26329
rect 7541 26226 7556 26272
rect 7602 26226 7617 26272
rect 7541 26169 7617 26226
rect 7541 26123 7556 26169
rect 7602 26123 7617 26169
rect 7541 26065 7617 26123
rect 7541 26019 7556 26065
rect 7602 26019 7617 26065
rect 7541 25791 7617 26019
rect 7785 26993 7861 27066
rect 7785 26947 7800 26993
rect 7846 26947 7861 26993
rect 7785 26890 7861 26947
rect 7785 26844 7800 26890
rect 7846 26844 7861 26890
rect 7785 26787 7861 26844
rect 7785 26741 7800 26787
rect 7846 26741 7861 26787
rect 7785 26684 7861 26741
rect 7785 26638 7800 26684
rect 7846 26638 7861 26684
rect 7785 26581 7861 26638
rect 7785 26535 7800 26581
rect 7846 26535 7861 26581
rect 7785 26478 7861 26535
rect 7785 26432 7800 26478
rect 7846 26432 7861 26478
rect 7785 26375 7861 26432
rect 7785 26329 7800 26375
rect 7846 26329 7861 26375
rect 7785 26272 7861 26329
rect 7785 26226 7800 26272
rect 7846 26226 7861 26272
rect 7785 26169 7861 26226
rect 7785 26123 7800 26169
rect 7846 26123 7861 26169
rect 7785 26065 7861 26123
rect 7785 26019 7800 26065
rect 7846 26019 7861 26065
rect 7785 25916 7861 26019
rect 8029 26993 8105 27006
rect 8029 26947 8044 26993
rect 8090 26947 8105 26993
rect 8029 26890 8105 26947
rect 8029 26844 8044 26890
rect 8090 26844 8105 26890
rect 8029 26787 8105 26844
rect 8029 26741 8044 26787
rect 8090 26741 8105 26787
rect 8029 26684 8105 26741
rect 8029 26638 8044 26684
rect 8090 26638 8105 26684
rect 8029 26581 8105 26638
rect 8029 26535 8044 26581
rect 8090 26535 8105 26581
rect 8029 26478 8105 26535
rect 8029 26432 8044 26478
rect 8090 26432 8105 26478
rect 8029 26375 8105 26432
rect 8029 26329 8044 26375
rect 8090 26329 8105 26375
rect 8029 26272 8105 26329
rect 8029 26226 8044 26272
rect 8090 26226 8105 26272
rect 8029 26169 8105 26226
rect 8029 26123 8044 26169
rect 8090 26123 8105 26169
rect 8029 26065 8105 26123
rect 8029 26019 8044 26065
rect 8090 26019 8105 26065
rect 8029 25791 8105 26019
rect 10622 25959 10634 27155
rect 10622 25947 10641 25959
rect 10630 25888 10641 25947
rect 10687 25888 10698 27156
rect 10630 25791 10698 25888
rect 6935 25780 10698 25791
rect 6935 25779 6975 25780
rect 7209 25779 7445 25780
rect 7679 25779 8009 25780
rect 6935 25727 6959 25779
rect 7219 25734 7445 25779
rect 7219 25727 7448 25734
rect 7708 25727 7963 25779
rect 10687 25734 10698 25780
rect 8847 25727 9282 25734
rect 10686 25727 10698 25734
rect 6935 25723 10698 25727
rect 6947 25715 7231 25723
rect 7436 25715 7720 25723
rect 7951 25715 8859 25723
rect 9270 25715 10698 25723
rect 1213 25597 11749 25617
rect 1213 25545 1233 25597
rect 1285 25545 1341 25597
rect 1393 25545 11569 25597
rect 11621 25545 11677 25597
rect 11729 25545 11749 25597
rect 1213 25489 11749 25545
rect 1213 25437 1233 25489
rect 1285 25437 1341 25489
rect 1393 25437 11569 25489
rect 11621 25437 11677 25489
rect 11729 25437 11749 25489
rect 1213 25417 11749 25437
<< via1 >>
rect 1493 45862 1545 45914
rect 1601 45862 1653 45914
rect 3863 45862 3915 45914
rect 3971 45862 4023 45914
rect 6239 45862 6291 45914
rect 6347 45862 6399 45914
rect 6455 45862 6507 45914
rect 6563 45862 6615 45914
rect 6671 45862 6723 45914
rect 8939 45862 8991 45914
rect 9047 45862 9099 45914
rect 11309 45862 11361 45914
rect 11417 45862 11469 45914
rect 1493 42122 1545 42174
rect 1601 42122 1653 42174
rect 3863 42122 3915 42174
rect 3971 42122 4023 42174
rect 6239 42122 6291 42174
rect 6347 42122 6399 42174
rect 6455 42122 6507 42174
rect 6563 42122 6615 42174
rect 6671 42122 6723 42174
rect 8939 42122 8991 42174
rect 9047 42122 9099 42174
rect 11309 42122 11361 42174
rect 11417 42122 11469 42174
rect 1760 41683 1812 41735
rect 1868 41683 1920 41735
rect 1976 41683 2028 41735
rect 2084 41683 2136 41735
rect 2192 41683 2244 41735
rect 2300 41683 2352 41735
rect 2408 41683 2460 41735
rect 2516 41683 2568 41735
rect 2624 41683 2676 41735
rect 2732 41683 2784 41735
rect 2840 41683 2892 41735
rect 2948 41683 3000 41735
rect 3056 41683 3108 41735
rect 3164 41683 3216 41735
rect 3272 41683 3324 41735
rect 3380 41683 3432 41735
rect 3488 41683 3540 41735
rect 3596 41683 3648 41735
rect 3704 41683 3756 41735
rect 1760 41575 1812 41627
rect 1868 41575 1920 41627
rect 1976 41575 2028 41627
rect 2084 41575 2136 41627
rect 2192 41575 2244 41627
rect 2300 41575 2352 41627
rect 2408 41575 2460 41627
rect 2516 41575 2568 41627
rect 2624 41575 2676 41627
rect 2732 41575 2784 41627
rect 2840 41575 2892 41627
rect 2948 41575 3000 41627
rect 3056 41575 3108 41627
rect 3164 41575 3216 41627
rect 3272 41575 3324 41627
rect 3380 41575 3432 41627
rect 3488 41575 3540 41627
rect 3596 41575 3648 41627
rect 3704 41575 3756 41627
rect 4130 41683 4182 41735
rect 4238 41683 4290 41735
rect 4346 41683 4398 41735
rect 4454 41683 4506 41735
rect 4562 41683 4614 41735
rect 4670 41683 4722 41735
rect 4778 41683 4830 41735
rect 4886 41683 4938 41735
rect 4994 41683 5046 41735
rect 5102 41683 5154 41735
rect 5210 41683 5262 41735
rect 5318 41683 5370 41735
rect 5426 41683 5478 41735
rect 5534 41683 5586 41735
rect 5642 41683 5694 41735
rect 5750 41683 5802 41735
rect 5858 41683 5910 41735
rect 5966 41683 6018 41735
rect 6074 41683 6126 41735
rect 4130 41575 4182 41627
rect 4238 41575 4290 41627
rect 4346 41575 4398 41627
rect 4454 41575 4506 41627
rect 4562 41575 4614 41627
rect 4670 41575 4722 41627
rect 4778 41575 4830 41627
rect 4886 41575 4938 41627
rect 4994 41575 5046 41627
rect 5102 41575 5154 41627
rect 5210 41575 5262 41627
rect 5318 41575 5370 41627
rect 5426 41575 5478 41627
rect 5534 41575 5586 41627
rect 5642 41575 5694 41627
rect 5750 41575 5802 41627
rect 5858 41575 5910 41627
rect 5966 41575 6018 41627
rect 6074 41575 6126 41627
rect 6836 41683 6888 41735
rect 6944 41683 6996 41735
rect 7052 41683 7104 41735
rect 7160 41683 7212 41735
rect 7268 41683 7320 41735
rect 7376 41683 7428 41735
rect 7484 41683 7536 41735
rect 7592 41683 7644 41735
rect 7700 41683 7752 41735
rect 7808 41683 7860 41735
rect 7916 41683 7968 41735
rect 8024 41683 8076 41735
rect 8132 41683 8184 41735
rect 8240 41683 8292 41735
rect 8348 41683 8400 41735
rect 8456 41683 8508 41735
rect 8564 41683 8616 41735
rect 8672 41683 8724 41735
rect 8780 41683 8832 41735
rect 6836 41575 6888 41627
rect 6944 41575 6996 41627
rect 7052 41575 7104 41627
rect 7160 41575 7212 41627
rect 7268 41575 7320 41627
rect 7376 41575 7428 41627
rect 7484 41575 7536 41627
rect 7592 41575 7644 41627
rect 7700 41575 7752 41627
rect 7808 41575 7860 41627
rect 7916 41575 7968 41627
rect 8024 41575 8076 41627
rect 8132 41575 8184 41627
rect 8240 41575 8292 41627
rect 8348 41575 8400 41627
rect 8456 41575 8508 41627
rect 8564 41575 8616 41627
rect 8672 41575 8724 41627
rect 8780 41575 8832 41627
rect 9206 41683 9258 41735
rect 9314 41683 9366 41735
rect 9422 41683 9474 41735
rect 9530 41683 9582 41735
rect 9638 41683 9690 41735
rect 9746 41683 9798 41735
rect 9854 41683 9906 41735
rect 9962 41683 10014 41735
rect 10070 41683 10122 41735
rect 10178 41683 10230 41735
rect 10286 41683 10338 41735
rect 10394 41683 10446 41735
rect 10502 41683 10554 41735
rect 10610 41683 10662 41735
rect 10718 41683 10770 41735
rect 10826 41683 10878 41735
rect 10934 41683 10986 41735
rect 11042 41683 11094 41735
rect 11150 41683 11202 41735
rect 9206 41575 9258 41627
rect 9314 41575 9366 41627
rect 9422 41575 9474 41627
rect 9530 41575 9582 41627
rect 9638 41575 9690 41627
rect 9746 41575 9798 41627
rect 9854 41575 9906 41627
rect 9962 41575 10014 41627
rect 10070 41575 10122 41627
rect 10178 41575 10230 41627
rect 10286 41575 10338 41627
rect 10394 41575 10446 41627
rect 10502 41575 10554 41627
rect 10610 41575 10662 41627
rect 10718 41575 10770 41627
rect 10826 41575 10878 41627
rect 10934 41575 10986 41627
rect 11042 41575 11094 41627
rect 11150 41575 11202 41627
rect 1802 35946 1854 35998
rect 1926 35946 1978 35998
rect 2050 35946 2102 35998
rect 2174 35946 2226 35998
rect 2298 35946 2350 35998
rect 2422 35946 2474 35998
rect 2546 35946 2598 35998
rect 2670 35946 2722 35998
rect 2794 35946 2846 35998
rect 2918 35946 2970 35998
rect 3042 35946 3094 35998
rect 3166 35946 3218 35998
rect 3290 35946 3342 35998
rect 3414 35946 3466 35998
rect 3538 35946 3590 35998
rect 3662 35946 3714 35998
rect 1802 35822 1854 35874
rect 1926 35822 1978 35874
rect 2050 35822 2102 35874
rect 2174 35822 2226 35874
rect 2298 35822 2350 35874
rect 2422 35822 2474 35874
rect 2546 35822 2598 35874
rect 2670 35822 2722 35874
rect 2794 35822 2846 35874
rect 2918 35822 2970 35874
rect 3042 35822 3094 35874
rect 3166 35822 3218 35874
rect 3290 35822 3342 35874
rect 3414 35822 3466 35874
rect 3538 35822 3590 35874
rect 3662 35822 3714 35874
rect 1802 35698 1854 35750
rect 1926 35698 1978 35750
rect 2050 35698 2102 35750
rect 2174 35698 2226 35750
rect 2298 35698 2350 35750
rect 2422 35698 2474 35750
rect 2546 35698 2598 35750
rect 2670 35698 2722 35750
rect 2794 35698 2846 35750
rect 2918 35698 2970 35750
rect 3042 35698 3094 35750
rect 3166 35698 3218 35750
rect 3290 35698 3342 35750
rect 3414 35698 3466 35750
rect 3538 35698 3590 35750
rect 3662 35698 3714 35750
rect 1802 35574 1854 35626
rect 1926 35574 1978 35626
rect 2050 35574 2102 35626
rect 2174 35574 2226 35626
rect 2298 35574 2350 35626
rect 2422 35574 2474 35626
rect 2546 35574 2598 35626
rect 2670 35574 2722 35626
rect 2794 35574 2846 35626
rect 2918 35574 2970 35626
rect 3042 35574 3094 35626
rect 3166 35574 3218 35626
rect 3290 35574 3342 35626
rect 3414 35574 3466 35626
rect 3538 35574 3590 35626
rect 3662 35574 3714 35626
rect 1802 35450 1854 35502
rect 1926 35450 1978 35502
rect 2050 35450 2102 35502
rect 2174 35450 2226 35502
rect 2298 35450 2350 35502
rect 2422 35450 2474 35502
rect 2546 35450 2598 35502
rect 2670 35450 2722 35502
rect 2794 35450 2846 35502
rect 2918 35450 2970 35502
rect 3042 35450 3094 35502
rect 3166 35450 3218 35502
rect 3290 35450 3342 35502
rect 3414 35450 3466 35502
rect 3538 35450 3590 35502
rect 3662 35450 3714 35502
rect 1802 35326 1854 35378
rect 1926 35326 1978 35378
rect 2050 35326 2102 35378
rect 2174 35326 2226 35378
rect 2298 35326 2350 35378
rect 2422 35326 2474 35378
rect 2546 35326 2598 35378
rect 2670 35326 2722 35378
rect 2794 35326 2846 35378
rect 2918 35326 2970 35378
rect 3042 35326 3094 35378
rect 3166 35326 3218 35378
rect 3290 35326 3342 35378
rect 3414 35326 3466 35378
rect 3538 35326 3590 35378
rect 3662 35326 3714 35378
rect 4172 35946 4224 35998
rect 4296 35946 4348 35998
rect 4420 35946 4472 35998
rect 4544 35946 4596 35998
rect 4668 35946 4720 35998
rect 4792 35946 4844 35998
rect 4916 35946 4968 35998
rect 5040 35946 5092 35998
rect 5164 35946 5216 35998
rect 5288 35946 5340 35998
rect 5412 35946 5464 35998
rect 5536 35946 5588 35998
rect 5660 35946 5712 35998
rect 5784 35946 5836 35998
rect 5908 35946 5960 35998
rect 6032 35946 6084 35998
rect 4172 35822 4224 35874
rect 4296 35822 4348 35874
rect 4420 35822 4472 35874
rect 4544 35822 4596 35874
rect 4668 35822 4720 35874
rect 4792 35822 4844 35874
rect 4916 35822 4968 35874
rect 5040 35822 5092 35874
rect 5164 35822 5216 35874
rect 5288 35822 5340 35874
rect 5412 35822 5464 35874
rect 5536 35822 5588 35874
rect 5660 35822 5712 35874
rect 5784 35822 5836 35874
rect 5908 35822 5960 35874
rect 6032 35822 6084 35874
rect 4172 35698 4224 35750
rect 4296 35698 4348 35750
rect 4420 35698 4472 35750
rect 4544 35698 4596 35750
rect 4668 35698 4720 35750
rect 4792 35698 4844 35750
rect 4916 35698 4968 35750
rect 5040 35698 5092 35750
rect 5164 35698 5216 35750
rect 5288 35698 5340 35750
rect 5412 35698 5464 35750
rect 5536 35698 5588 35750
rect 5660 35698 5712 35750
rect 5784 35698 5836 35750
rect 5908 35698 5960 35750
rect 6032 35698 6084 35750
rect 4172 35574 4224 35626
rect 4296 35574 4348 35626
rect 4420 35574 4472 35626
rect 4544 35574 4596 35626
rect 4668 35574 4720 35626
rect 4792 35574 4844 35626
rect 4916 35574 4968 35626
rect 5040 35574 5092 35626
rect 5164 35574 5216 35626
rect 5288 35574 5340 35626
rect 5412 35574 5464 35626
rect 5536 35574 5588 35626
rect 5660 35574 5712 35626
rect 5784 35574 5836 35626
rect 5908 35574 5960 35626
rect 6032 35574 6084 35626
rect 4172 35450 4224 35502
rect 4296 35450 4348 35502
rect 4420 35450 4472 35502
rect 4544 35450 4596 35502
rect 4668 35450 4720 35502
rect 4792 35450 4844 35502
rect 4916 35450 4968 35502
rect 5040 35450 5092 35502
rect 5164 35450 5216 35502
rect 5288 35450 5340 35502
rect 5412 35450 5464 35502
rect 5536 35450 5588 35502
rect 5660 35450 5712 35502
rect 5784 35450 5836 35502
rect 5908 35450 5960 35502
rect 6032 35450 6084 35502
rect 4172 35326 4224 35378
rect 4296 35326 4348 35378
rect 4420 35326 4472 35378
rect 4544 35326 4596 35378
rect 4668 35326 4720 35378
rect 4792 35326 4844 35378
rect 4916 35326 4968 35378
rect 5040 35326 5092 35378
rect 5164 35326 5216 35378
rect 5288 35326 5340 35378
rect 5412 35326 5464 35378
rect 5536 35326 5588 35378
rect 5660 35326 5712 35378
rect 5784 35326 5836 35378
rect 5908 35326 5960 35378
rect 6032 35326 6084 35378
rect 6878 35946 6930 35998
rect 7002 35946 7054 35998
rect 7126 35946 7178 35998
rect 7250 35946 7302 35998
rect 7374 35946 7426 35998
rect 7498 35946 7550 35998
rect 7622 35946 7674 35998
rect 7746 35946 7798 35998
rect 7870 35946 7922 35998
rect 7994 35946 8046 35998
rect 8118 35946 8170 35998
rect 8242 35946 8294 35998
rect 8366 35946 8418 35998
rect 8490 35946 8542 35998
rect 8614 35946 8666 35998
rect 8738 35946 8790 35998
rect 6878 35822 6930 35874
rect 7002 35822 7054 35874
rect 7126 35822 7178 35874
rect 7250 35822 7302 35874
rect 7374 35822 7426 35874
rect 7498 35822 7550 35874
rect 7622 35822 7674 35874
rect 7746 35822 7798 35874
rect 7870 35822 7922 35874
rect 7994 35822 8046 35874
rect 8118 35822 8170 35874
rect 8242 35822 8294 35874
rect 8366 35822 8418 35874
rect 8490 35822 8542 35874
rect 8614 35822 8666 35874
rect 8738 35822 8790 35874
rect 6878 35698 6930 35750
rect 7002 35698 7054 35750
rect 7126 35698 7178 35750
rect 7250 35698 7302 35750
rect 7374 35698 7426 35750
rect 7498 35698 7550 35750
rect 7622 35698 7674 35750
rect 7746 35698 7798 35750
rect 7870 35698 7922 35750
rect 7994 35698 8046 35750
rect 8118 35698 8170 35750
rect 8242 35698 8294 35750
rect 8366 35698 8418 35750
rect 8490 35698 8542 35750
rect 8614 35698 8666 35750
rect 8738 35698 8790 35750
rect 6878 35574 6930 35626
rect 7002 35574 7054 35626
rect 7126 35574 7178 35626
rect 7250 35574 7302 35626
rect 7374 35574 7426 35626
rect 7498 35574 7550 35626
rect 7622 35574 7674 35626
rect 7746 35574 7798 35626
rect 7870 35574 7922 35626
rect 7994 35574 8046 35626
rect 8118 35574 8170 35626
rect 8242 35574 8294 35626
rect 8366 35574 8418 35626
rect 8490 35574 8542 35626
rect 8614 35574 8666 35626
rect 8738 35574 8790 35626
rect 6878 35450 6930 35502
rect 7002 35450 7054 35502
rect 7126 35450 7178 35502
rect 7250 35450 7302 35502
rect 7374 35450 7426 35502
rect 7498 35450 7550 35502
rect 7622 35450 7674 35502
rect 7746 35450 7798 35502
rect 7870 35450 7922 35502
rect 7994 35450 8046 35502
rect 8118 35450 8170 35502
rect 8242 35450 8294 35502
rect 8366 35450 8418 35502
rect 8490 35450 8542 35502
rect 8614 35450 8666 35502
rect 8738 35450 8790 35502
rect 6878 35326 6930 35378
rect 7002 35326 7054 35378
rect 7126 35326 7178 35378
rect 7250 35326 7302 35378
rect 7374 35326 7426 35378
rect 7498 35326 7550 35378
rect 7622 35326 7674 35378
rect 7746 35326 7798 35378
rect 7870 35326 7922 35378
rect 7994 35326 8046 35378
rect 8118 35326 8170 35378
rect 8242 35326 8294 35378
rect 8366 35326 8418 35378
rect 8490 35326 8542 35378
rect 8614 35326 8666 35378
rect 8738 35326 8790 35378
rect 9248 35946 9300 35998
rect 9372 35946 9424 35998
rect 9496 35946 9548 35998
rect 9620 35946 9672 35998
rect 9744 35946 9796 35998
rect 9868 35946 9920 35998
rect 9992 35946 10044 35998
rect 10116 35946 10168 35998
rect 10240 35946 10292 35998
rect 10364 35946 10416 35998
rect 10488 35946 10540 35998
rect 10612 35946 10664 35998
rect 10736 35946 10788 35998
rect 10860 35946 10912 35998
rect 10984 35946 11036 35998
rect 11108 35946 11160 35998
rect 9248 35822 9300 35874
rect 9372 35822 9424 35874
rect 9496 35822 9548 35874
rect 9620 35822 9672 35874
rect 9744 35822 9796 35874
rect 9868 35822 9920 35874
rect 9992 35822 10044 35874
rect 10116 35822 10168 35874
rect 10240 35822 10292 35874
rect 10364 35822 10416 35874
rect 10488 35822 10540 35874
rect 10612 35822 10664 35874
rect 10736 35822 10788 35874
rect 10860 35822 10912 35874
rect 10984 35822 11036 35874
rect 11108 35822 11160 35874
rect 9248 35698 9300 35750
rect 9372 35698 9424 35750
rect 9496 35698 9548 35750
rect 9620 35698 9672 35750
rect 9744 35698 9796 35750
rect 9868 35698 9920 35750
rect 9992 35698 10044 35750
rect 10116 35698 10168 35750
rect 10240 35698 10292 35750
rect 10364 35698 10416 35750
rect 10488 35698 10540 35750
rect 10612 35698 10664 35750
rect 10736 35698 10788 35750
rect 10860 35698 10912 35750
rect 10984 35698 11036 35750
rect 11108 35698 11160 35750
rect 9248 35574 9300 35626
rect 9372 35574 9424 35626
rect 9496 35574 9548 35626
rect 9620 35574 9672 35626
rect 9744 35574 9796 35626
rect 9868 35574 9920 35626
rect 9992 35574 10044 35626
rect 10116 35574 10168 35626
rect 10240 35574 10292 35626
rect 10364 35574 10416 35626
rect 10488 35574 10540 35626
rect 10612 35574 10664 35626
rect 10736 35574 10788 35626
rect 10860 35574 10912 35626
rect 10984 35574 11036 35626
rect 11108 35574 11160 35626
rect 9248 35450 9300 35502
rect 9372 35450 9424 35502
rect 9496 35450 9548 35502
rect 9620 35450 9672 35502
rect 9744 35450 9796 35502
rect 9868 35450 9920 35502
rect 9992 35450 10044 35502
rect 10116 35450 10168 35502
rect 10240 35450 10292 35502
rect 10364 35450 10416 35502
rect 10488 35450 10540 35502
rect 10612 35450 10664 35502
rect 10736 35450 10788 35502
rect 10860 35450 10912 35502
rect 10984 35450 11036 35502
rect 11108 35450 11160 35502
rect 9248 35326 9300 35378
rect 9372 35326 9424 35378
rect 9496 35326 9548 35378
rect 9620 35326 9672 35378
rect 9744 35326 9796 35378
rect 9868 35326 9920 35378
rect 9992 35326 10044 35378
rect 10116 35326 10168 35378
rect 10240 35326 10292 35378
rect 10364 35326 10416 35378
rect 10488 35326 10540 35378
rect 10612 35326 10664 35378
rect 10736 35326 10788 35378
rect 10860 35326 10912 35378
rect 10984 35326 11036 35378
rect 11108 35326 11160 35378
rect 1760 29599 1812 29651
rect 1868 29599 1920 29651
rect 1976 29599 2028 29651
rect 2084 29599 2136 29651
rect 2192 29599 2244 29651
rect 2300 29599 2352 29651
rect 2408 29599 2460 29651
rect 2516 29599 2568 29651
rect 2624 29599 2676 29651
rect 2732 29599 2784 29651
rect 2840 29599 2892 29651
rect 2948 29599 3000 29651
rect 3056 29599 3108 29651
rect 3164 29599 3216 29651
rect 3272 29599 3324 29651
rect 3380 29599 3432 29651
rect 3488 29599 3540 29651
rect 3596 29599 3648 29651
rect 3704 29599 3756 29651
rect 1760 29491 1812 29543
rect 1868 29491 1920 29543
rect 1976 29491 2028 29543
rect 2084 29491 2136 29543
rect 2192 29491 2244 29543
rect 2300 29491 2352 29543
rect 2408 29491 2460 29543
rect 2516 29491 2568 29543
rect 2624 29491 2676 29543
rect 2732 29491 2784 29543
rect 2840 29491 2892 29543
rect 2948 29491 3000 29543
rect 3056 29491 3108 29543
rect 3164 29491 3216 29543
rect 3272 29491 3324 29543
rect 3380 29491 3432 29543
rect 3488 29491 3540 29543
rect 3596 29491 3648 29543
rect 3704 29491 3756 29543
rect 4130 29599 4182 29651
rect 4238 29599 4290 29651
rect 4346 29599 4398 29651
rect 4454 29599 4506 29651
rect 4562 29599 4614 29651
rect 4670 29599 4722 29651
rect 4778 29599 4830 29651
rect 4886 29599 4938 29651
rect 4994 29599 5046 29651
rect 5102 29599 5154 29651
rect 5210 29599 5262 29651
rect 5318 29599 5370 29651
rect 5426 29599 5478 29651
rect 5534 29599 5586 29651
rect 5642 29599 5694 29651
rect 5750 29599 5802 29651
rect 5858 29599 5910 29651
rect 5966 29599 6018 29651
rect 6074 29599 6126 29651
rect 4130 29491 4182 29543
rect 4238 29491 4290 29543
rect 4346 29491 4398 29543
rect 4454 29491 4506 29543
rect 4562 29491 4614 29543
rect 4670 29491 4722 29543
rect 4778 29491 4830 29543
rect 4886 29491 4938 29543
rect 4994 29491 5046 29543
rect 5102 29491 5154 29543
rect 5210 29491 5262 29543
rect 5318 29491 5370 29543
rect 5426 29491 5478 29543
rect 5534 29491 5586 29543
rect 5642 29491 5694 29543
rect 5750 29491 5802 29543
rect 5858 29491 5910 29543
rect 5966 29491 6018 29543
rect 6074 29491 6126 29543
rect 6836 29599 6888 29651
rect 6944 29599 6996 29651
rect 7052 29599 7104 29651
rect 7160 29599 7212 29651
rect 7268 29599 7320 29651
rect 7376 29599 7428 29651
rect 7484 29599 7536 29651
rect 7592 29599 7644 29651
rect 7700 29599 7752 29651
rect 7808 29599 7860 29651
rect 7916 29599 7968 29651
rect 8024 29599 8076 29651
rect 8132 29599 8184 29651
rect 8240 29599 8292 29651
rect 8348 29599 8400 29651
rect 8456 29599 8508 29651
rect 8564 29599 8616 29651
rect 8672 29599 8724 29651
rect 8780 29599 8832 29651
rect 6836 29491 6888 29543
rect 6944 29491 6996 29543
rect 7052 29491 7104 29543
rect 7160 29491 7212 29543
rect 7268 29491 7320 29543
rect 7376 29491 7428 29543
rect 7484 29491 7536 29543
rect 7592 29491 7644 29543
rect 7700 29491 7752 29543
rect 7808 29491 7860 29543
rect 7916 29491 7968 29543
rect 8024 29491 8076 29543
rect 8132 29491 8184 29543
rect 8240 29491 8292 29543
rect 8348 29491 8400 29543
rect 8456 29491 8508 29543
rect 8564 29491 8616 29543
rect 8672 29491 8724 29543
rect 8780 29491 8832 29543
rect 9206 29599 9258 29651
rect 9314 29599 9366 29651
rect 9422 29599 9474 29651
rect 9530 29599 9582 29651
rect 9638 29599 9690 29651
rect 9746 29599 9798 29651
rect 9854 29599 9906 29651
rect 9962 29599 10014 29651
rect 10070 29599 10122 29651
rect 10178 29599 10230 29651
rect 10286 29599 10338 29651
rect 10394 29599 10446 29651
rect 10502 29599 10554 29651
rect 10610 29599 10662 29651
rect 10718 29599 10770 29651
rect 10826 29599 10878 29651
rect 10934 29599 10986 29651
rect 11042 29599 11094 29651
rect 11150 29599 11202 29651
rect 9206 29491 9258 29543
rect 9314 29491 9366 29543
rect 9422 29491 9474 29543
rect 9530 29491 9582 29543
rect 9638 29491 9690 29543
rect 9746 29491 9798 29543
rect 9854 29491 9906 29543
rect 9962 29491 10014 29543
rect 10070 29491 10122 29543
rect 10178 29491 10230 29543
rect 10286 29491 10338 29543
rect 10394 29491 10446 29543
rect 10502 29491 10554 29543
rect 10610 29491 10662 29543
rect 10718 29491 10770 29543
rect 10826 29491 10878 29543
rect 10934 29491 10986 29543
rect 11042 29491 11094 29543
rect 11150 29491 11202 29543
rect 1495 29135 1651 29187
rect 3865 29142 4021 29187
rect 6247 29142 6715 29187
rect 8941 29142 9097 29187
rect 3865 29135 4021 29142
rect 6247 29135 6715 29142
rect 8941 29135 9097 29142
rect 11311 29135 11467 29187
rect 2276 25959 2321 27155
rect 2321 25959 2328 27155
rect 4166 27439 6090 27484
rect 4166 27432 6090 27439
rect 6872 27439 6889 27484
rect 6889 27439 8796 27484
rect 9236 27439 10224 27484
rect 6872 27432 8796 27439
rect 9236 27432 10224 27439
rect 2276 25734 3680 25779
rect 4166 25734 6090 25779
rect 2276 25727 3680 25734
rect 4166 25727 6090 25734
rect 10634 25959 10641 27155
rect 10641 25959 10686 27155
rect 6959 25734 6975 25779
rect 6975 25734 7209 25779
rect 7209 25734 7219 25779
rect 7448 25734 7679 25779
rect 7679 25734 7708 25779
rect 6959 25727 7219 25734
rect 7448 25727 7708 25734
rect 7963 25734 8009 25779
rect 8009 25734 8847 25779
rect 9282 25734 10686 25779
rect 7963 25727 8847 25734
rect 9282 25727 10686 25734
rect 1233 25545 1285 25597
rect 1341 25545 1393 25597
rect 11569 25545 11621 25597
rect 11677 25545 11729 25597
rect 1233 25437 1285 25489
rect 1341 25437 1393 25489
rect 11569 25437 11621 25489
rect 11677 25437 11729 25489
<< metal2 >>
rect -747 25617 1153 46134
rect 1473 45914 1673 46134
rect 1473 45862 1493 45914
rect 1545 45862 1601 45914
rect 1653 45862 1673 45914
rect 1473 42174 1673 45862
rect 1473 42122 1493 42174
rect 1545 42122 1601 42174
rect 1653 42122 1673 42174
rect 1473 29187 1673 42122
rect 1473 29135 1495 29187
rect 1651 29135 1673 29187
rect 1473 25617 1673 29135
rect 1733 41735 3783 46134
rect 1733 41683 1760 41735
rect 1812 41683 1868 41735
rect 1920 41683 1976 41735
rect 2028 41683 2084 41735
rect 2136 41683 2192 41735
rect 2244 41683 2300 41735
rect 2352 41683 2408 41735
rect 2460 41683 2516 41735
rect 2568 41683 2624 41735
rect 2676 41683 2732 41735
rect 2784 41683 2840 41735
rect 2892 41683 2948 41735
rect 3000 41683 3056 41735
rect 3108 41683 3164 41735
rect 3216 41683 3272 41735
rect 3324 41683 3380 41735
rect 3432 41683 3488 41735
rect 3540 41683 3596 41735
rect 3648 41683 3704 41735
rect 3756 41683 3783 41735
rect 1733 41627 3783 41683
rect 1733 41575 1760 41627
rect 1812 41575 1868 41627
rect 1920 41575 1976 41627
rect 2028 41575 2084 41627
rect 2136 41575 2192 41627
rect 2244 41575 2300 41627
rect 2352 41575 2408 41627
rect 2460 41575 2516 41627
rect 2568 41575 2624 41627
rect 2676 41575 2732 41627
rect 2784 41575 2840 41627
rect 2892 41575 2948 41627
rect 3000 41575 3056 41627
rect 3108 41575 3164 41627
rect 3216 41575 3272 41627
rect 3324 41575 3380 41627
rect 3432 41575 3488 41627
rect 3540 41575 3596 41627
rect 3648 41575 3704 41627
rect 3756 41575 3783 41627
rect 1733 35998 3783 41575
rect 1733 35946 1802 35998
rect 1854 35946 1926 35998
rect 1978 35946 2050 35998
rect 2102 35946 2174 35998
rect 2226 35946 2298 35998
rect 2350 35946 2422 35998
rect 2474 35946 2546 35998
rect 2598 35946 2670 35998
rect 2722 35946 2794 35998
rect 2846 35946 2918 35998
rect 2970 35946 3042 35998
rect 3094 35946 3166 35998
rect 3218 35946 3290 35998
rect 3342 35946 3414 35998
rect 3466 35946 3538 35998
rect 3590 35946 3662 35998
rect 3714 35946 3783 35998
rect 1733 35874 3783 35946
rect 1733 35822 1802 35874
rect 1854 35822 1926 35874
rect 1978 35822 2050 35874
rect 2102 35822 2174 35874
rect 2226 35822 2298 35874
rect 2350 35822 2422 35874
rect 2474 35822 2546 35874
rect 2598 35822 2670 35874
rect 2722 35822 2794 35874
rect 2846 35822 2918 35874
rect 2970 35822 3042 35874
rect 3094 35822 3166 35874
rect 3218 35822 3290 35874
rect 3342 35822 3414 35874
rect 3466 35822 3538 35874
rect 3590 35822 3662 35874
rect 3714 35822 3783 35874
rect 1733 35750 3783 35822
rect 1733 35698 1802 35750
rect 1854 35698 1926 35750
rect 1978 35698 2050 35750
rect 2102 35698 2174 35750
rect 2226 35698 2298 35750
rect 2350 35698 2422 35750
rect 2474 35698 2546 35750
rect 2598 35698 2670 35750
rect 2722 35698 2794 35750
rect 2846 35698 2918 35750
rect 2970 35698 3042 35750
rect 3094 35698 3166 35750
rect 3218 35698 3290 35750
rect 3342 35698 3414 35750
rect 3466 35698 3538 35750
rect 3590 35698 3662 35750
rect 3714 35698 3783 35750
rect 1733 35626 3783 35698
rect 1733 35574 1802 35626
rect 1854 35574 1926 35626
rect 1978 35574 2050 35626
rect 2102 35574 2174 35626
rect 2226 35574 2298 35626
rect 2350 35574 2422 35626
rect 2474 35574 2546 35626
rect 2598 35574 2670 35626
rect 2722 35574 2794 35626
rect 2846 35574 2918 35626
rect 2970 35574 3042 35626
rect 3094 35574 3166 35626
rect 3218 35574 3290 35626
rect 3342 35574 3414 35626
rect 3466 35574 3538 35626
rect 3590 35574 3662 35626
rect 3714 35574 3783 35626
rect 1733 35502 3783 35574
rect 1733 35450 1802 35502
rect 1854 35450 1926 35502
rect 1978 35450 2050 35502
rect 2102 35450 2174 35502
rect 2226 35450 2298 35502
rect 2350 35450 2422 35502
rect 2474 35450 2546 35502
rect 2598 35450 2670 35502
rect 2722 35450 2794 35502
rect 2846 35450 2918 35502
rect 2970 35450 3042 35502
rect 3094 35450 3166 35502
rect 3218 35450 3290 35502
rect 3342 35450 3414 35502
rect 3466 35450 3538 35502
rect 3590 35450 3662 35502
rect 3714 35450 3783 35502
rect 1733 35378 3783 35450
rect 1733 35326 1802 35378
rect 1854 35326 1926 35378
rect 1978 35326 2050 35378
rect 2102 35326 2174 35378
rect 2226 35326 2298 35378
rect 2350 35326 2422 35378
rect 2474 35326 2546 35378
rect 2598 35326 2670 35378
rect 2722 35326 2794 35378
rect 2846 35326 2918 35378
rect 2970 35326 3042 35378
rect 3094 35326 3166 35378
rect 3218 35326 3290 35378
rect 3342 35326 3414 35378
rect 3466 35326 3538 35378
rect 3590 35326 3662 35378
rect 3714 35326 3783 35378
rect 1733 29651 3783 35326
rect 1733 29599 1760 29651
rect 1812 29599 1868 29651
rect 1920 29599 1976 29651
rect 2028 29599 2084 29651
rect 2136 29599 2192 29651
rect 2244 29599 2300 29651
rect 2352 29599 2408 29651
rect 2460 29599 2516 29651
rect 2568 29599 2624 29651
rect 2676 29599 2732 29651
rect 2784 29599 2840 29651
rect 2892 29599 2948 29651
rect 3000 29599 3056 29651
rect 3108 29599 3164 29651
rect 3216 29599 3272 29651
rect 3324 29599 3380 29651
rect 3432 29599 3488 29651
rect 3540 29599 3596 29651
rect 3648 29599 3704 29651
rect 3756 29599 3783 29651
rect 1733 29543 3783 29599
rect 1733 29491 1760 29543
rect 1812 29491 1868 29543
rect 1920 29491 1976 29543
rect 2028 29491 2084 29543
rect 2136 29491 2192 29543
rect 2244 29491 2300 29543
rect 2352 29491 2408 29543
rect 2460 29491 2516 29543
rect 2568 29491 2624 29543
rect 2676 29491 2732 29543
rect 2784 29491 2840 29543
rect 2892 29491 2948 29543
rect 3000 29491 3056 29543
rect 3108 29491 3164 29543
rect 3216 29491 3272 29543
rect 3324 29491 3380 29543
rect 3432 29491 3488 29543
rect 3540 29491 3596 29543
rect 3648 29491 3704 29543
rect 3756 29491 3783 29543
rect 1733 27155 3783 29491
rect 1733 25959 2276 27155
rect 2328 25959 3783 27155
rect 1733 25779 3783 25959
rect 1733 25727 2276 25779
rect 3680 25727 3783 25779
rect 1733 25617 3783 25727
rect 3843 45914 4043 46134
rect 3843 45862 3863 45914
rect 3915 45862 3971 45914
rect 4023 45862 4043 45914
rect 3843 42174 4043 45862
rect 3843 42122 3863 42174
rect 3915 42122 3971 42174
rect 4023 42122 4043 42174
rect 3843 29187 4043 42122
rect 3843 29135 3865 29187
rect 4021 29135 4043 29187
rect 3843 25617 4043 29135
rect 4103 41735 6153 46134
rect 4103 41683 4130 41735
rect 4182 41683 4238 41735
rect 4290 41683 4346 41735
rect 4398 41683 4454 41735
rect 4506 41683 4562 41735
rect 4614 41683 4670 41735
rect 4722 41683 4778 41735
rect 4830 41683 4886 41735
rect 4938 41683 4994 41735
rect 5046 41683 5102 41735
rect 5154 41683 5210 41735
rect 5262 41683 5318 41735
rect 5370 41683 5426 41735
rect 5478 41683 5534 41735
rect 5586 41683 5642 41735
rect 5694 41683 5750 41735
rect 5802 41683 5858 41735
rect 5910 41683 5966 41735
rect 6018 41683 6074 41735
rect 6126 41683 6153 41735
rect 4103 41627 6153 41683
rect 4103 41575 4130 41627
rect 4182 41575 4238 41627
rect 4290 41575 4346 41627
rect 4398 41575 4454 41627
rect 4506 41575 4562 41627
rect 4614 41575 4670 41627
rect 4722 41575 4778 41627
rect 4830 41575 4886 41627
rect 4938 41575 4994 41627
rect 5046 41575 5102 41627
rect 5154 41575 5210 41627
rect 5262 41575 5318 41627
rect 5370 41575 5426 41627
rect 5478 41575 5534 41627
rect 5586 41575 5642 41627
rect 5694 41575 5750 41627
rect 5802 41575 5858 41627
rect 5910 41575 5966 41627
rect 6018 41575 6074 41627
rect 6126 41575 6153 41627
rect 4103 35998 6153 41575
rect 4103 35946 4172 35998
rect 4224 35946 4296 35998
rect 4348 35946 4420 35998
rect 4472 35946 4544 35998
rect 4596 35946 4668 35998
rect 4720 35946 4792 35998
rect 4844 35946 4916 35998
rect 4968 35946 5040 35998
rect 5092 35946 5164 35998
rect 5216 35946 5288 35998
rect 5340 35946 5412 35998
rect 5464 35946 5536 35998
rect 5588 35946 5660 35998
rect 5712 35946 5784 35998
rect 5836 35946 5908 35998
rect 5960 35946 6032 35998
rect 6084 35946 6153 35998
rect 4103 35874 6153 35946
rect 4103 35822 4172 35874
rect 4224 35822 4296 35874
rect 4348 35822 4420 35874
rect 4472 35822 4544 35874
rect 4596 35822 4668 35874
rect 4720 35822 4792 35874
rect 4844 35822 4916 35874
rect 4968 35822 5040 35874
rect 5092 35822 5164 35874
rect 5216 35822 5288 35874
rect 5340 35822 5412 35874
rect 5464 35822 5536 35874
rect 5588 35822 5660 35874
rect 5712 35822 5784 35874
rect 5836 35822 5908 35874
rect 5960 35822 6032 35874
rect 6084 35822 6153 35874
rect 4103 35750 6153 35822
rect 4103 35698 4172 35750
rect 4224 35698 4296 35750
rect 4348 35698 4420 35750
rect 4472 35698 4544 35750
rect 4596 35698 4668 35750
rect 4720 35698 4792 35750
rect 4844 35698 4916 35750
rect 4968 35698 5040 35750
rect 5092 35698 5164 35750
rect 5216 35698 5288 35750
rect 5340 35698 5412 35750
rect 5464 35698 5536 35750
rect 5588 35698 5660 35750
rect 5712 35698 5784 35750
rect 5836 35698 5908 35750
rect 5960 35698 6032 35750
rect 6084 35698 6153 35750
rect 4103 35626 6153 35698
rect 4103 35574 4172 35626
rect 4224 35574 4296 35626
rect 4348 35574 4420 35626
rect 4472 35574 4544 35626
rect 4596 35574 4668 35626
rect 4720 35574 4792 35626
rect 4844 35574 4916 35626
rect 4968 35574 5040 35626
rect 5092 35574 5164 35626
rect 5216 35574 5288 35626
rect 5340 35574 5412 35626
rect 5464 35574 5536 35626
rect 5588 35574 5660 35626
rect 5712 35574 5784 35626
rect 5836 35574 5908 35626
rect 5960 35574 6032 35626
rect 6084 35574 6153 35626
rect 4103 35502 6153 35574
rect 4103 35450 4172 35502
rect 4224 35450 4296 35502
rect 4348 35450 4420 35502
rect 4472 35450 4544 35502
rect 4596 35450 4668 35502
rect 4720 35450 4792 35502
rect 4844 35450 4916 35502
rect 4968 35450 5040 35502
rect 5092 35450 5164 35502
rect 5216 35450 5288 35502
rect 5340 35450 5412 35502
rect 5464 35450 5536 35502
rect 5588 35450 5660 35502
rect 5712 35450 5784 35502
rect 5836 35450 5908 35502
rect 5960 35450 6032 35502
rect 6084 35450 6153 35502
rect 4103 35378 6153 35450
rect 4103 35326 4172 35378
rect 4224 35326 4296 35378
rect 4348 35326 4420 35378
rect 4472 35326 4544 35378
rect 4596 35326 4668 35378
rect 4720 35326 4792 35378
rect 4844 35326 4916 35378
rect 4968 35326 5040 35378
rect 5092 35326 5164 35378
rect 5216 35326 5288 35378
rect 5340 35326 5412 35378
rect 5464 35326 5536 35378
rect 5588 35326 5660 35378
rect 5712 35326 5784 35378
rect 5836 35326 5908 35378
rect 5960 35326 6032 35378
rect 6084 35326 6153 35378
rect 4103 29651 6153 35326
rect 4103 29599 4130 29651
rect 4182 29599 4238 29651
rect 4290 29599 4346 29651
rect 4398 29599 4454 29651
rect 4506 29599 4562 29651
rect 4614 29599 4670 29651
rect 4722 29599 4778 29651
rect 4830 29599 4886 29651
rect 4938 29599 4994 29651
rect 5046 29599 5102 29651
rect 5154 29599 5210 29651
rect 5262 29599 5318 29651
rect 5370 29599 5426 29651
rect 5478 29599 5534 29651
rect 5586 29599 5642 29651
rect 5694 29599 5750 29651
rect 5802 29599 5858 29651
rect 5910 29599 5966 29651
rect 6018 29599 6074 29651
rect 6126 29599 6153 29651
rect 4103 29543 6153 29599
rect 4103 29491 4130 29543
rect 4182 29491 4238 29543
rect 4290 29491 4346 29543
rect 4398 29491 4454 29543
rect 4506 29491 4562 29543
rect 4614 29491 4670 29543
rect 4722 29491 4778 29543
rect 4830 29491 4886 29543
rect 4938 29491 4994 29543
rect 5046 29491 5102 29543
rect 5154 29491 5210 29543
rect 5262 29491 5318 29543
rect 5370 29491 5426 29543
rect 5478 29491 5534 29543
rect 5586 29491 5642 29543
rect 5694 29491 5750 29543
rect 5802 29491 5858 29543
rect 5910 29491 5966 29543
rect 6018 29491 6074 29543
rect 6126 29491 6153 29543
rect 4103 27484 6153 29491
rect 4103 27432 4166 27484
rect 6090 27432 6153 27484
rect 4103 25779 6153 27432
rect 4103 25727 4166 25779
rect 6090 25727 6153 25779
rect 4103 25617 6153 25727
rect 6213 45914 6749 46134
rect 6213 45862 6239 45914
rect 6291 45862 6347 45914
rect 6399 45862 6455 45914
rect 6507 45862 6563 45914
rect 6615 45862 6671 45914
rect 6723 45862 6749 45914
rect 6213 42174 6749 45862
rect 6213 42122 6239 42174
rect 6291 42122 6347 42174
rect 6399 42122 6455 42174
rect 6507 42122 6563 42174
rect 6615 42122 6671 42174
rect 6723 42122 6749 42174
rect 6213 29187 6749 42122
rect 6213 29135 6247 29187
rect 6715 29135 6749 29187
rect 6213 25617 6749 29135
rect 6809 41735 8859 46134
rect 6809 41683 6836 41735
rect 6888 41683 6944 41735
rect 6996 41683 7052 41735
rect 7104 41683 7160 41735
rect 7212 41683 7268 41735
rect 7320 41683 7376 41735
rect 7428 41683 7484 41735
rect 7536 41683 7592 41735
rect 7644 41683 7700 41735
rect 7752 41683 7808 41735
rect 7860 41683 7916 41735
rect 7968 41683 8024 41735
rect 8076 41683 8132 41735
rect 8184 41683 8240 41735
rect 8292 41683 8348 41735
rect 8400 41683 8456 41735
rect 8508 41683 8564 41735
rect 8616 41683 8672 41735
rect 8724 41683 8780 41735
rect 8832 41683 8859 41735
rect 6809 41627 8859 41683
rect 6809 41575 6836 41627
rect 6888 41575 6944 41627
rect 6996 41575 7052 41627
rect 7104 41575 7160 41627
rect 7212 41575 7268 41627
rect 7320 41575 7376 41627
rect 7428 41575 7484 41627
rect 7536 41575 7592 41627
rect 7644 41575 7700 41627
rect 7752 41575 7808 41627
rect 7860 41575 7916 41627
rect 7968 41575 8024 41627
rect 8076 41575 8132 41627
rect 8184 41575 8240 41627
rect 8292 41575 8348 41627
rect 8400 41575 8456 41627
rect 8508 41575 8564 41627
rect 8616 41575 8672 41627
rect 8724 41575 8780 41627
rect 8832 41575 8859 41627
rect 6809 35998 8859 41575
rect 6809 35946 6878 35998
rect 6930 35946 7002 35998
rect 7054 35946 7126 35998
rect 7178 35946 7250 35998
rect 7302 35946 7374 35998
rect 7426 35946 7498 35998
rect 7550 35946 7622 35998
rect 7674 35946 7746 35998
rect 7798 35946 7870 35998
rect 7922 35946 7994 35998
rect 8046 35946 8118 35998
rect 8170 35946 8242 35998
rect 8294 35946 8366 35998
rect 8418 35946 8490 35998
rect 8542 35946 8614 35998
rect 8666 35946 8738 35998
rect 8790 35946 8859 35998
rect 6809 35874 8859 35946
rect 6809 35822 6878 35874
rect 6930 35822 7002 35874
rect 7054 35822 7126 35874
rect 7178 35822 7250 35874
rect 7302 35822 7374 35874
rect 7426 35822 7498 35874
rect 7550 35822 7622 35874
rect 7674 35822 7746 35874
rect 7798 35822 7870 35874
rect 7922 35822 7994 35874
rect 8046 35822 8118 35874
rect 8170 35822 8242 35874
rect 8294 35822 8366 35874
rect 8418 35822 8490 35874
rect 8542 35822 8614 35874
rect 8666 35822 8738 35874
rect 8790 35822 8859 35874
rect 6809 35750 8859 35822
rect 6809 35698 6878 35750
rect 6930 35698 7002 35750
rect 7054 35698 7126 35750
rect 7178 35698 7250 35750
rect 7302 35698 7374 35750
rect 7426 35698 7498 35750
rect 7550 35698 7622 35750
rect 7674 35698 7746 35750
rect 7798 35698 7870 35750
rect 7922 35698 7994 35750
rect 8046 35698 8118 35750
rect 8170 35698 8242 35750
rect 8294 35698 8366 35750
rect 8418 35698 8490 35750
rect 8542 35698 8614 35750
rect 8666 35698 8738 35750
rect 8790 35698 8859 35750
rect 6809 35626 8859 35698
rect 6809 35574 6878 35626
rect 6930 35574 7002 35626
rect 7054 35574 7126 35626
rect 7178 35574 7250 35626
rect 7302 35574 7374 35626
rect 7426 35574 7498 35626
rect 7550 35574 7622 35626
rect 7674 35574 7746 35626
rect 7798 35574 7870 35626
rect 7922 35574 7994 35626
rect 8046 35574 8118 35626
rect 8170 35574 8242 35626
rect 8294 35574 8366 35626
rect 8418 35574 8490 35626
rect 8542 35574 8614 35626
rect 8666 35574 8738 35626
rect 8790 35574 8859 35626
rect 6809 35502 8859 35574
rect 6809 35450 6878 35502
rect 6930 35450 7002 35502
rect 7054 35450 7126 35502
rect 7178 35450 7250 35502
rect 7302 35450 7374 35502
rect 7426 35450 7498 35502
rect 7550 35450 7622 35502
rect 7674 35450 7746 35502
rect 7798 35450 7870 35502
rect 7922 35450 7994 35502
rect 8046 35450 8118 35502
rect 8170 35450 8242 35502
rect 8294 35450 8366 35502
rect 8418 35450 8490 35502
rect 8542 35450 8614 35502
rect 8666 35450 8738 35502
rect 8790 35450 8859 35502
rect 6809 35378 8859 35450
rect 6809 35326 6878 35378
rect 6930 35326 7002 35378
rect 7054 35326 7126 35378
rect 7178 35326 7250 35378
rect 7302 35326 7374 35378
rect 7426 35326 7498 35378
rect 7550 35326 7622 35378
rect 7674 35326 7746 35378
rect 7798 35326 7870 35378
rect 7922 35326 7994 35378
rect 8046 35326 8118 35378
rect 8170 35326 8242 35378
rect 8294 35326 8366 35378
rect 8418 35326 8490 35378
rect 8542 35326 8614 35378
rect 8666 35326 8738 35378
rect 8790 35326 8859 35378
rect 6809 29651 8859 35326
rect 6809 29599 6836 29651
rect 6888 29599 6944 29651
rect 6996 29599 7052 29651
rect 7104 29599 7160 29651
rect 7212 29599 7268 29651
rect 7320 29599 7376 29651
rect 7428 29599 7484 29651
rect 7536 29599 7592 29651
rect 7644 29599 7700 29651
rect 7752 29599 7808 29651
rect 7860 29599 7916 29651
rect 7968 29599 8024 29651
rect 8076 29599 8132 29651
rect 8184 29599 8240 29651
rect 8292 29599 8348 29651
rect 8400 29599 8456 29651
rect 8508 29599 8564 29651
rect 8616 29599 8672 29651
rect 8724 29599 8780 29651
rect 8832 29599 8859 29651
rect 6809 29543 8859 29599
rect 6809 29491 6836 29543
rect 6888 29491 6944 29543
rect 6996 29491 7052 29543
rect 7104 29491 7160 29543
rect 7212 29491 7268 29543
rect 7320 29491 7376 29543
rect 7428 29491 7484 29543
rect 7536 29491 7592 29543
rect 7644 29491 7700 29543
rect 7752 29491 7808 29543
rect 7860 29491 7916 29543
rect 7968 29491 8024 29543
rect 8076 29491 8132 29543
rect 8184 29491 8240 29543
rect 8292 29491 8348 29543
rect 8400 29491 8456 29543
rect 8508 29491 8564 29543
rect 8616 29491 8672 29543
rect 8724 29491 8780 29543
rect 8832 29491 8859 29543
rect 6809 27484 8859 29491
rect 6809 27432 6872 27484
rect 8796 27432 8859 27484
rect 6809 25779 8859 27432
rect 6809 25727 6959 25779
rect 7219 25727 7448 25779
rect 7708 25727 7963 25779
rect 8847 25727 8859 25779
rect 6809 25617 8859 25727
rect 8919 45914 9119 46134
rect 8919 45862 8939 45914
rect 8991 45862 9047 45914
rect 9099 45862 9119 45914
rect 8919 42174 9119 45862
rect 8919 42122 8939 42174
rect 8991 42122 9047 42174
rect 9099 42122 9119 42174
rect 8919 29187 9119 42122
rect 8919 29135 8941 29187
rect 9097 29135 9119 29187
rect 8919 25617 9119 29135
rect 9179 41735 11229 46134
rect 9179 41683 9206 41735
rect 9258 41683 9314 41735
rect 9366 41683 9422 41735
rect 9474 41683 9530 41735
rect 9582 41683 9638 41735
rect 9690 41683 9746 41735
rect 9798 41683 9854 41735
rect 9906 41683 9962 41735
rect 10014 41683 10070 41735
rect 10122 41683 10178 41735
rect 10230 41683 10286 41735
rect 10338 41683 10394 41735
rect 10446 41683 10502 41735
rect 10554 41683 10610 41735
rect 10662 41683 10718 41735
rect 10770 41683 10826 41735
rect 10878 41683 10934 41735
rect 10986 41683 11042 41735
rect 11094 41683 11150 41735
rect 11202 41683 11229 41735
rect 9179 41627 11229 41683
rect 9179 41575 9206 41627
rect 9258 41575 9314 41627
rect 9366 41575 9422 41627
rect 9474 41575 9530 41627
rect 9582 41575 9638 41627
rect 9690 41575 9746 41627
rect 9798 41575 9854 41627
rect 9906 41575 9962 41627
rect 10014 41575 10070 41627
rect 10122 41575 10178 41627
rect 10230 41575 10286 41627
rect 10338 41575 10394 41627
rect 10446 41575 10502 41627
rect 10554 41575 10610 41627
rect 10662 41575 10718 41627
rect 10770 41575 10826 41627
rect 10878 41575 10934 41627
rect 10986 41575 11042 41627
rect 11094 41575 11150 41627
rect 11202 41575 11229 41627
rect 9179 35998 11229 41575
rect 9179 35946 9248 35998
rect 9300 35946 9372 35998
rect 9424 35946 9496 35998
rect 9548 35946 9620 35998
rect 9672 35946 9744 35998
rect 9796 35946 9868 35998
rect 9920 35946 9992 35998
rect 10044 35946 10116 35998
rect 10168 35946 10240 35998
rect 10292 35946 10364 35998
rect 10416 35946 10488 35998
rect 10540 35946 10612 35998
rect 10664 35946 10736 35998
rect 10788 35946 10860 35998
rect 10912 35946 10984 35998
rect 11036 35946 11108 35998
rect 11160 35946 11229 35998
rect 9179 35874 11229 35946
rect 9179 35822 9248 35874
rect 9300 35822 9372 35874
rect 9424 35822 9496 35874
rect 9548 35822 9620 35874
rect 9672 35822 9744 35874
rect 9796 35822 9868 35874
rect 9920 35822 9992 35874
rect 10044 35822 10116 35874
rect 10168 35822 10240 35874
rect 10292 35822 10364 35874
rect 10416 35822 10488 35874
rect 10540 35822 10612 35874
rect 10664 35822 10736 35874
rect 10788 35822 10860 35874
rect 10912 35822 10984 35874
rect 11036 35822 11108 35874
rect 11160 35822 11229 35874
rect 9179 35750 11229 35822
rect 9179 35698 9248 35750
rect 9300 35698 9372 35750
rect 9424 35698 9496 35750
rect 9548 35698 9620 35750
rect 9672 35698 9744 35750
rect 9796 35698 9868 35750
rect 9920 35698 9992 35750
rect 10044 35698 10116 35750
rect 10168 35698 10240 35750
rect 10292 35698 10364 35750
rect 10416 35698 10488 35750
rect 10540 35698 10612 35750
rect 10664 35698 10736 35750
rect 10788 35698 10860 35750
rect 10912 35698 10984 35750
rect 11036 35698 11108 35750
rect 11160 35698 11229 35750
rect 9179 35626 11229 35698
rect 9179 35574 9248 35626
rect 9300 35574 9372 35626
rect 9424 35574 9496 35626
rect 9548 35574 9620 35626
rect 9672 35574 9744 35626
rect 9796 35574 9868 35626
rect 9920 35574 9992 35626
rect 10044 35574 10116 35626
rect 10168 35574 10240 35626
rect 10292 35574 10364 35626
rect 10416 35574 10488 35626
rect 10540 35574 10612 35626
rect 10664 35574 10736 35626
rect 10788 35574 10860 35626
rect 10912 35574 10984 35626
rect 11036 35574 11108 35626
rect 11160 35574 11229 35626
rect 9179 35502 11229 35574
rect 9179 35450 9248 35502
rect 9300 35450 9372 35502
rect 9424 35450 9496 35502
rect 9548 35450 9620 35502
rect 9672 35450 9744 35502
rect 9796 35450 9868 35502
rect 9920 35450 9992 35502
rect 10044 35450 10116 35502
rect 10168 35450 10240 35502
rect 10292 35450 10364 35502
rect 10416 35450 10488 35502
rect 10540 35450 10612 35502
rect 10664 35450 10736 35502
rect 10788 35450 10860 35502
rect 10912 35450 10984 35502
rect 11036 35450 11108 35502
rect 11160 35450 11229 35502
rect 9179 35378 11229 35450
rect 9179 35326 9248 35378
rect 9300 35326 9372 35378
rect 9424 35326 9496 35378
rect 9548 35326 9620 35378
rect 9672 35326 9744 35378
rect 9796 35326 9868 35378
rect 9920 35326 9992 35378
rect 10044 35326 10116 35378
rect 10168 35326 10240 35378
rect 10292 35326 10364 35378
rect 10416 35326 10488 35378
rect 10540 35326 10612 35378
rect 10664 35326 10736 35378
rect 10788 35326 10860 35378
rect 10912 35326 10984 35378
rect 11036 35326 11108 35378
rect 11160 35326 11229 35378
rect 9179 29651 11229 35326
rect 9179 29599 9206 29651
rect 9258 29599 9314 29651
rect 9366 29599 9422 29651
rect 9474 29599 9530 29651
rect 9582 29599 9638 29651
rect 9690 29599 9746 29651
rect 9798 29599 9854 29651
rect 9906 29599 9962 29651
rect 10014 29599 10070 29651
rect 10122 29599 10178 29651
rect 10230 29599 10286 29651
rect 10338 29599 10394 29651
rect 10446 29599 10502 29651
rect 10554 29599 10610 29651
rect 10662 29599 10718 29651
rect 10770 29599 10826 29651
rect 10878 29599 10934 29651
rect 10986 29599 11042 29651
rect 11094 29599 11150 29651
rect 11202 29599 11229 29651
rect 9179 29543 11229 29599
rect 9179 29491 9206 29543
rect 9258 29491 9314 29543
rect 9366 29491 9422 29543
rect 9474 29491 9530 29543
rect 9582 29491 9638 29543
rect 9690 29491 9746 29543
rect 9798 29491 9854 29543
rect 9906 29491 9962 29543
rect 10014 29491 10070 29543
rect 10122 29491 10178 29543
rect 10230 29491 10286 29543
rect 10338 29491 10394 29543
rect 10446 29491 10502 29543
rect 10554 29491 10610 29543
rect 10662 29491 10718 29543
rect 10770 29491 10826 29543
rect 10878 29491 10934 29543
rect 10986 29491 11042 29543
rect 11094 29491 11150 29543
rect 11202 29491 11229 29543
rect 9179 27484 11229 29491
rect 9179 27432 9236 27484
rect 10224 27432 11229 27484
rect 9179 27155 11229 27432
rect 9179 25959 10634 27155
rect 10686 25959 11229 27155
rect 9179 25779 11229 25959
rect 9179 25727 9282 25779
rect 10686 25727 11229 25779
rect 9179 25617 11229 25727
rect 11289 45914 11489 46134
rect 11289 45862 11309 45914
rect 11361 45862 11417 45914
rect 11469 45862 11489 45914
rect 11289 42174 11489 45862
rect 11289 42122 11309 42174
rect 11361 42122 11417 42174
rect 11469 42122 11489 42174
rect 11289 29187 11489 42122
rect 11289 29135 11311 29187
rect 11467 29135 11489 29187
rect 11289 25617 11489 29135
rect 11809 25617 13709 46134
rect 1221 25597 1405 25609
rect 1221 25545 1233 25597
rect 1285 25545 1341 25597
rect 1393 25545 1405 25597
rect 1221 25489 1405 25545
rect 1221 25437 1233 25489
rect 1285 25437 1341 25489
rect 1393 25437 1405 25489
rect 1221 25425 1405 25437
rect 11557 25597 11741 25609
rect 11557 25545 11569 25597
rect 11621 25545 11677 25597
rect 11729 25545 11741 25597
rect 11557 25489 11741 25545
rect 11557 25437 11569 25489
rect 11621 25437 11677 25489
rect 11729 25437 11741 25489
rect 11557 25425 11741 25437
use comp018green_esd_rc_v5p0  comp018green_esd_rc_v5p0_0
timestamp 1758726819
transform 1 0 -356 0 -1 46507
box -51 491 13725 17038
use nmos_clamp_20_50_4_DVSS  nmos_clamp_20_50_4_DVSS_0
timestamp 1764277680
transform 1 0 0 0 1 0
box -747 -51 13709 25617
<< end >>
