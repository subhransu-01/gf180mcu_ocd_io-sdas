magic
tech gf180mcuD
magscale 1 10
timestamp 1764347740
<< nwell >>
rect -51 491 13725 4487
<< pwell >>
rect 2092 11351 4268 16351
rect 4528 11351 6704 16351
rect 6964 11351 9140 16351
rect 9400 11351 11576 16351
rect 2092 5339 4268 10339
rect 4528 5339 6704 10339
rect 6964 5339 9140 10339
rect 9400 5339 11576 10339
<< mvndiff >>
rect 2092 16314 2180 16351
rect 2092 11388 2105 16314
rect 2151 11388 2180 16314
rect 2092 11351 2180 11388
rect 4180 16314 4268 16351
rect 4180 11388 4209 16314
rect 4255 11388 4268 16314
rect 4180 11351 4268 11388
rect 4528 16314 4616 16351
rect 4528 11388 4541 16314
rect 4587 11388 4616 16314
rect 4528 11351 4616 11388
rect 6616 16314 6704 16351
rect 6616 11388 6645 16314
rect 6691 11388 6704 16314
rect 6616 11351 6704 11388
rect 6964 16314 7052 16351
rect 6964 11388 6977 16314
rect 7023 11388 7052 16314
rect 6964 11351 7052 11388
rect 9052 16314 9140 16351
rect 9052 11388 9081 16314
rect 9127 11388 9140 16314
rect 9052 11351 9140 11388
rect 9400 16314 9488 16351
rect 9400 11388 9413 16314
rect 9459 11388 9488 16314
rect 9400 11351 9488 11388
rect 11488 16314 11576 16351
rect 11488 11388 11517 16314
rect 11563 11388 11576 16314
rect 11488 11351 11576 11388
rect 2092 10302 2180 10339
rect 2092 5376 2105 10302
rect 2151 5376 2180 10302
rect 2092 5339 2180 5376
rect 4180 10302 4268 10339
rect 4180 5376 4209 10302
rect 4255 5376 4268 10302
rect 4180 5339 4268 5376
rect 4528 10302 4616 10339
rect 4528 5376 4541 10302
rect 4587 5376 4616 10302
rect 4528 5339 4616 5376
rect 6616 10302 6704 10339
rect 6616 5376 6645 10302
rect 6691 5376 6704 10302
rect 6616 5339 6704 5376
rect 6964 10302 7052 10339
rect 6964 5376 6977 10302
rect 7023 5376 7052 10302
rect 6964 5339 7052 5376
rect 9052 10302 9140 10339
rect 9052 5376 9081 10302
rect 9127 5376 9140 10302
rect 9052 5339 9140 5376
rect 9400 10302 9488 10339
rect 9400 5376 9413 10302
rect 9459 5376 9488 10302
rect 9400 5339 9488 5376
rect 11488 10302 11576 10339
rect 11488 5376 11517 10302
rect 11563 5376 11576 10302
rect 11488 5339 11576 5376
<< mvndiffc >>
rect 2105 11388 2151 16314
rect 4209 11388 4255 16314
rect 4541 11388 4587 16314
rect 6645 11388 6691 16314
rect 6977 11388 7023 16314
rect 9081 11388 9127 16314
rect 9413 11388 9459 16314
rect 11517 11388 11563 16314
rect 2105 5376 2151 10302
rect 4209 5376 4255 10302
rect 4541 5376 4587 10302
rect 6645 5376 6691 10302
rect 6977 5376 7023 10302
rect 9081 5376 9127 10302
rect 9413 5376 9459 10302
rect 11517 5376 11563 10302
<< psubdiff >>
rect 1565 17016 12109 17038
rect 1565 16970 1587 17016
rect 1633 16970 1701 17016
rect 1747 16970 1855 17016
rect 1901 16970 1969 17016
rect 2015 16970 2083 17016
rect 2129 16970 2197 17016
rect 2243 16970 2311 17016
rect 2357 16970 2425 17016
rect 2471 16970 2539 17016
rect 2585 16970 2653 17016
rect 2699 16970 2767 17016
rect 2813 16970 2881 17016
rect 2927 16970 2995 17016
rect 3041 16970 3109 17016
rect 3155 16970 3223 17016
rect 3269 16970 3337 17016
rect 3383 16970 3451 17016
rect 3497 16970 3565 17016
rect 3611 16970 3679 17016
rect 3725 16970 3793 17016
rect 3839 16970 3907 17016
rect 3953 16970 4021 17016
rect 4067 16970 4135 17016
rect 4181 16970 4249 17016
rect 4295 16970 4363 17016
rect 4409 16970 4477 17016
rect 4523 16970 4591 17016
rect 4637 16970 4705 17016
rect 4751 16970 4819 17016
rect 4865 16970 4933 17016
rect 4979 16970 5047 17016
rect 5093 16970 5161 17016
rect 5207 16970 5275 17016
rect 5321 16970 5389 17016
rect 5435 16970 5503 17016
rect 5549 16970 5617 17016
rect 5663 16970 5731 17016
rect 5777 16970 5845 17016
rect 5891 16970 5959 17016
rect 6005 16970 6073 17016
rect 6119 16970 6187 17016
rect 6233 16970 6301 17016
rect 6347 16970 6415 17016
rect 6461 16970 6529 17016
rect 6575 16970 6643 17016
rect 6689 16970 6757 17016
rect 6803 16970 6871 17016
rect 6917 16970 6985 17016
rect 7031 16970 7099 17016
rect 7145 16970 7213 17016
rect 7259 16970 7327 17016
rect 7373 16970 7441 17016
rect 7487 16970 7555 17016
rect 7601 16970 7669 17016
rect 7715 16970 7783 17016
rect 7829 16970 7897 17016
rect 7943 16970 8011 17016
rect 8057 16970 8125 17016
rect 8171 16970 8239 17016
rect 8285 16970 8353 17016
rect 8399 16970 8467 17016
rect 8513 16970 8581 17016
rect 8627 16970 8695 17016
rect 8741 16970 8809 17016
rect 8855 16970 8923 17016
rect 8969 16970 9037 17016
rect 9083 16970 9151 17016
rect 9197 16970 9265 17016
rect 9311 16970 9379 17016
rect 9425 16970 9493 17016
rect 9539 16970 9607 17016
rect 9653 16970 9721 17016
rect 9767 16970 9835 17016
rect 9881 16970 9949 17016
rect 9995 16970 10063 17016
rect 10109 16970 10177 17016
rect 10223 16970 10291 17016
rect 10337 16970 10405 17016
rect 10451 16970 10519 17016
rect 10565 16970 10633 17016
rect 10679 16970 10747 17016
rect 10793 16970 10861 17016
rect 10907 16970 10975 17016
rect 11021 16970 11089 17016
rect 11135 16970 11203 17016
rect 11249 16970 11317 17016
rect 11363 16970 11431 17016
rect 11477 16970 11545 17016
rect 11591 16970 11659 17016
rect 11705 16970 11773 17016
rect 11819 16970 11927 17016
rect 11973 16970 12041 17016
rect 12087 16970 12109 17016
rect 1565 16902 12109 16970
rect 1565 16856 1587 16902
rect 1633 16856 1701 16902
rect 1747 16856 1855 16902
rect 1901 16856 1969 16902
rect 2015 16856 2083 16902
rect 2129 16856 2197 16902
rect 2243 16856 2311 16902
rect 2357 16856 2425 16902
rect 2471 16856 2539 16902
rect 2585 16856 2653 16902
rect 2699 16856 2767 16902
rect 2813 16856 2881 16902
rect 2927 16856 2995 16902
rect 3041 16856 3109 16902
rect 3155 16856 3223 16902
rect 3269 16856 3337 16902
rect 3383 16856 3451 16902
rect 3497 16856 3565 16902
rect 3611 16856 3679 16902
rect 3725 16856 3793 16902
rect 3839 16856 3907 16902
rect 3953 16856 4021 16902
rect 4067 16856 4135 16902
rect 4181 16856 4249 16902
rect 4295 16856 4363 16902
rect 4409 16856 4477 16902
rect 4523 16856 4591 16902
rect 4637 16856 4705 16902
rect 4751 16856 4819 16902
rect 4865 16856 4933 16902
rect 4979 16856 5047 16902
rect 5093 16856 5161 16902
rect 5207 16856 5275 16902
rect 5321 16856 5389 16902
rect 5435 16856 5503 16902
rect 5549 16856 5617 16902
rect 5663 16856 5731 16902
rect 5777 16856 5845 16902
rect 5891 16856 5959 16902
rect 6005 16856 6073 16902
rect 6119 16856 6187 16902
rect 6233 16856 6301 16902
rect 6347 16856 6415 16902
rect 6461 16856 6529 16902
rect 6575 16856 6643 16902
rect 6689 16856 6757 16902
rect 6803 16856 6871 16902
rect 6917 16856 6985 16902
rect 7031 16856 7099 16902
rect 7145 16856 7213 16902
rect 7259 16856 7327 16902
rect 7373 16856 7441 16902
rect 7487 16856 7555 16902
rect 7601 16856 7669 16902
rect 7715 16856 7783 16902
rect 7829 16856 7897 16902
rect 7943 16856 8011 16902
rect 8057 16856 8125 16902
rect 8171 16856 8239 16902
rect 8285 16856 8353 16902
rect 8399 16856 8467 16902
rect 8513 16856 8581 16902
rect 8627 16856 8695 16902
rect 8741 16856 8809 16902
rect 8855 16856 8923 16902
rect 8969 16856 9037 16902
rect 9083 16856 9151 16902
rect 9197 16856 9265 16902
rect 9311 16856 9379 16902
rect 9425 16856 9493 16902
rect 9539 16856 9607 16902
rect 9653 16856 9721 16902
rect 9767 16856 9835 16902
rect 9881 16856 9949 16902
rect 9995 16856 10063 16902
rect 10109 16856 10177 16902
rect 10223 16856 10291 16902
rect 10337 16856 10405 16902
rect 10451 16856 10519 16902
rect 10565 16856 10633 16902
rect 10679 16856 10747 16902
rect 10793 16856 10861 16902
rect 10907 16856 10975 16902
rect 11021 16856 11089 16902
rect 11135 16856 11203 16902
rect 11249 16856 11317 16902
rect 11363 16856 11431 16902
rect 11477 16856 11545 16902
rect 11591 16856 11659 16902
rect 11705 16856 11773 16902
rect 11819 16856 11927 16902
rect 11973 16856 12041 16902
rect 12087 16856 12109 16902
rect 1565 16834 12109 16856
rect 1565 16788 1769 16834
rect 1565 16742 1587 16788
rect 1633 16742 1701 16788
rect 1747 16742 1769 16788
rect 1565 16218 1769 16742
rect 11905 16788 12109 16834
rect 11905 16742 11927 16788
rect 11973 16742 12041 16788
rect 12087 16742 12109 16788
rect 11905 16674 12109 16742
rect 11905 16628 11927 16674
rect 11973 16628 12041 16674
rect 12087 16628 12109 16674
rect 11905 16560 12109 16628
rect 11905 16514 11927 16560
rect 11973 16514 12041 16560
rect 12087 16514 12109 16560
rect 11905 16446 12109 16514
rect 11905 16400 11927 16446
rect 11973 16400 12041 16446
rect 12087 16400 12109 16446
rect 1565 16172 1587 16218
rect 1633 16172 1701 16218
rect 1747 16172 1769 16218
rect 1565 16104 1769 16172
rect 1565 16058 1587 16104
rect 1633 16058 1701 16104
rect 1747 16058 1769 16104
rect 1565 15990 1769 16058
rect 1565 15944 1587 15990
rect 1633 15944 1701 15990
rect 1747 15944 1769 15990
rect 1565 15876 1769 15944
rect 1565 15830 1587 15876
rect 1633 15830 1701 15876
rect 1747 15830 1769 15876
rect 1565 15762 1769 15830
rect 1565 15716 1587 15762
rect 1633 15716 1701 15762
rect 1747 15716 1769 15762
rect 1565 15648 1769 15716
rect 1565 15602 1587 15648
rect 1633 15602 1701 15648
rect 1747 15602 1769 15648
rect 1565 15534 1769 15602
rect 1565 15488 1587 15534
rect 1633 15488 1701 15534
rect 1747 15488 1769 15534
rect 1565 15420 1769 15488
rect 1565 15374 1587 15420
rect 1633 15374 1701 15420
rect 1747 15374 1769 15420
rect 1565 15306 1769 15374
rect 1565 15260 1587 15306
rect 1633 15260 1701 15306
rect 1747 15260 1769 15306
rect 1565 15192 1769 15260
rect 1565 15146 1587 15192
rect 1633 15146 1701 15192
rect 1747 15146 1769 15192
rect 1565 15078 1769 15146
rect 1565 15032 1587 15078
rect 1633 15032 1701 15078
rect 1747 15032 1769 15078
rect 1565 14964 1769 15032
rect 1565 14918 1587 14964
rect 1633 14918 1701 14964
rect 1747 14918 1769 14964
rect 1565 14850 1769 14918
rect 1565 14804 1587 14850
rect 1633 14804 1701 14850
rect 1747 14804 1769 14850
rect 1565 14736 1769 14804
rect 1565 14690 1587 14736
rect 1633 14690 1701 14736
rect 1747 14690 1769 14736
rect 1565 14622 1769 14690
rect 1565 14576 1587 14622
rect 1633 14576 1701 14622
rect 1747 14576 1769 14622
rect 1565 14508 1769 14576
rect 1565 14462 1587 14508
rect 1633 14462 1701 14508
rect 1747 14462 1769 14508
rect 1565 14394 1769 14462
rect 1565 14348 1587 14394
rect 1633 14348 1701 14394
rect 1747 14348 1769 14394
rect 1565 14280 1769 14348
rect 1565 14234 1587 14280
rect 1633 14234 1701 14280
rect 1747 14234 1769 14280
rect 1565 14166 1769 14234
rect 1565 14120 1587 14166
rect 1633 14120 1701 14166
rect 1747 14120 1769 14166
rect 1565 14052 1769 14120
rect 1565 14006 1587 14052
rect 1633 14006 1701 14052
rect 1747 14006 1769 14052
rect 1565 13938 1769 14006
rect 1565 13892 1587 13938
rect 1633 13892 1701 13938
rect 1747 13892 1769 13938
rect 1565 13824 1769 13892
rect 1565 13778 1587 13824
rect 1633 13778 1701 13824
rect 1747 13778 1769 13824
rect 1565 13710 1769 13778
rect 1565 13664 1587 13710
rect 1633 13664 1701 13710
rect 1747 13664 1769 13710
rect 1565 13596 1769 13664
rect 1565 13550 1587 13596
rect 1633 13550 1701 13596
rect 1747 13550 1769 13596
rect 1565 13482 1769 13550
rect 1565 13436 1587 13482
rect 1633 13436 1701 13482
rect 1747 13436 1769 13482
rect 1565 13368 1769 13436
rect 1565 13322 1587 13368
rect 1633 13322 1701 13368
rect 1747 13322 1769 13368
rect 1565 13254 1769 13322
rect 1565 13208 1587 13254
rect 1633 13208 1701 13254
rect 1747 13208 1769 13254
rect 1565 13140 1769 13208
rect 1565 13094 1587 13140
rect 1633 13094 1701 13140
rect 1747 13094 1769 13140
rect 1565 13026 1769 13094
rect 1565 12980 1587 13026
rect 1633 12980 1701 13026
rect 1747 12980 1769 13026
rect 1565 12912 1769 12980
rect 1565 12866 1587 12912
rect 1633 12866 1701 12912
rect 1747 12866 1769 12912
rect 1565 12798 1769 12866
rect 1565 12752 1587 12798
rect 1633 12752 1701 12798
rect 1747 12752 1769 12798
rect 1565 12684 1769 12752
rect 1565 12638 1587 12684
rect 1633 12638 1701 12684
rect 1747 12638 1769 12684
rect 1565 12570 1769 12638
rect 1565 12524 1587 12570
rect 1633 12524 1701 12570
rect 1747 12524 1769 12570
rect 1565 12456 1769 12524
rect 1565 12410 1587 12456
rect 1633 12410 1701 12456
rect 1747 12410 1769 12456
rect 1565 12342 1769 12410
rect 1565 12296 1587 12342
rect 1633 12296 1701 12342
rect 1747 12296 1769 12342
rect 1565 12228 1769 12296
rect 1565 12182 1587 12228
rect 1633 12182 1701 12228
rect 1747 12182 1769 12228
rect 1565 12114 1769 12182
rect 1565 12068 1587 12114
rect 1633 12068 1701 12114
rect 1747 12068 1769 12114
rect 1565 12000 1769 12068
rect 1565 11954 1587 12000
rect 1633 11954 1701 12000
rect 1747 11954 1769 12000
rect 1565 11886 1769 11954
rect 1565 11840 1587 11886
rect 1633 11840 1701 11886
rect 1747 11840 1769 11886
rect 1565 11772 1769 11840
rect 1565 11726 1587 11772
rect 1633 11726 1701 11772
rect 1747 11726 1769 11772
rect 1565 11658 1769 11726
rect 1565 11612 1587 11658
rect 1633 11612 1701 11658
rect 1747 11612 1769 11658
rect 1565 11544 1769 11612
rect 1565 11498 1587 11544
rect 1633 11498 1701 11544
rect 1747 11498 1769 11544
rect 1565 11430 1769 11498
rect 1565 11384 1587 11430
rect 1633 11384 1701 11430
rect 1747 11384 1769 11430
rect 1565 11316 1769 11384
rect 11905 16332 12109 16400
rect 11905 16286 11927 16332
rect 11973 16286 12041 16332
rect 12087 16286 12109 16332
rect 11905 16218 12109 16286
rect 11905 16172 11927 16218
rect 11973 16172 12041 16218
rect 12087 16172 12109 16218
rect 11905 16104 12109 16172
rect 11905 16058 11927 16104
rect 11973 16058 12041 16104
rect 12087 16058 12109 16104
rect 11905 15990 12109 16058
rect 11905 15944 11927 15990
rect 11973 15944 12041 15990
rect 12087 15944 12109 15990
rect 11905 15876 12109 15944
rect 11905 15830 11927 15876
rect 11973 15830 12041 15876
rect 12087 15830 12109 15876
rect 11905 15762 12109 15830
rect 11905 15716 11927 15762
rect 11973 15716 12041 15762
rect 12087 15716 12109 15762
rect 11905 15648 12109 15716
rect 11905 15602 11927 15648
rect 11973 15602 12041 15648
rect 12087 15602 12109 15648
rect 11905 15534 12109 15602
rect 11905 15488 11927 15534
rect 11973 15488 12041 15534
rect 12087 15488 12109 15534
rect 11905 15420 12109 15488
rect 11905 15374 11927 15420
rect 11973 15374 12041 15420
rect 12087 15374 12109 15420
rect 11905 15306 12109 15374
rect 11905 15260 11927 15306
rect 11973 15260 12041 15306
rect 12087 15260 12109 15306
rect 11905 15192 12109 15260
rect 11905 15146 11927 15192
rect 11973 15146 12041 15192
rect 12087 15146 12109 15192
rect 11905 15078 12109 15146
rect 11905 15032 11927 15078
rect 11973 15032 12041 15078
rect 12087 15032 12109 15078
rect 11905 14964 12109 15032
rect 11905 14918 11927 14964
rect 11973 14918 12041 14964
rect 12087 14918 12109 14964
rect 11905 14850 12109 14918
rect 11905 14804 11927 14850
rect 11973 14804 12041 14850
rect 12087 14804 12109 14850
rect 11905 14736 12109 14804
rect 11905 14690 11927 14736
rect 11973 14690 12041 14736
rect 12087 14690 12109 14736
rect 11905 14622 12109 14690
rect 11905 14576 11927 14622
rect 11973 14576 12041 14622
rect 12087 14576 12109 14622
rect 11905 14508 12109 14576
rect 11905 14462 11927 14508
rect 11973 14462 12041 14508
rect 12087 14462 12109 14508
rect 11905 14394 12109 14462
rect 11905 14348 11927 14394
rect 11973 14348 12041 14394
rect 12087 14348 12109 14394
rect 11905 14280 12109 14348
rect 11905 14234 11927 14280
rect 11973 14234 12041 14280
rect 12087 14234 12109 14280
rect 11905 14166 12109 14234
rect 11905 14120 11927 14166
rect 11973 14120 12041 14166
rect 12087 14120 12109 14166
rect 11905 14052 12109 14120
rect 11905 14006 11927 14052
rect 11973 14006 12041 14052
rect 12087 14006 12109 14052
rect 11905 13938 12109 14006
rect 11905 13892 11927 13938
rect 11973 13892 12041 13938
rect 12087 13892 12109 13938
rect 11905 13824 12109 13892
rect 11905 13778 11927 13824
rect 11973 13778 12041 13824
rect 12087 13778 12109 13824
rect 11905 13710 12109 13778
rect 11905 13664 11927 13710
rect 11973 13664 12041 13710
rect 12087 13664 12109 13710
rect 11905 13596 12109 13664
rect 11905 13550 11927 13596
rect 11973 13550 12041 13596
rect 12087 13550 12109 13596
rect 11905 13482 12109 13550
rect 11905 13436 11927 13482
rect 11973 13436 12041 13482
rect 12087 13436 12109 13482
rect 11905 13368 12109 13436
rect 11905 13322 11927 13368
rect 11973 13322 12041 13368
rect 12087 13322 12109 13368
rect 11905 13254 12109 13322
rect 11905 13208 11927 13254
rect 11973 13208 12041 13254
rect 12087 13208 12109 13254
rect 11905 13140 12109 13208
rect 11905 13094 11927 13140
rect 11973 13094 12041 13140
rect 12087 13094 12109 13140
rect 11905 13026 12109 13094
rect 11905 12980 11927 13026
rect 11973 12980 12041 13026
rect 12087 12980 12109 13026
rect 11905 12912 12109 12980
rect 11905 12866 11927 12912
rect 11973 12866 12041 12912
rect 12087 12866 12109 12912
rect 11905 12798 12109 12866
rect 11905 12752 11927 12798
rect 11973 12752 12041 12798
rect 12087 12752 12109 12798
rect 11905 12684 12109 12752
rect 11905 12638 11927 12684
rect 11973 12638 12041 12684
rect 12087 12638 12109 12684
rect 11905 12570 12109 12638
rect 11905 12524 11927 12570
rect 11973 12524 12041 12570
rect 12087 12524 12109 12570
rect 11905 12456 12109 12524
rect 11905 12410 11927 12456
rect 11973 12410 12041 12456
rect 12087 12410 12109 12456
rect 11905 12342 12109 12410
rect 11905 12296 11927 12342
rect 11973 12296 12041 12342
rect 12087 12296 12109 12342
rect 11905 12228 12109 12296
rect 11905 12182 11927 12228
rect 11973 12182 12041 12228
rect 12087 12182 12109 12228
rect 11905 12114 12109 12182
rect 11905 12068 11927 12114
rect 11973 12068 12041 12114
rect 12087 12068 12109 12114
rect 11905 12000 12109 12068
rect 11905 11954 11927 12000
rect 11973 11954 12041 12000
rect 12087 11954 12109 12000
rect 11905 11886 12109 11954
rect 11905 11840 11927 11886
rect 11973 11840 12041 11886
rect 12087 11840 12109 11886
rect 11905 11772 12109 11840
rect 11905 11726 11927 11772
rect 11973 11726 12041 11772
rect 12087 11726 12109 11772
rect 11905 11658 12109 11726
rect 11905 11612 11927 11658
rect 11973 11612 12041 11658
rect 12087 11612 12109 11658
rect 11905 11544 12109 11612
rect 11905 11498 11927 11544
rect 11973 11498 12041 11544
rect 12087 11498 12109 11544
rect 11905 11430 12109 11498
rect 11905 11384 11927 11430
rect 11973 11384 12041 11430
rect 12087 11384 12109 11430
rect 1565 11270 1587 11316
rect 1633 11270 1701 11316
rect 1747 11270 1769 11316
rect 1565 11202 1769 11270
rect 11905 11316 12109 11384
rect 11905 11270 11927 11316
rect 11973 11270 12041 11316
rect 12087 11270 12109 11316
rect 1565 11156 1587 11202
rect 1633 11156 1701 11202
rect 1747 11156 1769 11202
rect 1565 11088 1769 11156
rect 1565 11042 1587 11088
rect 1633 11042 1701 11088
rect 1747 11042 1769 11088
rect 1565 10974 1769 11042
rect 1565 10928 1587 10974
rect 1633 10928 1701 10974
rect 1747 10947 1769 10974
rect 11905 11202 12109 11270
rect 11905 11156 11927 11202
rect 11973 11156 12041 11202
rect 12087 11156 12109 11202
rect 11905 11088 12109 11156
rect 11905 11042 11927 11088
rect 11973 11042 12041 11088
rect 12087 11042 12109 11088
rect 11905 10974 12109 11042
rect 11905 10947 11927 10974
rect 1747 10928 11927 10947
rect 11973 10928 12041 10974
rect 12087 10928 12109 10974
rect 1565 10925 12109 10928
rect 1565 10879 1855 10925
rect 1901 10879 1969 10925
rect 2015 10879 2083 10925
rect 2129 10879 2197 10925
rect 2243 10879 2311 10925
rect 2357 10879 2425 10925
rect 2471 10879 2539 10925
rect 2585 10879 2653 10925
rect 2699 10879 2767 10925
rect 2813 10879 2881 10925
rect 2927 10879 2995 10925
rect 3041 10879 3109 10925
rect 3155 10879 3223 10925
rect 3269 10879 3337 10925
rect 3383 10879 3451 10925
rect 3497 10879 3565 10925
rect 3611 10879 3679 10925
rect 3725 10879 3793 10925
rect 3839 10879 3907 10925
rect 3953 10879 4021 10925
rect 4067 10879 4135 10925
rect 4181 10879 4249 10925
rect 4295 10879 4363 10925
rect 4409 10879 4477 10925
rect 4523 10879 4591 10925
rect 4637 10879 4705 10925
rect 4751 10879 4819 10925
rect 4865 10879 4933 10925
rect 4979 10879 5047 10925
rect 5093 10879 5161 10925
rect 5207 10879 5275 10925
rect 5321 10879 5389 10925
rect 5435 10879 5503 10925
rect 5549 10879 5617 10925
rect 5663 10879 5731 10925
rect 5777 10879 5845 10925
rect 5891 10879 5959 10925
rect 6005 10879 6073 10925
rect 6119 10879 6187 10925
rect 6233 10879 6301 10925
rect 6347 10879 6415 10925
rect 6461 10879 6529 10925
rect 6575 10879 6643 10925
rect 6689 10879 6757 10925
rect 6803 10879 6871 10925
rect 6917 10879 6985 10925
rect 7031 10879 7099 10925
rect 7145 10879 7213 10925
rect 7259 10879 7327 10925
rect 7373 10879 7441 10925
rect 7487 10879 7555 10925
rect 7601 10879 7669 10925
rect 7715 10879 7783 10925
rect 7829 10879 7897 10925
rect 7943 10879 8011 10925
rect 8057 10879 8125 10925
rect 8171 10879 8239 10925
rect 8285 10879 8353 10925
rect 8399 10879 8467 10925
rect 8513 10879 8581 10925
rect 8627 10879 8695 10925
rect 8741 10879 8809 10925
rect 8855 10879 8923 10925
rect 8969 10879 9037 10925
rect 9083 10879 9151 10925
rect 9197 10879 9265 10925
rect 9311 10879 9379 10925
rect 9425 10879 9493 10925
rect 9539 10879 9607 10925
rect 9653 10879 9721 10925
rect 9767 10879 9835 10925
rect 9881 10879 9949 10925
rect 9995 10879 10063 10925
rect 10109 10879 10177 10925
rect 10223 10879 10291 10925
rect 10337 10879 10405 10925
rect 10451 10879 10519 10925
rect 10565 10879 10633 10925
rect 10679 10879 10747 10925
rect 10793 10879 10861 10925
rect 10907 10879 10975 10925
rect 11021 10879 11089 10925
rect 11135 10879 11203 10925
rect 11249 10879 11317 10925
rect 11363 10879 11431 10925
rect 11477 10879 11545 10925
rect 11591 10879 11659 10925
rect 11705 10879 11773 10925
rect 11819 10879 12109 10925
rect 1565 10860 12109 10879
rect 1565 10814 1587 10860
rect 1633 10814 1701 10860
rect 1747 10814 11927 10860
rect 11973 10814 12041 10860
rect 12087 10814 12109 10860
rect 1565 10811 12109 10814
rect 1565 10765 1855 10811
rect 1901 10765 1969 10811
rect 2015 10765 2083 10811
rect 2129 10765 2197 10811
rect 2243 10765 2311 10811
rect 2357 10765 2425 10811
rect 2471 10765 2539 10811
rect 2585 10765 2653 10811
rect 2699 10765 2767 10811
rect 2813 10765 2881 10811
rect 2927 10765 2995 10811
rect 3041 10765 3109 10811
rect 3155 10765 3223 10811
rect 3269 10765 3337 10811
rect 3383 10765 3451 10811
rect 3497 10765 3565 10811
rect 3611 10765 3679 10811
rect 3725 10765 3793 10811
rect 3839 10765 3907 10811
rect 3953 10765 4021 10811
rect 4067 10765 4135 10811
rect 4181 10765 4249 10811
rect 4295 10765 4363 10811
rect 4409 10765 4477 10811
rect 4523 10765 4591 10811
rect 4637 10765 4705 10811
rect 4751 10765 4819 10811
rect 4865 10765 4933 10811
rect 4979 10765 5047 10811
rect 5093 10765 5161 10811
rect 5207 10765 5275 10811
rect 5321 10765 5389 10811
rect 5435 10765 5503 10811
rect 5549 10765 5617 10811
rect 5663 10765 5731 10811
rect 5777 10765 5845 10811
rect 5891 10765 5959 10811
rect 6005 10765 6073 10811
rect 6119 10765 6187 10811
rect 6233 10765 6301 10811
rect 6347 10765 6415 10811
rect 6461 10765 6529 10811
rect 6575 10765 6643 10811
rect 6689 10765 6757 10811
rect 6803 10765 6871 10811
rect 6917 10765 6985 10811
rect 7031 10765 7099 10811
rect 7145 10765 7213 10811
rect 7259 10765 7327 10811
rect 7373 10765 7441 10811
rect 7487 10765 7555 10811
rect 7601 10765 7669 10811
rect 7715 10765 7783 10811
rect 7829 10765 7897 10811
rect 7943 10765 8011 10811
rect 8057 10765 8125 10811
rect 8171 10765 8239 10811
rect 8285 10765 8353 10811
rect 8399 10765 8467 10811
rect 8513 10765 8581 10811
rect 8627 10765 8695 10811
rect 8741 10765 8809 10811
rect 8855 10765 8923 10811
rect 8969 10765 9037 10811
rect 9083 10765 9151 10811
rect 9197 10765 9265 10811
rect 9311 10765 9379 10811
rect 9425 10765 9493 10811
rect 9539 10765 9607 10811
rect 9653 10765 9721 10811
rect 9767 10765 9835 10811
rect 9881 10765 9949 10811
rect 9995 10765 10063 10811
rect 10109 10765 10177 10811
rect 10223 10765 10291 10811
rect 10337 10765 10405 10811
rect 10451 10765 10519 10811
rect 10565 10765 10633 10811
rect 10679 10765 10747 10811
rect 10793 10765 10861 10811
rect 10907 10765 10975 10811
rect 11021 10765 11089 10811
rect 11135 10765 11203 10811
rect 11249 10765 11317 10811
rect 11363 10765 11431 10811
rect 11477 10765 11545 10811
rect 11591 10765 11659 10811
rect 11705 10765 11773 10811
rect 11819 10765 12109 10811
rect 1565 10746 12109 10765
rect 1565 10700 1587 10746
rect 1633 10700 1701 10746
rect 1747 10743 11927 10746
rect 1747 10700 1769 10743
rect 1565 10632 1769 10700
rect 1565 10586 1587 10632
rect 1633 10586 1701 10632
rect 1747 10586 1769 10632
rect 1565 10518 1769 10586
rect 1565 10472 1587 10518
rect 1633 10472 1701 10518
rect 1747 10472 1769 10518
rect 1565 10404 1769 10472
rect 11905 10700 11927 10743
rect 11973 10700 12041 10746
rect 12087 10700 12109 10746
rect 11905 10632 12109 10700
rect 11905 10586 11927 10632
rect 11973 10586 12041 10632
rect 12087 10586 12109 10632
rect 11905 10518 12109 10586
rect 11905 10472 11927 10518
rect 11973 10472 12041 10518
rect 12087 10472 12109 10518
rect 1565 10358 1587 10404
rect 1633 10358 1701 10404
rect 1747 10358 1769 10404
rect 1565 10290 1769 10358
rect 11905 10404 12109 10472
rect 11905 10358 11927 10404
rect 11973 10358 12041 10404
rect 12087 10358 12109 10404
rect 1565 10244 1587 10290
rect 1633 10244 1701 10290
rect 1747 10244 1769 10290
rect 1565 10176 1769 10244
rect 1565 10130 1587 10176
rect 1633 10130 1701 10176
rect 1747 10130 1769 10176
rect 1565 10062 1769 10130
rect 1565 10016 1587 10062
rect 1633 10016 1701 10062
rect 1747 10016 1769 10062
rect 1565 9948 1769 10016
rect 1565 9902 1587 9948
rect 1633 9902 1701 9948
rect 1747 9902 1769 9948
rect 1565 9834 1769 9902
rect 1565 9788 1587 9834
rect 1633 9788 1701 9834
rect 1747 9788 1769 9834
rect 1565 9720 1769 9788
rect 1565 9674 1587 9720
rect 1633 9674 1701 9720
rect 1747 9674 1769 9720
rect 1565 9606 1769 9674
rect 1565 9560 1587 9606
rect 1633 9560 1701 9606
rect 1747 9560 1769 9606
rect 1565 9492 1769 9560
rect 1565 9446 1587 9492
rect 1633 9446 1701 9492
rect 1747 9446 1769 9492
rect 1565 9378 1769 9446
rect 1565 9332 1587 9378
rect 1633 9332 1701 9378
rect 1747 9332 1769 9378
rect 1565 9264 1769 9332
rect 1565 9218 1587 9264
rect 1633 9218 1701 9264
rect 1747 9218 1769 9264
rect 1565 9150 1769 9218
rect 1565 9104 1587 9150
rect 1633 9104 1701 9150
rect 1747 9104 1769 9150
rect 1565 9036 1769 9104
rect 1565 8990 1587 9036
rect 1633 8990 1701 9036
rect 1747 8990 1769 9036
rect 1565 8922 1769 8990
rect 1565 8876 1587 8922
rect 1633 8876 1701 8922
rect 1747 8876 1769 8922
rect 1565 8808 1769 8876
rect 1565 8762 1587 8808
rect 1633 8762 1701 8808
rect 1747 8762 1769 8808
rect 1565 8694 1769 8762
rect 1565 8648 1587 8694
rect 1633 8648 1701 8694
rect 1747 8648 1769 8694
rect 1565 8580 1769 8648
rect 1565 8534 1587 8580
rect 1633 8534 1701 8580
rect 1747 8534 1769 8580
rect 1565 8466 1769 8534
rect 1565 8420 1587 8466
rect 1633 8420 1701 8466
rect 1747 8420 1769 8466
rect 1565 8352 1769 8420
rect 1565 8306 1587 8352
rect 1633 8306 1701 8352
rect 1747 8306 1769 8352
rect 1565 8238 1769 8306
rect 1565 8192 1587 8238
rect 1633 8192 1701 8238
rect 1747 8192 1769 8238
rect 1565 8124 1769 8192
rect 1565 8078 1587 8124
rect 1633 8078 1701 8124
rect 1747 8078 1769 8124
rect 1565 8010 1769 8078
rect 1565 7964 1587 8010
rect 1633 7964 1701 8010
rect 1747 7964 1769 8010
rect 1565 7896 1769 7964
rect 1565 7850 1587 7896
rect 1633 7850 1701 7896
rect 1747 7850 1769 7896
rect 1565 7782 1769 7850
rect 1565 7736 1587 7782
rect 1633 7736 1701 7782
rect 1747 7736 1769 7782
rect 1565 7668 1769 7736
rect 1565 7622 1587 7668
rect 1633 7622 1701 7668
rect 1747 7622 1769 7668
rect 1565 7554 1769 7622
rect 1565 7508 1587 7554
rect 1633 7508 1701 7554
rect 1747 7508 1769 7554
rect 1565 7440 1769 7508
rect 1565 7394 1587 7440
rect 1633 7394 1701 7440
rect 1747 7394 1769 7440
rect 1565 7326 1769 7394
rect 1565 7280 1587 7326
rect 1633 7280 1701 7326
rect 1747 7280 1769 7326
rect 1565 7212 1769 7280
rect 1565 7166 1587 7212
rect 1633 7166 1701 7212
rect 1747 7166 1769 7212
rect 1565 7098 1769 7166
rect 1565 7052 1587 7098
rect 1633 7052 1701 7098
rect 1747 7052 1769 7098
rect 1565 6984 1769 7052
rect 1565 6938 1587 6984
rect 1633 6938 1701 6984
rect 1747 6938 1769 6984
rect 1565 6870 1769 6938
rect 1565 6824 1587 6870
rect 1633 6824 1701 6870
rect 1747 6824 1769 6870
rect 1565 6756 1769 6824
rect 1565 6710 1587 6756
rect 1633 6710 1701 6756
rect 1747 6710 1769 6756
rect 1565 6642 1769 6710
rect 1565 6596 1587 6642
rect 1633 6596 1701 6642
rect 1747 6596 1769 6642
rect 1565 6528 1769 6596
rect 1565 6482 1587 6528
rect 1633 6482 1701 6528
rect 1747 6482 1769 6528
rect 1565 6414 1769 6482
rect 1565 6368 1587 6414
rect 1633 6368 1701 6414
rect 1747 6368 1769 6414
rect 1565 6300 1769 6368
rect 1565 6254 1587 6300
rect 1633 6254 1701 6300
rect 1747 6254 1769 6300
rect 1565 6186 1769 6254
rect 1565 6140 1587 6186
rect 1633 6140 1701 6186
rect 1747 6140 1769 6186
rect 1565 6072 1769 6140
rect 1565 6026 1587 6072
rect 1633 6026 1701 6072
rect 1747 6026 1769 6072
rect 1565 5958 1769 6026
rect 1565 5912 1587 5958
rect 1633 5912 1701 5958
rect 1747 5912 1769 5958
rect 1565 5844 1769 5912
rect 1565 5798 1587 5844
rect 1633 5798 1701 5844
rect 1747 5798 1769 5844
rect 1565 5730 1769 5798
rect 1565 5684 1587 5730
rect 1633 5684 1701 5730
rect 1747 5684 1769 5730
rect 1565 5616 1769 5684
rect 1565 5570 1587 5616
rect 1633 5570 1701 5616
rect 1747 5570 1769 5616
rect 1565 5502 1769 5570
rect 1565 5456 1587 5502
rect 1633 5456 1701 5502
rect 1747 5456 1769 5502
rect 1565 5046 1769 5456
rect 11905 10290 12109 10358
rect 11905 10244 11927 10290
rect 11973 10244 12041 10290
rect 12087 10244 12109 10290
rect 11905 10176 12109 10244
rect 11905 10130 11927 10176
rect 11973 10130 12041 10176
rect 12087 10130 12109 10176
rect 11905 10062 12109 10130
rect 11905 10016 11927 10062
rect 11973 10016 12041 10062
rect 12087 10016 12109 10062
rect 11905 9948 12109 10016
rect 11905 9902 11927 9948
rect 11973 9902 12041 9948
rect 12087 9902 12109 9948
rect 11905 9834 12109 9902
rect 11905 9788 11927 9834
rect 11973 9788 12041 9834
rect 12087 9788 12109 9834
rect 11905 9720 12109 9788
rect 11905 9674 11927 9720
rect 11973 9674 12041 9720
rect 12087 9674 12109 9720
rect 11905 9606 12109 9674
rect 11905 9560 11927 9606
rect 11973 9560 12041 9606
rect 12087 9560 12109 9606
rect 11905 9492 12109 9560
rect 11905 9446 11927 9492
rect 11973 9446 12041 9492
rect 12087 9446 12109 9492
rect 11905 9378 12109 9446
rect 11905 9332 11927 9378
rect 11973 9332 12041 9378
rect 12087 9332 12109 9378
rect 11905 9264 12109 9332
rect 11905 9218 11927 9264
rect 11973 9218 12041 9264
rect 12087 9218 12109 9264
rect 11905 9150 12109 9218
rect 11905 9104 11927 9150
rect 11973 9104 12041 9150
rect 12087 9104 12109 9150
rect 11905 9036 12109 9104
rect 11905 8990 11927 9036
rect 11973 8990 12041 9036
rect 12087 8990 12109 9036
rect 11905 8922 12109 8990
rect 11905 8876 11927 8922
rect 11973 8876 12041 8922
rect 12087 8876 12109 8922
rect 11905 8808 12109 8876
rect 11905 8762 11927 8808
rect 11973 8762 12041 8808
rect 12087 8762 12109 8808
rect 11905 8694 12109 8762
rect 11905 8648 11927 8694
rect 11973 8648 12041 8694
rect 12087 8648 12109 8694
rect 11905 8580 12109 8648
rect 11905 8534 11927 8580
rect 11973 8534 12041 8580
rect 12087 8534 12109 8580
rect 11905 8466 12109 8534
rect 11905 8420 11927 8466
rect 11973 8420 12041 8466
rect 12087 8420 12109 8466
rect 11905 8352 12109 8420
rect 11905 8306 11927 8352
rect 11973 8306 12041 8352
rect 12087 8306 12109 8352
rect 11905 8238 12109 8306
rect 11905 8192 11927 8238
rect 11973 8192 12041 8238
rect 12087 8192 12109 8238
rect 11905 8124 12109 8192
rect 11905 8078 11927 8124
rect 11973 8078 12041 8124
rect 12087 8078 12109 8124
rect 11905 8010 12109 8078
rect 11905 7964 11927 8010
rect 11973 7964 12041 8010
rect 12087 7964 12109 8010
rect 11905 7896 12109 7964
rect 11905 7850 11927 7896
rect 11973 7850 12041 7896
rect 12087 7850 12109 7896
rect 11905 7782 12109 7850
rect 11905 7736 11927 7782
rect 11973 7736 12041 7782
rect 12087 7736 12109 7782
rect 11905 7668 12109 7736
rect 11905 7622 11927 7668
rect 11973 7622 12041 7668
rect 12087 7622 12109 7668
rect 11905 7554 12109 7622
rect 11905 7508 11927 7554
rect 11973 7508 12041 7554
rect 12087 7508 12109 7554
rect 11905 7440 12109 7508
rect 11905 7394 11927 7440
rect 11973 7394 12041 7440
rect 12087 7394 12109 7440
rect 11905 7326 12109 7394
rect 11905 7280 11927 7326
rect 11973 7280 12041 7326
rect 12087 7280 12109 7326
rect 11905 7212 12109 7280
rect 11905 7166 11927 7212
rect 11973 7166 12041 7212
rect 12087 7166 12109 7212
rect 11905 7098 12109 7166
rect 11905 7052 11927 7098
rect 11973 7052 12041 7098
rect 12087 7052 12109 7098
rect 11905 6984 12109 7052
rect 11905 6938 11927 6984
rect 11973 6938 12041 6984
rect 12087 6938 12109 6984
rect 11905 6870 12109 6938
rect 11905 6824 11927 6870
rect 11973 6824 12041 6870
rect 12087 6824 12109 6870
rect 11905 6756 12109 6824
rect 11905 6710 11927 6756
rect 11973 6710 12041 6756
rect 12087 6710 12109 6756
rect 11905 6642 12109 6710
rect 11905 6596 11927 6642
rect 11973 6596 12041 6642
rect 12087 6596 12109 6642
rect 11905 6528 12109 6596
rect 11905 6482 11927 6528
rect 11973 6482 12041 6528
rect 12087 6482 12109 6528
rect 11905 6414 12109 6482
rect 11905 6368 11927 6414
rect 11973 6368 12041 6414
rect 12087 6368 12109 6414
rect 11905 6300 12109 6368
rect 11905 6254 11927 6300
rect 11973 6254 12041 6300
rect 12087 6254 12109 6300
rect 11905 6186 12109 6254
rect 11905 6140 11927 6186
rect 11973 6140 12041 6186
rect 12087 6140 12109 6186
rect 11905 6072 12109 6140
rect 11905 6026 11927 6072
rect 11973 6026 12041 6072
rect 12087 6026 12109 6072
rect 11905 5958 12109 6026
rect 11905 5912 11927 5958
rect 11973 5912 12041 5958
rect 12087 5912 12109 5958
rect 11905 5844 12109 5912
rect 11905 5798 11927 5844
rect 11973 5798 12041 5844
rect 12087 5798 12109 5844
rect 11905 5730 12109 5798
rect 11905 5684 11927 5730
rect 11973 5684 12041 5730
rect 12087 5684 12109 5730
rect 11905 5616 12109 5684
rect 11905 5570 11927 5616
rect 11973 5570 12041 5616
rect 12087 5570 12109 5616
rect 11905 5502 12109 5570
rect 11905 5456 11927 5502
rect 11973 5456 12041 5502
rect 12087 5456 12109 5502
rect 11905 5388 12109 5456
rect 11905 5342 11927 5388
rect 11973 5342 12041 5388
rect 12087 5342 12109 5388
rect 11905 5274 12109 5342
rect 1565 5000 1587 5046
rect 1633 5000 1701 5046
rect 1747 5000 1769 5046
rect 1565 4954 1769 5000
rect 11905 5228 11927 5274
rect 11973 5228 12041 5274
rect 12087 5228 12109 5274
rect 11905 5160 12109 5228
rect 11905 5114 11927 5160
rect 11973 5114 12041 5160
rect 12087 5114 12109 5160
rect 11905 5046 12109 5114
rect 11905 5000 11927 5046
rect 11973 5000 12041 5046
rect 12087 5000 12109 5046
rect 11905 4954 12109 5000
rect 1565 4932 12109 4954
rect 1565 4886 1587 4932
rect 1633 4886 1701 4932
rect 1747 4886 1855 4932
rect 1901 4886 1969 4932
rect 2015 4886 2083 4932
rect 2129 4886 2197 4932
rect 2243 4886 2311 4932
rect 2357 4886 2425 4932
rect 2471 4886 2539 4932
rect 2585 4886 2653 4932
rect 2699 4886 2767 4932
rect 2813 4886 2881 4932
rect 2927 4886 2995 4932
rect 3041 4886 3109 4932
rect 3155 4886 3223 4932
rect 3269 4886 3337 4932
rect 3383 4886 3451 4932
rect 3497 4886 3565 4932
rect 3611 4886 3679 4932
rect 3725 4886 3793 4932
rect 3839 4886 3907 4932
rect 3953 4886 4021 4932
rect 4067 4886 4135 4932
rect 4181 4886 4249 4932
rect 4295 4886 4363 4932
rect 4409 4886 4477 4932
rect 4523 4886 4591 4932
rect 4637 4886 4705 4932
rect 4751 4886 4819 4932
rect 4865 4886 4933 4932
rect 4979 4886 5047 4932
rect 5093 4886 5161 4932
rect 5207 4886 5275 4932
rect 5321 4886 5389 4932
rect 5435 4886 5503 4932
rect 5549 4886 5617 4932
rect 5663 4886 5731 4932
rect 5777 4886 5845 4932
rect 5891 4886 5959 4932
rect 6005 4886 6073 4932
rect 6119 4886 6187 4932
rect 6233 4886 6301 4932
rect 6347 4886 6415 4932
rect 6461 4886 6529 4932
rect 6575 4886 6643 4932
rect 6689 4886 6757 4932
rect 6803 4886 6871 4932
rect 6917 4886 6985 4932
rect 7031 4886 7099 4932
rect 7145 4886 7213 4932
rect 7259 4886 7327 4932
rect 7373 4886 7441 4932
rect 7487 4886 7555 4932
rect 7601 4886 7669 4932
rect 7715 4886 7783 4932
rect 7829 4886 7897 4932
rect 7943 4886 8011 4932
rect 8057 4886 8125 4932
rect 8171 4886 8239 4932
rect 8285 4886 8353 4932
rect 8399 4886 8467 4932
rect 8513 4886 8581 4932
rect 8627 4886 8695 4932
rect 8741 4886 8809 4932
rect 8855 4886 8923 4932
rect 8969 4886 9037 4932
rect 9083 4886 9151 4932
rect 9197 4886 9265 4932
rect 9311 4886 9379 4932
rect 9425 4886 9493 4932
rect 9539 4886 9607 4932
rect 9653 4886 9721 4932
rect 9767 4886 9835 4932
rect 9881 4886 9949 4932
rect 9995 4886 10063 4932
rect 10109 4886 10177 4932
rect 10223 4886 10291 4932
rect 10337 4886 10405 4932
rect 10451 4886 10519 4932
rect 10565 4886 10633 4932
rect 10679 4886 10747 4932
rect 10793 4886 10861 4932
rect 10907 4886 10975 4932
rect 11021 4886 11089 4932
rect 11135 4886 11203 4932
rect 11249 4886 11317 4932
rect 11363 4886 11431 4932
rect 11477 4886 11545 4932
rect 11591 4886 11659 4932
rect 11705 4886 11773 4932
rect 11819 4886 11927 4932
rect 11973 4886 12041 4932
rect 12087 4886 12109 4932
rect 1565 4818 12109 4886
rect 1565 4772 1587 4818
rect 1633 4772 1701 4818
rect 1747 4772 1855 4818
rect 1901 4772 1969 4818
rect 2015 4772 2083 4818
rect 2129 4772 2197 4818
rect 2243 4772 2311 4818
rect 2357 4772 2425 4818
rect 2471 4772 2539 4818
rect 2585 4772 2653 4818
rect 2699 4772 2767 4818
rect 2813 4772 2881 4818
rect 2927 4772 2995 4818
rect 3041 4772 3109 4818
rect 3155 4772 3223 4818
rect 3269 4772 3337 4818
rect 3383 4772 3451 4818
rect 3497 4772 3565 4818
rect 3611 4772 3679 4818
rect 3725 4772 3793 4818
rect 3839 4772 3907 4818
rect 3953 4772 4021 4818
rect 4067 4772 4135 4818
rect 4181 4772 4249 4818
rect 4295 4772 4363 4818
rect 4409 4772 4477 4818
rect 4523 4772 4591 4818
rect 4637 4772 4705 4818
rect 4751 4772 4819 4818
rect 4865 4772 4933 4818
rect 4979 4772 5047 4818
rect 5093 4772 5161 4818
rect 5207 4772 5275 4818
rect 5321 4772 5389 4818
rect 5435 4772 5503 4818
rect 5549 4772 5617 4818
rect 5663 4772 5731 4818
rect 5777 4772 5845 4818
rect 5891 4772 5959 4818
rect 6005 4772 6073 4818
rect 6119 4772 6187 4818
rect 6233 4772 6301 4818
rect 6347 4772 6415 4818
rect 6461 4772 6529 4818
rect 6575 4772 6643 4818
rect 6689 4772 6757 4818
rect 6803 4772 6871 4818
rect 6917 4772 6985 4818
rect 7031 4772 7099 4818
rect 7145 4772 7213 4818
rect 7259 4772 7327 4818
rect 7373 4772 7441 4818
rect 7487 4772 7555 4818
rect 7601 4772 7669 4818
rect 7715 4772 7783 4818
rect 7829 4772 7897 4818
rect 7943 4772 8011 4818
rect 8057 4772 8125 4818
rect 8171 4772 8239 4818
rect 8285 4772 8353 4818
rect 8399 4772 8467 4818
rect 8513 4772 8581 4818
rect 8627 4772 8695 4818
rect 8741 4772 8809 4818
rect 8855 4772 8923 4818
rect 8969 4772 9037 4818
rect 9083 4772 9151 4818
rect 9197 4772 9265 4818
rect 9311 4772 9379 4818
rect 9425 4772 9493 4818
rect 9539 4772 9607 4818
rect 9653 4772 9721 4818
rect 9767 4772 9835 4818
rect 9881 4772 9949 4818
rect 9995 4772 10063 4818
rect 10109 4772 10177 4818
rect 10223 4772 10291 4818
rect 10337 4772 10405 4818
rect 10451 4772 10519 4818
rect 10565 4772 10633 4818
rect 10679 4772 10747 4818
rect 10793 4772 10861 4818
rect 10907 4772 10975 4818
rect 11021 4772 11089 4818
rect 11135 4772 11203 4818
rect 11249 4772 11317 4818
rect 11363 4772 11431 4818
rect 11477 4772 11545 4818
rect 11591 4772 11659 4818
rect 11705 4772 11773 4818
rect 11819 4772 11927 4818
rect 11973 4772 12041 4818
rect 12087 4772 12109 4818
rect 1565 4750 12109 4772
<< nsubdiff >>
rect 32 4382 13642 4404
rect 32 4336 54 4382
rect 100 4336 158 4382
rect 204 4336 574 4382
rect 620 4336 678 4382
rect 724 4336 782 4382
rect 828 4336 886 4382
rect 932 4336 990 4382
rect 1036 4336 1094 4382
rect 1140 4336 1198 4382
rect 1244 4336 1302 4382
rect 1348 4336 1406 4382
rect 1452 4336 1510 4382
rect 1556 4336 1614 4382
rect 1660 4336 1718 4382
rect 1764 4336 1822 4382
rect 1868 4336 1926 4382
rect 1972 4336 2030 4382
rect 2076 4336 2134 4382
rect 2180 4336 2238 4382
rect 2284 4336 2342 4382
rect 2388 4336 2446 4382
rect 2492 4336 2550 4382
rect 2596 4336 2654 4382
rect 2700 4336 2758 4382
rect 2804 4336 2862 4382
rect 2908 4336 2966 4382
rect 3012 4336 3070 4382
rect 3116 4336 3174 4382
rect 3220 4336 3278 4382
rect 3324 4336 3382 4382
rect 3428 4336 3486 4382
rect 3532 4336 3590 4382
rect 3636 4336 3694 4382
rect 3740 4336 3798 4382
rect 3844 4336 3902 4382
rect 3948 4336 4006 4382
rect 4052 4336 4110 4382
rect 4156 4336 4214 4382
rect 4260 4336 4318 4382
rect 4364 4336 4422 4382
rect 4468 4336 4526 4382
rect 4572 4336 4630 4382
rect 4676 4336 4734 4382
rect 4780 4336 4838 4382
rect 4884 4336 4942 4382
rect 4988 4336 5046 4382
rect 5092 4336 5150 4382
rect 5196 4336 5254 4382
rect 5300 4336 5358 4382
rect 5404 4336 5462 4382
rect 5508 4336 5566 4382
rect 5612 4336 5670 4382
rect 5716 4336 5774 4382
rect 5820 4336 5878 4382
rect 5924 4336 5982 4382
rect 6028 4336 6086 4382
rect 6132 4336 6190 4382
rect 6236 4336 6294 4382
rect 6340 4336 6398 4382
rect 6444 4336 6502 4382
rect 6548 4336 6606 4382
rect 6652 4336 6710 4382
rect 6756 4336 6814 4382
rect 6860 4336 6918 4382
rect 6964 4336 7022 4382
rect 7068 4336 7126 4382
rect 7172 4336 7230 4382
rect 7276 4336 7334 4382
rect 7380 4336 7438 4382
rect 7484 4336 7542 4382
rect 7588 4336 7646 4382
rect 7692 4336 7750 4382
rect 7796 4336 7854 4382
rect 7900 4336 7958 4382
rect 8004 4336 8062 4382
rect 8108 4336 8166 4382
rect 8212 4336 8270 4382
rect 8316 4336 8374 4382
rect 8420 4336 8478 4382
rect 8524 4336 8582 4382
rect 8628 4336 8686 4382
rect 8732 4336 8790 4382
rect 8836 4336 8894 4382
rect 8940 4336 8998 4382
rect 9044 4336 9102 4382
rect 9148 4336 9206 4382
rect 9252 4336 9310 4382
rect 9356 4336 9414 4382
rect 9460 4336 9518 4382
rect 9564 4336 9622 4382
rect 9668 4336 9726 4382
rect 9772 4336 9830 4382
rect 9876 4336 9934 4382
rect 9980 4336 10038 4382
rect 10084 4336 10142 4382
rect 10188 4336 10246 4382
rect 10292 4336 10350 4382
rect 10396 4336 10454 4382
rect 10500 4336 10558 4382
rect 10604 4336 10662 4382
rect 10708 4336 10766 4382
rect 10812 4336 10870 4382
rect 10916 4336 10974 4382
rect 11020 4336 11078 4382
rect 11124 4336 11182 4382
rect 11228 4336 11286 4382
rect 11332 4336 11390 4382
rect 11436 4336 11494 4382
rect 11540 4336 11598 4382
rect 11644 4336 11702 4382
rect 11748 4336 11806 4382
rect 11852 4336 11910 4382
rect 11956 4336 12014 4382
rect 12060 4336 12118 4382
rect 12164 4336 12222 4382
rect 12268 4336 12326 4382
rect 12372 4336 12430 4382
rect 12476 4336 12534 4382
rect 12580 4336 12638 4382
rect 12684 4336 12742 4382
rect 12788 4336 12846 4382
rect 12892 4336 12950 4382
rect 12996 4336 13054 4382
rect 13100 4336 13158 4382
rect 13204 4336 13262 4382
rect 13308 4336 13366 4382
rect 13412 4336 13470 4382
rect 13516 4336 13574 4382
rect 13620 4336 13642 4382
rect 32 4314 13642 4336
rect 32 4228 122 4314
rect 32 4182 54 4228
rect 100 4182 122 4228
rect 32 4124 122 4182
rect 32 4078 54 4124
rect 100 4078 122 4124
rect 13552 4228 13642 4314
rect 13552 4182 13574 4228
rect 13620 4182 13642 4228
rect 13552 4124 13642 4182
rect 32 4020 122 4078
rect 32 3974 54 4020
rect 100 3974 122 4020
rect 32 3916 122 3974
rect 13552 4078 13574 4124
rect 13620 4078 13642 4124
rect 13552 4020 13642 4078
rect 13552 3974 13574 4020
rect 13620 3974 13642 4020
rect 32 3870 54 3916
rect 100 3870 122 3916
rect 32 3812 122 3870
rect 13552 3916 13642 3974
rect 13552 3870 13574 3916
rect 13620 3870 13642 3916
rect 32 3766 54 3812
rect 100 3766 122 3812
rect 32 3708 122 3766
rect 32 3662 54 3708
rect 100 3662 122 3708
rect 13552 3812 13642 3870
rect 13552 3766 13574 3812
rect 13620 3766 13642 3812
rect 13552 3708 13642 3766
rect 32 3604 122 3662
rect 32 3558 54 3604
rect 100 3558 122 3604
rect 32 3500 122 3558
rect 13552 3662 13574 3708
rect 13620 3662 13642 3708
rect 13552 3604 13642 3662
rect 13552 3558 13574 3604
rect 13620 3558 13642 3604
rect 32 3454 54 3500
rect 100 3454 122 3500
rect 32 3396 122 3454
rect 32 3350 54 3396
rect 100 3350 122 3396
rect 13552 3500 13642 3558
rect 13552 3454 13574 3500
rect 13620 3454 13642 3500
rect 13552 3396 13642 3454
rect 32 3292 122 3350
rect 32 3246 54 3292
rect 100 3246 122 3292
rect 13552 3350 13574 3396
rect 13620 3350 13642 3396
rect 13552 3292 13642 3350
rect 32 3188 122 3246
rect 32 3142 54 3188
rect 100 3142 122 3188
rect 32 3084 122 3142
rect 13552 3246 13574 3292
rect 13620 3246 13642 3292
rect 13552 3188 13642 3246
rect 13552 3142 13574 3188
rect 13620 3142 13642 3188
rect 32 3038 54 3084
rect 100 3038 122 3084
rect 32 2980 122 3038
rect 13552 3084 13642 3142
rect 13552 3038 13574 3084
rect 13620 3038 13642 3084
rect 32 2934 54 2980
rect 100 2934 122 2980
rect 32 2876 122 2934
rect 32 2830 54 2876
rect 100 2830 122 2876
rect 32 2772 122 2830
rect 13552 2980 13642 3038
rect 13552 2934 13574 2980
rect 13620 2934 13642 2980
rect 13552 2876 13642 2934
rect 13552 2830 13574 2876
rect 13620 2830 13642 2876
rect 32 2726 54 2772
rect 100 2726 122 2772
rect 32 2668 122 2726
rect 13552 2772 13642 2830
rect 13552 2726 13574 2772
rect 13620 2726 13642 2772
rect 32 2622 54 2668
rect 100 2622 122 2668
rect 32 2564 122 2622
rect 32 2518 54 2564
rect 100 2518 122 2564
rect 13552 2668 13642 2726
rect 13552 2622 13574 2668
rect 13620 2622 13642 2668
rect 13552 2564 13642 2622
rect 32 2460 122 2518
rect 32 2414 54 2460
rect 100 2414 122 2460
rect 13552 2518 13574 2564
rect 13620 2518 13642 2564
rect 13552 2460 13642 2518
rect 32 2356 122 2414
rect 32 2310 54 2356
rect 100 2310 122 2356
rect 32 2252 122 2310
rect 13552 2414 13574 2460
rect 13620 2414 13642 2460
rect 13552 2356 13642 2414
rect 13552 2310 13574 2356
rect 13620 2310 13642 2356
rect 32 2206 54 2252
rect 100 2206 122 2252
rect 32 2148 122 2206
rect 13552 2252 13642 2310
rect 13552 2206 13574 2252
rect 13620 2206 13642 2252
rect 32 2102 54 2148
rect 100 2102 122 2148
rect 32 2044 122 2102
rect 32 1998 54 2044
rect 100 1998 122 2044
rect 32 1940 122 1998
rect 13552 2148 13642 2206
rect 13552 2102 13574 2148
rect 13620 2102 13642 2148
rect 13552 2044 13642 2102
rect 13552 1998 13574 2044
rect 13620 1998 13642 2044
rect 32 1894 54 1940
rect 100 1894 122 1940
rect 32 1836 122 1894
rect 13552 1940 13642 1998
rect 13552 1894 13574 1940
rect 13620 1894 13642 1940
rect 32 1790 54 1836
rect 100 1790 122 1836
rect 32 1732 122 1790
rect 32 1686 54 1732
rect 100 1686 122 1732
rect 13552 1836 13642 1894
rect 13552 1790 13574 1836
rect 13620 1790 13642 1836
rect 13552 1732 13642 1790
rect 32 1628 122 1686
rect 32 1582 54 1628
rect 100 1582 122 1628
rect 13552 1686 13574 1732
rect 13620 1686 13642 1732
rect 13552 1628 13642 1686
rect 32 1524 122 1582
rect 32 1478 54 1524
rect 100 1478 122 1524
rect 32 1420 122 1478
rect 13552 1582 13574 1628
rect 13620 1582 13642 1628
rect 13552 1524 13642 1582
rect 13552 1478 13574 1524
rect 13620 1478 13642 1524
rect 32 1374 54 1420
rect 100 1374 122 1420
rect 32 1316 122 1374
rect 32 1270 54 1316
rect 100 1270 122 1316
rect 13552 1420 13642 1478
rect 13552 1374 13574 1420
rect 13620 1374 13642 1420
rect 13552 1316 13642 1374
rect 32 1212 122 1270
rect 32 1166 54 1212
rect 100 1166 122 1212
rect 32 1108 122 1166
rect 13552 1270 13574 1316
rect 13620 1270 13642 1316
rect 13552 1212 13642 1270
rect 13552 1166 13574 1212
rect 13620 1166 13642 1212
rect 32 1062 54 1108
rect 100 1062 122 1108
rect 32 1004 122 1062
rect 13552 1108 13642 1166
rect 13552 1062 13574 1108
rect 13620 1062 13642 1108
rect 32 958 54 1004
rect 100 958 122 1004
rect 32 900 122 958
rect 32 854 54 900
rect 100 854 122 900
rect 13552 1004 13642 1062
rect 13552 958 13574 1004
rect 13620 958 13642 1004
rect 13552 900 13642 958
rect 32 796 122 854
rect 32 750 54 796
rect 100 750 122 796
rect 32 664 122 750
rect 13552 854 13574 900
rect 13620 854 13642 900
rect 13552 796 13642 854
rect 13552 750 13574 796
rect 13620 750 13642 796
rect 13552 664 13642 750
rect 32 642 13642 664
rect 32 596 54 642
rect 100 596 158 642
rect 204 596 262 642
rect 308 596 366 642
rect 412 596 470 642
rect 516 596 574 642
rect 620 596 678 642
rect 724 596 782 642
rect 828 596 886 642
rect 932 596 990 642
rect 1036 596 1094 642
rect 1140 596 1198 642
rect 1244 596 1302 642
rect 1348 596 1406 642
rect 1452 596 1510 642
rect 1556 596 1614 642
rect 1660 596 1718 642
rect 1764 596 1822 642
rect 1868 596 1926 642
rect 1972 596 2030 642
rect 2076 596 2134 642
rect 2180 596 2238 642
rect 2284 596 2342 642
rect 2388 596 2446 642
rect 2492 596 2550 642
rect 2596 596 2654 642
rect 2700 596 2758 642
rect 2804 596 2862 642
rect 2908 596 2966 642
rect 3012 596 3070 642
rect 3116 596 3174 642
rect 3220 596 3278 642
rect 3324 596 3382 642
rect 3428 596 3486 642
rect 3532 596 3590 642
rect 3636 596 3694 642
rect 3740 596 3798 642
rect 3844 596 3902 642
rect 3948 596 4006 642
rect 4052 596 4110 642
rect 4156 596 4214 642
rect 4260 596 4318 642
rect 4364 596 4422 642
rect 4468 596 4526 642
rect 4572 596 4630 642
rect 4676 596 4734 642
rect 4780 596 4838 642
rect 4884 596 4942 642
rect 4988 596 5046 642
rect 5092 596 5150 642
rect 5196 596 5254 642
rect 5300 596 5358 642
rect 5404 596 5462 642
rect 5508 596 5566 642
rect 5612 596 5670 642
rect 5716 596 5774 642
rect 5820 596 5878 642
rect 5924 596 5982 642
rect 6028 596 6086 642
rect 6132 596 6190 642
rect 6236 596 6294 642
rect 6340 596 6398 642
rect 6444 596 6502 642
rect 6548 596 6606 642
rect 6652 596 6710 642
rect 6756 596 6814 642
rect 6860 596 6918 642
rect 6964 596 7022 642
rect 7068 596 7126 642
rect 7172 596 7230 642
rect 7276 596 7334 642
rect 7380 596 7438 642
rect 7484 596 7542 642
rect 7588 596 7646 642
rect 7692 596 7750 642
rect 7796 596 7854 642
rect 7900 596 7958 642
rect 8004 596 8062 642
rect 8108 596 8166 642
rect 8212 596 8270 642
rect 8316 596 8374 642
rect 8420 596 8478 642
rect 8524 596 8582 642
rect 8628 596 8686 642
rect 8732 596 8790 642
rect 8836 596 8894 642
rect 8940 596 8998 642
rect 9044 596 9102 642
rect 9148 596 9206 642
rect 9252 596 9310 642
rect 9356 596 9414 642
rect 9460 596 9518 642
rect 9564 596 9622 642
rect 9668 596 9726 642
rect 9772 596 9830 642
rect 9876 596 9934 642
rect 9980 596 10038 642
rect 10084 596 10142 642
rect 10188 596 10246 642
rect 10292 596 10350 642
rect 10396 596 10454 642
rect 10500 596 10558 642
rect 10604 596 10662 642
rect 10708 596 10766 642
rect 10812 596 10870 642
rect 10916 596 10974 642
rect 11020 596 11078 642
rect 11124 596 11182 642
rect 11228 596 11286 642
rect 11332 596 11390 642
rect 11436 596 11494 642
rect 11540 596 11598 642
rect 11644 596 11702 642
rect 11748 596 11806 642
rect 11852 596 11910 642
rect 11956 596 12014 642
rect 12060 596 12118 642
rect 12164 596 12222 642
rect 12268 596 12326 642
rect 12372 596 12430 642
rect 12476 596 12534 642
rect 12580 596 12638 642
rect 12684 596 12742 642
rect 12788 596 12846 642
rect 12892 596 12950 642
rect 12996 596 13054 642
rect 13100 596 13158 642
rect 13204 596 13262 642
rect 13308 596 13366 642
rect 13412 596 13470 642
rect 13516 596 13574 642
rect 13620 596 13642 642
rect 32 574 13642 596
<< psubdiffcont >>
rect 1587 16970 1633 17016
rect 1701 16970 1747 17016
rect 1855 16970 1901 17016
rect 1969 16970 2015 17016
rect 2083 16970 2129 17016
rect 2197 16970 2243 17016
rect 2311 16970 2357 17016
rect 2425 16970 2471 17016
rect 2539 16970 2585 17016
rect 2653 16970 2699 17016
rect 2767 16970 2813 17016
rect 2881 16970 2927 17016
rect 2995 16970 3041 17016
rect 3109 16970 3155 17016
rect 3223 16970 3269 17016
rect 3337 16970 3383 17016
rect 3451 16970 3497 17016
rect 3565 16970 3611 17016
rect 3679 16970 3725 17016
rect 3793 16970 3839 17016
rect 3907 16970 3953 17016
rect 4021 16970 4067 17016
rect 4135 16970 4181 17016
rect 4249 16970 4295 17016
rect 4363 16970 4409 17016
rect 4477 16970 4523 17016
rect 4591 16970 4637 17016
rect 4705 16970 4751 17016
rect 4819 16970 4865 17016
rect 4933 16970 4979 17016
rect 5047 16970 5093 17016
rect 5161 16970 5207 17016
rect 5275 16970 5321 17016
rect 5389 16970 5435 17016
rect 5503 16970 5549 17016
rect 5617 16970 5663 17016
rect 5731 16970 5777 17016
rect 5845 16970 5891 17016
rect 5959 16970 6005 17016
rect 6073 16970 6119 17016
rect 6187 16970 6233 17016
rect 6301 16970 6347 17016
rect 6415 16970 6461 17016
rect 6529 16970 6575 17016
rect 6643 16970 6689 17016
rect 6757 16970 6803 17016
rect 6871 16970 6917 17016
rect 6985 16970 7031 17016
rect 7099 16970 7145 17016
rect 7213 16970 7259 17016
rect 7327 16970 7373 17016
rect 7441 16970 7487 17016
rect 7555 16970 7601 17016
rect 7669 16970 7715 17016
rect 7783 16970 7829 17016
rect 7897 16970 7943 17016
rect 8011 16970 8057 17016
rect 8125 16970 8171 17016
rect 8239 16970 8285 17016
rect 8353 16970 8399 17016
rect 8467 16970 8513 17016
rect 8581 16970 8627 17016
rect 8695 16970 8741 17016
rect 8809 16970 8855 17016
rect 8923 16970 8969 17016
rect 9037 16970 9083 17016
rect 9151 16970 9197 17016
rect 9265 16970 9311 17016
rect 9379 16970 9425 17016
rect 9493 16970 9539 17016
rect 9607 16970 9653 17016
rect 9721 16970 9767 17016
rect 9835 16970 9881 17016
rect 9949 16970 9995 17016
rect 10063 16970 10109 17016
rect 10177 16970 10223 17016
rect 10291 16970 10337 17016
rect 10405 16970 10451 17016
rect 10519 16970 10565 17016
rect 10633 16970 10679 17016
rect 10747 16970 10793 17016
rect 10861 16970 10907 17016
rect 10975 16970 11021 17016
rect 11089 16970 11135 17016
rect 11203 16970 11249 17016
rect 11317 16970 11363 17016
rect 11431 16970 11477 17016
rect 11545 16970 11591 17016
rect 11659 16970 11705 17016
rect 11773 16970 11819 17016
rect 11927 16970 11973 17016
rect 12041 16970 12087 17016
rect 1587 16856 1633 16902
rect 1701 16856 1747 16902
rect 1855 16856 1901 16902
rect 1969 16856 2015 16902
rect 2083 16856 2129 16902
rect 2197 16856 2243 16902
rect 2311 16856 2357 16902
rect 2425 16856 2471 16902
rect 2539 16856 2585 16902
rect 2653 16856 2699 16902
rect 2767 16856 2813 16902
rect 2881 16856 2927 16902
rect 2995 16856 3041 16902
rect 3109 16856 3155 16902
rect 3223 16856 3269 16902
rect 3337 16856 3383 16902
rect 3451 16856 3497 16902
rect 3565 16856 3611 16902
rect 3679 16856 3725 16902
rect 3793 16856 3839 16902
rect 3907 16856 3953 16902
rect 4021 16856 4067 16902
rect 4135 16856 4181 16902
rect 4249 16856 4295 16902
rect 4363 16856 4409 16902
rect 4477 16856 4523 16902
rect 4591 16856 4637 16902
rect 4705 16856 4751 16902
rect 4819 16856 4865 16902
rect 4933 16856 4979 16902
rect 5047 16856 5093 16902
rect 5161 16856 5207 16902
rect 5275 16856 5321 16902
rect 5389 16856 5435 16902
rect 5503 16856 5549 16902
rect 5617 16856 5663 16902
rect 5731 16856 5777 16902
rect 5845 16856 5891 16902
rect 5959 16856 6005 16902
rect 6073 16856 6119 16902
rect 6187 16856 6233 16902
rect 6301 16856 6347 16902
rect 6415 16856 6461 16902
rect 6529 16856 6575 16902
rect 6643 16856 6689 16902
rect 6757 16856 6803 16902
rect 6871 16856 6917 16902
rect 6985 16856 7031 16902
rect 7099 16856 7145 16902
rect 7213 16856 7259 16902
rect 7327 16856 7373 16902
rect 7441 16856 7487 16902
rect 7555 16856 7601 16902
rect 7669 16856 7715 16902
rect 7783 16856 7829 16902
rect 7897 16856 7943 16902
rect 8011 16856 8057 16902
rect 8125 16856 8171 16902
rect 8239 16856 8285 16902
rect 8353 16856 8399 16902
rect 8467 16856 8513 16902
rect 8581 16856 8627 16902
rect 8695 16856 8741 16902
rect 8809 16856 8855 16902
rect 8923 16856 8969 16902
rect 9037 16856 9083 16902
rect 9151 16856 9197 16902
rect 9265 16856 9311 16902
rect 9379 16856 9425 16902
rect 9493 16856 9539 16902
rect 9607 16856 9653 16902
rect 9721 16856 9767 16902
rect 9835 16856 9881 16902
rect 9949 16856 9995 16902
rect 10063 16856 10109 16902
rect 10177 16856 10223 16902
rect 10291 16856 10337 16902
rect 10405 16856 10451 16902
rect 10519 16856 10565 16902
rect 10633 16856 10679 16902
rect 10747 16856 10793 16902
rect 10861 16856 10907 16902
rect 10975 16856 11021 16902
rect 11089 16856 11135 16902
rect 11203 16856 11249 16902
rect 11317 16856 11363 16902
rect 11431 16856 11477 16902
rect 11545 16856 11591 16902
rect 11659 16856 11705 16902
rect 11773 16856 11819 16902
rect 11927 16856 11973 16902
rect 12041 16856 12087 16902
rect 1587 16742 1633 16788
rect 1701 16742 1747 16788
rect 11927 16742 11973 16788
rect 12041 16742 12087 16788
rect 11927 16628 11973 16674
rect 12041 16628 12087 16674
rect 11927 16514 11973 16560
rect 12041 16514 12087 16560
rect 11927 16400 11973 16446
rect 12041 16400 12087 16446
rect 1587 16172 1633 16218
rect 1701 16172 1747 16218
rect 1587 16058 1633 16104
rect 1701 16058 1747 16104
rect 1587 15944 1633 15990
rect 1701 15944 1747 15990
rect 1587 15830 1633 15876
rect 1701 15830 1747 15876
rect 1587 15716 1633 15762
rect 1701 15716 1747 15762
rect 1587 15602 1633 15648
rect 1701 15602 1747 15648
rect 1587 15488 1633 15534
rect 1701 15488 1747 15534
rect 1587 15374 1633 15420
rect 1701 15374 1747 15420
rect 1587 15260 1633 15306
rect 1701 15260 1747 15306
rect 1587 15146 1633 15192
rect 1701 15146 1747 15192
rect 1587 15032 1633 15078
rect 1701 15032 1747 15078
rect 1587 14918 1633 14964
rect 1701 14918 1747 14964
rect 1587 14804 1633 14850
rect 1701 14804 1747 14850
rect 1587 14690 1633 14736
rect 1701 14690 1747 14736
rect 1587 14576 1633 14622
rect 1701 14576 1747 14622
rect 1587 14462 1633 14508
rect 1701 14462 1747 14508
rect 1587 14348 1633 14394
rect 1701 14348 1747 14394
rect 1587 14234 1633 14280
rect 1701 14234 1747 14280
rect 1587 14120 1633 14166
rect 1701 14120 1747 14166
rect 1587 14006 1633 14052
rect 1701 14006 1747 14052
rect 1587 13892 1633 13938
rect 1701 13892 1747 13938
rect 1587 13778 1633 13824
rect 1701 13778 1747 13824
rect 1587 13664 1633 13710
rect 1701 13664 1747 13710
rect 1587 13550 1633 13596
rect 1701 13550 1747 13596
rect 1587 13436 1633 13482
rect 1701 13436 1747 13482
rect 1587 13322 1633 13368
rect 1701 13322 1747 13368
rect 1587 13208 1633 13254
rect 1701 13208 1747 13254
rect 1587 13094 1633 13140
rect 1701 13094 1747 13140
rect 1587 12980 1633 13026
rect 1701 12980 1747 13026
rect 1587 12866 1633 12912
rect 1701 12866 1747 12912
rect 1587 12752 1633 12798
rect 1701 12752 1747 12798
rect 1587 12638 1633 12684
rect 1701 12638 1747 12684
rect 1587 12524 1633 12570
rect 1701 12524 1747 12570
rect 1587 12410 1633 12456
rect 1701 12410 1747 12456
rect 1587 12296 1633 12342
rect 1701 12296 1747 12342
rect 1587 12182 1633 12228
rect 1701 12182 1747 12228
rect 1587 12068 1633 12114
rect 1701 12068 1747 12114
rect 1587 11954 1633 12000
rect 1701 11954 1747 12000
rect 1587 11840 1633 11886
rect 1701 11840 1747 11886
rect 1587 11726 1633 11772
rect 1701 11726 1747 11772
rect 1587 11612 1633 11658
rect 1701 11612 1747 11658
rect 1587 11498 1633 11544
rect 1701 11498 1747 11544
rect 1587 11384 1633 11430
rect 1701 11384 1747 11430
rect 11927 16286 11973 16332
rect 12041 16286 12087 16332
rect 11927 16172 11973 16218
rect 12041 16172 12087 16218
rect 11927 16058 11973 16104
rect 12041 16058 12087 16104
rect 11927 15944 11973 15990
rect 12041 15944 12087 15990
rect 11927 15830 11973 15876
rect 12041 15830 12087 15876
rect 11927 15716 11973 15762
rect 12041 15716 12087 15762
rect 11927 15602 11973 15648
rect 12041 15602 12087 15648
rect 11927 15488 11973 15534
rect 12041 15488 12087 15534
rect 11927 15374 11973 15420
rect 12041 15374 12087 15420
rect 11927 15260 11973 15306
rect 12041 15260 12087 15306
rect 11927 15146 11973 15192
rect 12041 15146 12087 15192
rect 11927 15032 11973 15078
rect 12041 15032 12087 15078
rect 11927 14918 11973 14964
rect 12041 14918 12087 14964
rect 11927 14804 11973 14850
rect 12041 14804 12087 14850
rect 11927 14690 11973 14736
rect 12041 14690 12087 14736
rect 11927 14576 11973 14622
rect 12041 14576 12087 14622
rect 11927 14462 11973 14508
rect 12041 14462 12087 14508
rect 11927 14348 11973 14394
rect 12041 14348 12087 14394
rect 11927 14234 11973 14280
rect 12041 14234 12087 14280
rect 11927 14120 11973 14166
rect 12041 14120 12087 14166
rect 11927 14006 11973 14052
rect 12041 14006 12087 14052
rect 11927 13892 11973 13938
rect 12041 13892 12087 13938
rect 11927 13778 11973 13824
rect 12041 13778 12087 13824
rect 11927 13664 11973 13710
rect 12041 13664 12087 13710
rect 11927 13550 11973 13596
rect 12041 13550 12087 13596
rect 11927 13436 11973 13482
rect 12041 13436 12087 13482
rect 11927 13322 11973 13368
rect 12041 13322 12087 13368
rect 11927 13208 11973 13254
rect 12041 13208 12087 13254
rect 11927 13094 11973 13140
rect 12041 13094 12087 13140
rect 11927 12980 11973 13026
rect 12041 12980 12087 13026
rect 11927 12866 11973 12912
rect 12041 12866 12087 12912
rect 11927 12752 11973 12798
rect 12041 12752 12087 12798
rect 11927 12638 11973 12684
rect 12041 12638 12087 12684
rect 11927 12524 11973 12570
rect 12041 12524 12087 12570
rect 11927 12410 11973 12456
rect 12041 12410 12087 12456
rect 11927 12296 11973 12342
rect 12041 12296 12087 12342
rect 11927 12182 11973 12228
rect 12041 12182 12087 12228
rect 11927 12068 11973 12114
rect 12041 12068 12087 12114
rect 11927 11954 11973 12000
rect 12041 11954 12087 12000
rect 11927 11840 11973 11886
rect 12041 11840 12087 11886
rect 11927 11726 11973 11772
rect 12041 11726 12087 11772
rect 11927 11612 11973 11658
rect 12041 11612 12087 11658
rect 11927 11498 11973 11544
rect 12041 11498 12087 11544
rect 11927 11384 11973 11430
rect 12041 11384 12087 11430
rect 1587 11270 1633 11316
rect 1701 11270 1747 11316
rect 11927 11270 11973 11316
rect 12041 11270 12087 11316
rect 1587 11156 1633 11202
rect 1701 11156 1747 11202
rect 1587 11042 1633 11088
rect 1701 11042 1747 11088
rect 1587 10928 1633 10974
rect 1701 10928 1747 10974
rect 11927 11156 11973 11202
rect 12041 11156 12087 11202
rect 11927 11042 11973 11088
rect 12041 11042 12087 11088
rect 11927 10928 11973 10974
rect 12041 10928 12087 10974
rect 1855 10879 1901 10925
rect 1969 10879 2015 10925
rect 2083 10879 2129 10925
rect 2197 10879 2243 10925
rect 2311 10879 2357 10925
rect 2425 10879 2471 10925
rect 2539 10879 2585 10925
rect 2653 10879 2699 10925
rect 2767 10879 2813 10925
rect 2881 10879 2927 10925
rect 2995 10879 3041 10925
rect 3109 10879 3155 10925
rect 3223 10879 3269 10925
rect 3337 10879 3383 10925
rect 3451 10879 3497 10925
rect 3565 10879 3611 10925
rect 3679 10879 3725 10925
rect 3793 10879 3839 10925
rect 3907 10879 3953 10925
rect 4021 10879 4067 10925
rect 4135 10879 4181 10925
rect 4249 10879 4295 10925
rect 4363 10879 4409 10925
rect 4477 10879 4523 10925
rect 4591 10879 4637 10925
rect 4705 10879 4751 10925
rect 4819 10879 4865 10925
rect 4933 10879 4979 10925
rect 5047 10879 5093 10925
rect 5161 10879 5207 10925
rect 5275 10879 5321 10925
rect 5389 10879 5435 10925
rect 5503 10879 5549 10925
rect 5617 10879 5663 10925
rect 5731 10879 5777 10925
rect 5845 10879 5891 10925
rect 5959 10879 6005 10925
rect 6073 10879 6119 10925
rect 6187 10879 6233 10925
rect 6301 10879 6347 10925
rect 6415 10879 6461 10925
rect 6529 10879 6575 10925
rect 6643 10879 6689 10925
rect 6757 10879 6803 10925
rect 6871 10879 6917 10925
rect 6985 10879 7031 10925
rect 7099 10879 7145 10925
rect 7213 10879 7259 10925
rect 7327 10879 7373 10925
rect 7441 10879 7487 10925
rect 7555 10879 7601 10925
rect 7669 10879 7715 10925
rect 7783 10879 7829 10925
rect 7897 10879 7943 10925
rect 8011 10879 8057 10925
rect 8125 10879 8171 10925
rect 8239 10879 8285 10925
rect 8353 10879 8399 10925
rect 8467 10879 8513 10925
rect 8581 10879 8627 10925
rect 8695 10879 8741 10925
rect 8809 10879 8855 10925
rect 8923 10879 8969 10925
rect 9037 10879 9083 10925
rect 9151 10879 9197 10925
rect 9265 10879 9311 10925
rect 9379 10879 9425 10925
rect 9493 10879 9539 10925
rect 9607 10879 9653 10925
rect 9721 10879 9767 10925
rect 9835 10879 9881 10925
rect 9949 10879 9995 10925
rect 10063 10879 10109 10925
rect 10177 10879 10223 10925
rect 10291 10879 10337 10925
rect 10405 10879 10451 10925
rect 10519 10879 10565 10925
rect 10633 10879 10679 10925
rect 10747 10879 10793 10925
rect 10861 10879 10907 10925
rect 10975 10879 11021 10925
rect 11089 10879 11135 10925
rect 11203 10879 11249 10925
rect 11317 10879 11363 10925
rect 11431 10879 11477 10925
rect 11545 10879 11591 10925
rect 11659 10879 11705 10925
rect 11773 10879 11819 10925
rect 1587 10814 1633 10860
rect 1701 10814 1747 10860
rect 11927 10814 11973 10860
rect 12041 10814 12087 10860
rect 1855 10765 1901 10811
rect 1969 10765 2015 10811
rect 2083 10765 2129 10811
rect 2197 10765 2243 10811
rect 2311 10765 2357 10811
rect 2425 10765 2471 10811
rect 2539 10765 2585 10811
rect 2653 10765 2699 10811
rect 2767 10765 2813 10811
rect 2881 10765 2927 10811
rect 2995 10765 3041 10811
rect 3109 10765 3155 10811
rect 3223 10765 3269 10811
rect 3337 10765 3383 10811
rect 3451 10765 3497 10811
rect 3565 10765 3611 10811
rect 3679 10765 3725 10811
rect 3793 10765 3839 10811
rect 3907 10765 3953 10811
rect 4021 10765 4067 10811
rect 4135 10765 4181 10811
rect 4249 10765 4295 10811
rect 4363 10765 4409 10811
rect 4477 10765 4523 10811
rect 4591 10765 4637 10811
rect 4705 10765 4751 10811
rect 4819 10765 4865 10811
rect 4933 10765 4979 10811
rect 5047 10765 5093 10811
rect 5161 10765 5207 10811
rect 5275 10765 5321 10811
rect 5389 10765 5435 10811
rect 5503 10765 5549 10811
rect 5617 10765 5663 10811
rect 5731 10765 5777 10811
rect 5845 10765 5891 10811
rect 5959 10765 6005 10811
rect 6073 10765 6119 10811
rect 6187 10765 6233 10811
rect 6301 10765 6347 10811
rect 6415 10765 6461 10811
rect 6529 10765 6575 10811
rect 6643 10765 6689 10811
rect 6757 10765 6803 10811
rect 6871 10765 6917 10811
rect 6985 10765 7031 10811
rect 7099 10765 7145 10811
rect 7213 10765 7259 10811
rect 7327 10765 7373 10811
rect 7441 10765 7487 10811
rect 7555 10765 7601 10811
rect 7669 10765 7715 10811
rect 7783 10765 7829 10811
rect 7897 10765 7943 10811
rect 8011 10765 8057 10811
rect 8125 10765 8171 10811
rect 8239 10765 8285 10811
rect 8353 10765 8399 10811
rect 8467 10765 8513 10811
rect 8581 10765 8627 10811
rect 8695 10765 8741 10811
rect 8809 10765 8855 10811
rect 8923 10765 8969 10811
rect 9037 10765 9083 10811
rect 9151 10765 9197 10811
rect 9265 10765 9311 10811
rect 9379 10765 9425 10811
rect 9493 10765 9539 10811
rect 9607 10765 9653 10811
rect 9721 10765 9767 10811
rect 9835 10765 9881 10811
rect 9949 10765 9995 10811
rect 10063 10765 10109 10811
rect 10177 10765 10223 10811
rect 10291 10765 10337 10811
rect 10405 10765 10451 10811
rect 10519 10765 10565 10811
rect 10633 10765 10679 10811
rect 10747 10765 10793 10811
rect 10861 10765 10907 10811
rect 10975 10765 11021 10811
rect 11089 10765 11135 10811
rect 11203 10765 11249 10811
rect 11317 10765 11363 10811
rect 11431 10765 11477 10811
rect 11545 10765 11591 10811
rect 11659 10765 11705 10811
rect 11773 10765 11819 10811
rect 1587 10700 1633 10746
rect 1701 10700 1747 10746
rect 1587 10586 1633 10632
rect 1701 10586 1747 10632
rect 1587 10472 1633 10518
rect 1701 10472 1747 10518
rect 11927 10700 11973 10746
rect 12041 10700 12087 10746
rect 11927 10586 11973 10632
rect 12041 10586 12087 10632
rect 11927 10472 11973 10518
rect 12041 10472 12087 10518
rect 1587 10358 1633 10404
rect 1701 10358 1747 10404
rect 11927 10358 11973 10404
rect 12041 10358 12087 10404
rect 1587 10244 1633 10290
rect 1701 10244 1747 10290
rect 1587 10130 1633 10176
rect 1701 10130 1747 10176
rect 1587 10016 1633 10062
rect 1701 10016 1747 10062
rect 1587 9902 1633 9948
rect 1701 9902 1747 9948
rect 1587 9788 1633 9834
rect 1701 9788 1747 9834
rect 1587 9674 1633 9720
rect 1701 9674 1747 9720
rect 1587 9560 1633 9606
rect 1701 9560 1747 9606
rect 1587 9446 1633 9492
rect 1701 9446 1747 9492
rect 1587 9332 1633 9378
rect 1701 9332 1747 9378
rect 1587 9218 1633 9264
rect 1701 9218 1747 9264
rect 1587 9104 1633 9150
rect 1701 9104 1747 9150
rect 1587 8990 1633 9036
rect 1701 8990 1747 9036
rect 1587 8876 1633 8922
rect 1701 8876 1747 8922
rect 1587 8762 1633 8808
rect 1701 8762 1747 8808
rect 1587 8648 1633 8694
rect 1701 8648 1747 8694
rect 1587 8534 1633 8580
rect 1701 8534 1747 8580
rect 1587 8420 1633 8466
rect 1701 8420 1747 8466
rect 1587 8306 1633 8352
rect 1701 8306 1747 8352
rect 1587 8192 1633 8238
rect 1701 8192 1747 8238
rect 1587 8078 1633 8124
rect 1701 8078 1747 8124
rect 1587 7964 1633 8010
rect 1701 7964 1747 8010
rect 1587 7850 1633 7896
rect 1701 7850 1747 7896
rect 1587 7736 1633 7782
rect 1701 7736 1747 7782
rect 1587 7622 1633 7668
rect 1701 7622 1747 7668
rect 1587 7508 1633 7554
rect 1701 7508 1747 7554
rect 1587 7394 1633 7440
rect 1701 7394 1747 7440
rect 1587 7280 1633 7326
rect 1701 7280 1747 7326
rect 1587 7166 1633 7212
rect 1701 7166 1747 7212
rect 1587 7052 1633 7098
rect 1701 7052 1747 7098
rect 1587 6938 1633 6984
rect 1701 6938 1747 6984
rect 1587 6824 1633 6870
rect 1701 6824 1747 6870
rect 1587 6710 1633 6756
rect 1701 6710 1747 6756
rect 1587 6596 1633 6642
rect 1701 6596 1747 6642
rect 1587 6482 1633 6528
rect 1701 6482 1747 6528
rect 1587 6368 1633 6414
rect 1701 6368 1747 6414
rect 1587 6254 1633 6300
rect 1701 6254 1747 6300
rect 1587 6140 1633 6186
rect 1701 6140 1747 6186
rect 1587 6026 1633 6072
rect 1701 6026 1747 6072
rect 1587 5912 1633 5958
rect 1701 5912 1747 5958
rect 1587 5798 1633 5844
rect 1701 5798 1747 5844
rect 1587 5684 1633 5730
rect 1701 5684 1747 5730
rect 1587 5570 1633 5616
rect 1701 5570 1747 5616
rect 1587 5456 1633 5502
rect 1701 5456 1747 5502
rect 11927 10244 11973 10290
rect 12041 10244 12087 10290
rect 11927 10130 11973 10176
rect 12041 10130 12087 10176
rect 11927 10016 11973 10062
rect 12041 10016 12087 10062
rect 11927 9902 11973 9948
rect 12041 9902 12087 9948
rect 11927 9788 11973 9834
rect 12041 9788 12087 9834
rect 11927 9674 11973 9720
rect 12041 9674 12087 9720
rect 11927 9560 11973 9606
rect 12041 9560 12087 9606
rect 11927 9446 11973 9492
rect 12041 9446 12087 9492
rect 11927 9332 11973 9378
rect 12041 9332 12087 9378
rect 11927 9218 11973 9264
rect 12041 9218 12087 9264
rect 11927 9104 11973 9150
rect 12041 9104 12087 9150
rect 11927 8990 11973 9036
rect 12041 8990 12087 9036
rect 11927 8876 11973 8922
rect 12041 8876 12087 8922
rect 11927 8762 11973 8808
rect 12041 8762 12087 8808
rect 11927 8648 11973 8694
rect 12041 8648 12087 8694
rect 11927 8534 11973 8580
rect 12041 8534 12087 8580
rect 11927 8420 11973 8466
rect 12041 8420 12087 8466
rect 11927 8306 11973 8352
rect 12041 8306 12087 8352
rect 11927 8192 11973 8238
rect 12041 8192 12087 8238
rect 11927 8078 11973 8124
rect 12041 8078 12087 8124
rect 11927 7964 11973 8010
rect 12041 7964 12087 8010
rect 11927 7850 11973 7896
rect 12041 7850 12087 7896
rect 11927 7736 11973 7782
rect 12041 7736 12087 7782
rect 11927 7622 11973 7668
rect 12041 7622 12087 7668
rect 11927 7508 11973 7554
rect 12041 7508 12087 7554
rect 11927 7394 11973 7440
rect 12041 7394 12087 7440
rect 11927 7280 11973 7326
rect 12041 7280 12087 7326
rect 11927 7166 11973 7212
rect 12041 7166 12087 7212
rect 11927 7052 11973 7098
rect 12041 7052 12087 7098
rect 11927 6938 11973 6984
rect 12041 6938 12087 6984
rect 11927 6824 11973 6870
rect 12041 6824 12087 6870
rect 11927 6710 11973 6756
rect 12041 6710 12087 6756
rect 11927 6596 11973 6642
rect 12041 6596 12087 6642
rect 11927 6482 11973 6528
rect 12041 6482 12087 6528
rect 11927 6368 11973 6414
rect 12041 6368 12087 6414
rect 11927 6254 11973 6300
rect 12041 6254 12087 6300
rect 11927 6140 11973 6186
rect 12041 6140 12087 6186
rect 11927 6026 11973 6072
rect 12041 6026 12087 6072
rect 11927 5912 11973 5958
rect 12041 5912 12087 5958
rect 11927 5798 11973 5844
rect 12041 5798 12087 5844
rect 11927 5684 11973 5730
rect 12041 5684 12087 5730
rect 11927 5570 11973 5616
rect 12041 5570 12087 5616
rect 11927 5456 11973 5502
rect 12041 5456 12087 5502
rect 11927 5342 11973 5388
rect 12041 5342 12087 5388
rect 1587 5000 1633 5046
rect 1701 5000 1747 5046
rect 11927 5228 11973 5274
rect 12041 5228 12087 5274
rect 11927 5114 11973 5160
rect 12041 5114 12087 5160
rect 11927 5000 11973 5046
rect 12041 5000 12087 5046
rect 1587 4886 1633 4932
rect 1701 4886 1747 4932
rect 1855 4886 1901 4932
rect 1969 4886 2015 4932
rect 2083 4886 2129 4932
rect 2197 4886 2243 4932
rect 2311 4886 2357 4932
rect 2425 4886 2471 4932
rect 2539 4886 2585 4932
rect 2653 4886 2699 4932
rect 2767 4886 2813 4932
rect 2881 4886 2927 4932
rect 2995 4886 3041 4932
rect 3109 4886 3155 4932
rect 3223 4886 3269 4932
rect 3337 4886 3383 4932
rect 3451 4886 3497 4932
rect 3565 4886 3611 4932
rect 3679 4886 3725 4932
rect 3793 4886 3839 4932
rect 3907 4886 3953 4932
rect 4021 4886 4067 4932
rect 4135 4886 4181 4932
rect 4249 4886 4295 4932
rect 4363 4886 4409 4932
rect 4477 4886 4523 4932
rect 4591 4886 4637 4932
rect 4705 4886 4751 4932
rect 4819 4886 4865 4932
rect 4933 4886 4979 4932
rect 5047 4886 5093 4932
rect 5161 4886 5207 4932
rect 5275 4886 5321 4932
rect 5389 4886 5435 4932
rect 5503 4886 5549 4932
rect 5617 4886 5663 4932
rect 5731 4886 5777 4932
rect 5845 4886 5891 4932
rect 5959 4886 6005 4932
rect 6073 4886 6119 4932
rect 6187 4886 6233 4932
rect 6301 4886 6347 4932
rect 6415 4886 6461 4932
rect 6529 4886 6575 4932
rect 6643 4886 6689 4932
rect 6757 4886 6803 4932
rect 6871 4886 6917 4932
rect 6985 4886 7031 4932
rect 7099 4886 7145 4932
rect 7213 4886 7259 4932
rect 7327 4886 7373 4932
rect 7441 4886 7487 4932
rect 7555 4886 7601 4932
rect 7669 4886 7715 4932
rect 7783 4886 7829 4932
rect 7897 4886 7943 4932
rect 8011 4886 8057 4932
rect 8125 4886 8171 4932
rect 8239 4886 8285 4932
rect 8353 4886 8399 4932
rect 8467 4886 8513 4932
rect 8581 4886 8627 4932
rect 8695 4886 8741 4932
rect 8809 4886 8855 4932
rect 8923 4886 8969 4932
rect 9037 4886 9083 4932
rect 9151 4886 9197 4932
rect 9265 4886 9311 4932
rect 9379 4886 9425 4932
rect 9493 4886 9539 4932
rect 9607 4886 9653 4932
rect 9721 4886 9767 4932
rect 9835 4886 9881 4932
rect 9949 4886 9995 4932
rect 10063 4886 10109 4932
rect 10177 4886 10223 4932
rect 10291 4886 10337 4932
rect 10405 4886 10451 4932
rect 10519 4886 10565 4932
rect 10633 4886 10679 4932
rect 10747 4886 10793 4932
rect 10861 4886 10907 4932
rect 10975 4886 11021 4932
rect 11089 4886 11135 4932
rect 11203 4886 11249 4932
rect 11317 4886 11363 4932
rect 11431 4886 11477 4932
rect 11545 4886 11591 4932
rect 11659 4886 11705 4932
rect 11773 4886 11819 4932
rect 11927 4886 11973 4932
rect 12041 4886 12087 4932
rect 1587 4772 1633 4818
rect 1701 4772 1747 4818
rect 1855 4772 1901 4818
rect 1969 4772 2015 4818
rect 2083 4772 2129 4818
rect 2197 4772 2243 4818
rect 2311 4772 2357 4818
rect 2425 4772 2471 4818
rect 2539 4772 2585 4818
rect 2653 4772 2699 4818
rect 2767 4772 2813 4818
rect 2881 4772 2927 4818
rect 2995 4772 3041 4818
rect 3109 4772 3155 4818
rect 3223 4772 3269 4818
rect 3337 4772 3383 4818
rect 3451 4772 3497 4818
rect 3565 4772 3611 4818
rect 3679 4772 3725 4818
rect 3793 4772 3839 4818
rect 3907 4772 3953 4818
rect 4021 4772 4067 4818
rect 4135 4772 4181 4818
rect 4249 4772 4295 4818
rect 4363 4772 4409 4818
rect 4477 4772 4523 4818
rect 4591 4772 4637 4818
rect 4705 4772 4751 4818
rect 4819 4772 4865 4818
rect 4933 4772 4979 4818
rect 5047 4772 5093 4818
rect 5161 4772 5207 4818
rect 5275 4772 5321 4818
rect 5389 4772 5435 4818
rect 5503 4772 5549 4818
rect 5617 4772 5663 4818
rect 5731 4772 5777 4818
rect 5845 4772 5891 4818
rect 5959 4772 6005 4818
rect 6073 4772 6119 4818
rect 6187 4772 6233 4818
rect 6301 4772 6347 4818
rect 6415 4772 6461 4818
rect 6529 4772 6575 4818
rect 6643 4772 6689 4818
rect 6757 4772 6803 4818
rect 6871 4772 6917 4818
rect 6985 4772 7031 4818
rect 7099 4772 7145 4818
rect 7213 4772 7259 4818
rect 7327 4772 7373 4818
rect 7441 4772 7487 4818
rect 7555 4772 7601 4818
rect 7669 4772 7715 4818
rect 7783 4772 7829 4818
rect 7897 4772 7943 4818
rect 8011 4772 8057 4818
rect 8125 4772 8171 4818
rect 8239 4772 8285 4818
rect 8353 4772 8399 4818
rect 8467 4772 8513 4818
rect 8581 4772 8627 4818
rect 8695 4772 8741 4818
rect 8809 4772 8855 4818
rect 8923 4772 8969 4818
rect 9037 4772 9083 4818
rect 9151 4772 9197 4818
rect 9265 4772 9311 4818
rect 9379 4772 9425 4818
rect 9493 4772 9539 4818
rect 9607 4772 9653 4818
rect 9721 4772 9767 4818
rect 9835 4772 9881 4818
rect 9949 4772 9995 4818
rect 10063 4772 10109 4818
rect 10177 4772 10223 4818
rect 10291 4772 10337 4818
rect 10405 4772 10451 4818
rect 10519 4772 10565 4818
rect 10633 4772 10679 4818
rect 10747 4772 10793 4818
rect 10861 4772 10907 4818
rect 10975 4772 11021 4818
rect 11089 4772 11135 4818
rect 11203 4772 11249 4818
rect 11317 4772 11363 4818
rect 11431 4772 11477 4818
rect 11545 4772 11591 4818
rect 11659 4772 11705 4818
rect 11773 4772 11819 4818
rect 11927 4772 11973 4818
rect 12041 4772 12087 4818
<< nsubdiffcont >>
rect 54 4336 100 4382
rect 158 4336 204 4382
rect 574 4336 620 4382
rect 678 4336 724 4382
rect 782 4336 828 4382
rect 886 4336 932 4382
rect 990 4336 1036 4382
rect 1094 4336 1140 4382
rect 1198 4336 1244 4382
rect 1302 4336 1348 4382
rect 1406 4336 1452 4382
rect 1510 4336 1556 4382
rect 1614 4336 1660 4382
rect 1718 4336 1764 4382
rect 1822 4336 1868 4382
rect 1926 4336 1972 4382
rect 2030 4336 2076 4382
rect 2134 4336 2180 4382
rect 2238 4336 2284 4382
rect 2342 4336 2388 4382
rect 2446 4336 2492 4382
rect 2550 4336 2596 4382
rect 2654 4336 2700 4382
rect 2758 4336 2804 4382
rect 2862 4336 2908 4382
rect 2966 4336 3012 4382
rect 3070 4336 3116 4382
rect 3174 4336 3220 4382
rect 3278 4336 3324 4382
rect 3382 4336 3428 4382
rect 3486 4336 3532 4382
rect 3590 4336 3636 4382
rect 3694 4336 3740 4382
rect 3798 4336 3844 4382
rect 3902 4336 3948 4382
rect 4006 4336 4052 4382
rect 4110 4336 4156 4382
rect 4214 4336 4260 4382
rect 4318 4336 4364 4382
rect 4422 4336 4468 4382
rect 4526 4336 4572 4382
rect 4630 4336 4676 4382
rect 4734 4336 4780 4382
rect 4838 4336 4884 4382
rect 4942 4336 4988 4382
rect 5046 4336 5092 4382
rect 5150 4336 5196 4382
rect 5254 4336 5300 4382
rect 5358 4336 5404 4382
rect 5462 4336 5508 4382
rect 5566 4336 5612 4382
rect 5670 4336 5716 4382
rect 5774 4336 5820 4382
rect 5878 4336 5924 4382
rect 5982 4336 6028 4382
rect 6086 4336 6132 4382
rect 6190 4336 6236 4382
rect 6294 4336 6340 4382
rect 6398 4336 6444 4382
rect 6502 4336 6548 4382
rect 6606 4336 6652 4382
rect 6710 4336 6756 4382
rect 6814 4336 6860 4382
rect 6918 4336 6964 4382
rect 7022 4336 7068 4382
rect 7126 4336 7172 4382
rect 7230 4336 7276 4382
rect 7334 4336 7380 4382
rect 7438 4336 7484 4382
rect 7542 4336 7588 4382
rect 7646 4336 7692 4382
rect 7750 4336 7796 4382
rect 7854 4336 7900 4382
rect 7958 4336 8004 4382
rect 8062 4336 8108 4382
rect 8166 4336 8212 4382
rect 8270 4336 8316 4382
rect 8374 4336 8420 4382
rect 8478 4336 8524 4382
rect 8582 4336 8628 4382
rect 8686 4336 8732 4382
rect 8790 4336 8836 4382
rect 8894 4336 8940 4382
rect 8998 4336 9044 4382
rect 9102 4336 9148 4382
rect 9206 4336 9252 4382
rect 9310 4336 9356 4382
rect 9414 4336 9460 4382
rect 9518 4336 9564 4382
rect 9622 4336 9668 4382
rect 9726 4336 9772 4382
rect 9830 4336 9876 4382
rect 9934 4336 9980 4382
rect 10038 4336 10084 4382
rect 10142 4336 10188 4382
rect 10246 4336 10292 4382
rect 10350 4336 10396 4382
rect 10454 4336 10500 4382
rect 10558 4336 10604 4382
rect 10662 4336 10708 4382
rect 10766 4336 10812 4382
rect 10870 4336 10916 4382
rect 10974 4336 11020 4382
rect 11078 4336 11124 4382
rect 11182 4336 11228 4382
rect 11286 4336 11332 4382
rect 11390 4336 11436 4382
rect 11494 4336 11540 4382
rect 11598 4336 11644 4382
rect 11702 4336 11748 4382
rect 11806 4336 11852 4382
rect 11910 4336 11956 4382
rect 12014 4336 12060 4382
rect 12118 4336 12164 4382
rect 12222 4336 12268 4382
rect 12326 4336 12372 4382
rect 12430 4336 12476 4382
rect 12534 4336 12580 4382
rect 12638 4336 12684 4382
rect 12742 4336 12788 4382
rect 12846 4336 12892 4382
rect 12950 4336 12996 4382
rect 13054 4336 13100 4382
rect 13158 4336 13204 4382
rect 13262 4336 13308 4382
rect 13366 4336 13412 4382
rect 13470 4336 13516 4382
rect 13574 4336 13620 4382
rect 54 4182 100 4228
rect 54 4078 100 4124
rect 13574 4182 13620 4228
rect 54 3974 100 4020
rect 13574 4078 13620 4124
rect 13574 3974 13620 4020
rect 54 3870 100 3916
rect 13574 3870 13620 3916
rect 54 3766 100 3812
rect 54 3662 100 3708
rect 13574 3766 13620 3812
rect 54 3558 100 3604
rect 13574 3662 13620 3708
rect 13574 3558 13620 3604
rect 54 3454 100 3500
rect 54 3350 100 3396
rect 13574 3454 13620 3500
rect 54 3246 100 3292
rect 13574 3350 13620 3396
rect 54 3142 100 3188
rect 13574 3246 13620 3292
rect 13574 3142 13620 3188
rect 54 3038 100 3084
rect 13574 3038 13620 3084
rect 54 2934 100 2980
rect 54 2830 100 2876
rect 13574 2934 13620 2980
rect 13574 2830 13620 2876
rect 54 2726 100 2772
rect 13574 2726 13620 2772
rect 54 2622 100 2668
rect 54 2518 100 2564
rect 13574 2622 13620 2668
rect 54 2414 100 2460
rect 13574 2518 13620 2564
rect 54 2310 100 2356
rect 13574 2414 13620 2460
rect 13574 2310 13620 2356
rect 54 2206 100 2252
rect 13574 2206 13620 2252
rect 54 2102 100 2148
rect 54 1998 100 2044
rect 13574 2102 13620 2148
rect 13574 1998 13620 2044
rect 54 1894 100 1940
rect 13574 1894 13620 1940
rect 54 1790 100 1836
rect 54 1686 100 1732
rect 13574 1790 13620 1836
rect 54 1582 100 1628
rect 13574 1686 13620 1732
rect 54 1478 100 1524
rect 13574 1582 13620 1628
rect 13574 1478 13620 1524
rect 54 1374 100 1420
rect 54 1270 100 1316
rect 13574 1374 13620 1420
rect 54 1166 100 1212
rect 13574 1270 13620 1316
rect 13574 1166 13620 1212
rect 54 1062 100 1108
rect 13574 1062 13620 1108
rect 54 958 100 1004
rect 54 854 100 900
rect 13574 958 13620 1004
rect 54 750 100 796
rect 13574 854 13620 900
rect 13574 750 13620 796
rect 54 596 100 642
rect 158 596 204 642
rect 262 596 308 642
rect 366 596 412 642
rect 470 596 516 642
rect 574 596 620 642
rect 678 596 724 642
rect 782 596 828 642
rect 886 596 932 642
rect 990 596 1036 642
rect 1094 596 1140 642
rect 1198 596 1244 642
rect 1302 596 1348 642
rect 1406 596 1452 642
rect 1510 596 1556 642
rect 1614 596 1660 642
rect 1718 596 1764 642
rect 1822 596 1868 642
rect 1926 596 1972 642
rect 2030 596 2076 642
rect 2134 596 2180 642
rect 2238 596 2284 642
rect 2342 596 2388 642
rect 2446 596 2492 642
rect 2550 596 2596 642
rect 2654 596 2700 642
rect 2758 596 2804 642
rect 2862 596 2908 642
rect 2966 596 3012 642
rect 3070 596 3116 642
rect 3174 596 3220 642
rect 3278 596 3324 642
rect 3382 596 3428 642
rect 3486 596 3532 642
rect 3590 596 3636 642
rect 3694 596 3740 642
rect 3798 596 3844 642
rect 3902 596 3948 642
rect 4006 596 4052 642
rect 4110 596 4156 642
rect 4214 596 4260 642
rect 4318 596 4364 642
rect 4422 596 4468 642
rect 4526 596 4572 642
rect 4630 596 4676 642
rect 4734 596 4780 642
rect 4838 596 4884 642
rect 4942 596 4988 642
rect 5046 596 5092 642
rect 5150 596 5196 642
rect 5254 596 5300 642
rect 5358 596 5404 642
rect 5462 596 5508 642
rect 5566 596 5612 642
rect 5670 596 5716 642
rect 5774 596 5820 642
rect 5878 596 5924 642
rect 5982 596 6028 642
rect 6086 596 6132 642
rect 6190 596 6236 642
rect 6294 596 6340 642
rect 6398 596 6444 642
rect 6502 596 6548 642
rect 6606 596 6652 642
rect 6710 596 6756 642
rect 6814 596 6860 642
rect 6918 596 6964 642
rect 7022 596 7068 642
rect 7126 596 7172 642
rect 7230 596 7276 642
rect 7334 596 7380 642
rect 7438 596 7484 642
rect 7542 596 7588 642
rect 7646 596 7692 642
rect 7750 596 7796 642
rect 7854 596 7900 642
rect 7958 596 8004 642
rect 8062 596 8108 642
rect 8166 596 8212 642
rect 8270 596 8316 642
rect 8374 596 8420 642
rect 8478 596 8524 642
rect 8582 596 8628 642
rect 8686 596 8732 642
rect 8790 596 8836 642
rect 8894 596 8940 642
rect 8998 596 9044 642
rect 9102 596 9148 642
rect 9206 596 9252 642
rect 9310 596 9356 642
rect 9414 596 9460 642
rect 9518 596 9564 642
rect 9622 596 9668 642
rect 9726 596 9772 642
rect 9830 596 9876 642
rect 9934 596 9980 642
rect 10038 596 10084 642
rect 10142 596 10188 642
rect 10246 596 10292 642
rect 10350 596 10396 642
rect 10454 596 10500 642
rect 10558 596 10604 642
rect 10662 596 10708 642
rect 10766 596 10812 642
rect 10870 596 10916 642
rect 10974 596 11020 642
rect 11078 596 11124 642
rect 11182 596 11228 642
rect 11286 596 11332 642
rect 11390 596 11436 642
rect 11494 596 11540 642
rect 11598 596 11644 642
rect 11702 596 11748 642
rect 11806 596 11852 642
rect 11910 596 11956 642
rect 12014 596 12060 642
rect 12118 596 12164 642
rect 12222 596 12268 642
rect 12326 596 12372 642
rect 12430 596 12476 642
rect 12534 596 12580 642
rect 12638 596 12684 642
rect 12742 596 12788 642
rect 12846 596 12892 642
rect 12950 596 12996 642
rect 13054 596 13100 642
rect 13158 596 13204 642
rect 13262 596 13308 642
rect 13366 596 13412 642
rect 13470 596 13516 642
rect 13574 596 13620 642
<< mvnmoscap >>
rect 2180 11351 4180 16351
rect 4616 11351 6616 16351
rect 7052 11351 9052 16351
rect 9488 11351 11488 16351
rect 2180 5339 4180 10339
rect 4616 5339 6616 10339
rect 7052 5339 9052 10339
rect 9488 5339 11488 10339
<< polysilicon >>
rect 2180 16430 4180 16443
rect 2180 16384 2233 16430
rect 4127 16384 4180 16430
rect 2180 16351 4180 16384
rect 4616 16430 6616 16443
rect 4616 16384 4669 16430
rect 6563 16384 6616 16430
rect 4616 16351 6616 16384
rect 7052 16430 9052 16443
rect 7052 16384 7105 16430
rect 8999 16384 9052 16430
rect 7052 16351 9052 16384
rect 9488 16430 11488 16443
rect 9488 16384 9541 16430
rect 11435 16384 11488 16430
rect 9488 16351 11488 16384
rect 2180 11318 4180 11351
rect 2180 11272 2233 11318
rect 4127 11272 4180 11318
rect 2180 11259 4180 11272
rect 4616 11318 6616 11351
rect 4616 11272 4669 11318
rect 6563 11272 6616 11318
rect 4616 11259 6616 11272
rect 7052 11318 9052 11351
rect 7052 11272 7105 11318
rect 8999 11272 9052 11318
rect 7052 11259 9052 11272
rect 9488 11318 11488 11351
rect 9488 11272 9541 11318
rect 11435 11272 11488 11318
rect 9488 11259 11488 11272
rect 2180 10418 4180 10431
rect 2180 10372 2233 10418
rect 4127 10372 4180 10418
rect 2180 10339 4180 10372
rect 4616 10418 6616 10431
rect 4616 10372 4669 10418
rect 6563 10372 6616 10418
rect 4616 10339 6616 10372
rect 7052 10418 9052 10431
rect 7052 10372 7105 10418
rect 8999 10372 9052 10418
rect 7052 10339 9052 10372
rect 9488 10418 11488 10431
rect 9488 10372 9541 10418
rect 11435 10372 11488 10418
rect 9488 10339 11488 10372
rect 2180 5306 4180 5339
rect 2180 5260 2233 5306
rect 4127 5260 4180 5306
rect 2180 5247 4180 5260
rect 4616 5306 6616 5339
rect 4616 5260 4669 5306
rect 6563 5260 6616 5306
rect 4616 5247 6616 5260
rect 7052 5306 9052 5339
rect 7052 5260 7105 5306
rect 8999 5260 9052 5306
rect 7052 5247 9052 5260
rect 9488 5306 11488 5339
rect 9488 5260 9541 5306
rect 11435 5260 11488 5306
rect 9488 5247 11488 5260
rect 353 4052 455 4109
rect 353 4006 366 4052
rect 412 4006 455 4052
rect 353 3949 455 4006
rect 13226 4052 13328 4109
rect 13226 4006 13269 4052
rect 13315 4006 13328 4052
rect 13226 3949 13328 4006
rect 353 3772 455 3829
rect 353 3726 366 3772
rect 412 3726 455 3772
rect 353 3669 455 3726
rect 13226 3772 13328 3829
rect 13226 3726 13269 3772
rect 13315 3726 13328 3772
rect 13226 3669 13328 3726
rect 353 3492 455 3549
rect 353 3446 366 3492
rect 412 3446 455 3492
rect 353 3389 455 3446
rect 13226 3492 13328 3549
rect 13226 3446 13269 3492
rect 13315 3446 13328 3492
rect 13226 3389 13328 3446
rect 353 3212 455 3269
rect 353 3166 366 3212
rect 412 3166 455 3212
rect 353 3109 455 3166
rect 13226 3212 13328 3269
rect 13226 3166 13269 3212
rect 13315 3166 13328 3212
rect 13226 3109 13328 3166
rect 353 2932 455 2989
rect 353 2886 366 2932
rect 412 2886 455 2932
rect 353 2829 455 2886
rect 13226 2932 13328 2989
rect 13226 2886 13269 2932
rect 13315 2886 13328 2932
rect 13226 2829 13328 2886
rect 353 2652 455 2709
rect 353 2606 366 2652
rect 412 2606 455 2652
rect 353 2549 455 2606
rect 13226 2652 13328 2709
rect 13226 2606 13269 2652
rect 13315 2606 13328 2652
rect 13226 2549 13328 2606
rect 353 2372 455 2429
rect 353 2326 366 2372
rect 412 2326 455 2372
rect 353 2269 455 2326
rect 13226 2372 13328 2429
rect 13226 2326 13269 2372
rect 13315 2326 13328 2372
rect 13226 2269 13328 2326
rect 353 2092 455 2149
rect 353 2046 366 2092
rect 412 2046 455 2092
rect 353 1989 455 2046
rect 13226 2092 13328 2149
rect 13226 2046 13269 2092
rect 13315 2046 13328 2092
rect 13226 1989 13328 2046
rect 353 1812 455 1869
rect 353 1766 366 1812
rect 412 1766 455 1812
rect 353 1709 455 1766
rect 13226 1812 13328 1869
rect 13226 1766 13269 1812
rect 13315 1766 13328 1812
rect 13226 1709 13328 1766
rect 353 1532 455 1589
rect 353 1486 366 1532
rect 412 1486 455 1532
rect 353 1429 455 1486
rect 13226 1532 13328 1589
rect 13226 1486 13269 1532
rect 13315 1486 13328 1532
rect 13226 1429 13328 1486
rect 353 1252 455 1309
rect 353 1206 366 1252
rect 412 1206 455 1252
rect 353 1149 455 1206
rect 13226 1252 13328 1309
rect 13226 1206 13269 1252
rect 13315 1206 13328 1252
rect 13226 1149 13328 1206
rect 353 972 455 1029
rect 353 926 366 972
rect 412 926 455 972
rect 353 869 455 926
rect 13226 972 13328 1029
rect 13226 926 13269 972
rect 13315 926 13328 972
rect 13226 869 13328 926
<< polycontact >>
rect 2233 16384 4127 16430
rect 4669 16384 6563 16430
rect 7105 16384 8999 16430
rect 9541 16384 11435 16430
rect 2233 11272 4127 11318
rect 4669 11272 6563 11318
rect 7105 11272 8999 11318
rect 9541 11272 11435 11318
rect 2233 10372 4127 10418
rect 4669 10372 6563 10418
rect 7105 10372 8999 10418
rect 9541 10372 11435 10418
rect 2233 5260 4127 5306
rect 4669 5260 6563 5306
rect 7105 5260 8999 5306
rect 9541 5260 11435 5306
rect 366 4006 412 4052
rect 13269 4006 13315 4052
rect 366 3726 412 3772
rect 13269 3726 13315 3772
rect 366 3446 412 3492
rect 13269 3446 13315 3492
rect 366 3166 412 3212
rect 13269 3166 13315 3212
rect 366 2886 412 2932
rect 13269 2886 13315 2932
rect 366 2606 412 2652
rect 13269 2606 13315 2652
rect 366 2326 412 2372
rect 13269 2326 13315 2372
rect 366 2046 412 2092
rect 13269 2046 13315 2092
rect 366 1766 412 1812
rect 13269 1766 13315 1812
rect 366 1486 412 1532
rect 13269 1486 13315 1532
rect 366 1206 412 1252
rect 13269 1206 13315 1252
rect 366 926 412 972
rect 13269 926 13315 972
<< ppolyres >>
rect 455 3949 13226 4109
rect 455 3669 13226 3829
rect 455 3389 13226 3549
rect 455 3109 13226 3269
rect 455 2829 13226 2989
rect 455 2549 13226 2709
rect 455 2269 13226 2429
rect 455 1989 13226 2149
rect 455 1709 13226 1869
rect 455 1429 13226 1589
rect 455 1149 13226 1309
rect 455 869 13226 1029
<< metal1 >>
rect 1576 17016 12098 17028
rect 1576 16970 1587 17016
rect 1633 16970 1701 17016
rect 1747 16970 1855 17016
rect 1901 16970 1969 17016
rect 2015 16970 2083 17016
rect 2129 16970 2197 17016
rect 2243 16970 2311 17016
rect 2357 16970 2425 17016
rect 2471 16970 2539 17016
rect 2585 16970 2653 17016
rect 2699 16970 2767 17016
rect 2813 16970 2881 17016
rect 2927 16970 2995 17016
rect 3041 16970 3109 17016
rect 3155 16970 3223 17016
rect 3269 16970 3337 17016
rect 3383 16970 3451 17016
rect 3497 16970 3565 17016
rect 3611 16970 3679 17016
rect 3725 16970 3793 17016
rect 3839 16970 3907 17016
rect 3953 16970 4021 17016
rect 4067 16970 4135 17016
rect 4181 16970 4249 17016
rect 4295 16970 4363 17016
rect 4409 16970 4477 17016
rect 4523 16970 4591 17016
rect 4637 16970 4705 17016
rect 4751 16970 4819 17016
rect 4865 16970 4933 17016
rect 4979 16970 5047 17016
rect 5093 16970 5161 17016
rect 5207 16970 5275 17016
rect 5321 16970 5389 17016
rect 5435 16970 5503 17016
rect 5549 16970 5617 17016
rect 5663 16970 5731 17016
rect 5777 16970 5845 17016
rect 5891 16970 5959 17016
rect 6005 16970 6073 17016
rect 6119 16970 6187 17016
rect 6233 16970 6301 17016
rect 6347 16970 6415 17016
rect 6461 16970 6529 17016
rect 6575 16970 6643 17016
rect 6689 16970 6757 17016
rect 6803 16970 6871 17016
rect 6917 16970 6985 17016
rect 7031 16970 7099 17016
rect 7145 16970 7213 17016
rect 7259 16970 7327 17016
rect 7373 16970 7441 17016
rect 7487 16970 7555 17016
rect 7601 16970 7669 17016
rect 7715 16970 7783 17016
rect 7829 16970 7897 17016
rect 7943 16970 8011 17016
rect 8057 16970 8125 17016
rect 8171 16970 8239 17016
rect 8285 16970 8353 17016
rect 8399 16970 8467 17016
rect 8513 16970 8581 17016
rect 8627 16970 8695 17016
rect 8741 16970 8809 17016
rect 8855 16970 8923 17016
rect 8969 16970 9037 17016
rect 9083 16970 9151 17016
rect 9197 16970 9265 17016
rect 9311 16970 9379 17016
rect 9425 16970 9493 17016
rect 9539 16970 9607 17016
rect 9653 16970 9721 17016
rect 9767 16970 9835 17016
rect 9881 16970 9949 17016
rect 9995 16970 10063 17016
rect 10109 16970 10177 17016
rect 10223 16970 10291 17016
rect 10337 16970 10405 17016
rect 10451 16970 10519 17016
rect 10565 16970 10633 17016
rect 10679 16970 10747 17016
rect 10793 16970 10861 17016
rect 10907 16970 10975 17016
rect 11021 16970 11089 17016
rect 11135 16970 11203 17016
rect 11249 16970 11317 17016
rect 11363 16970 11431 17016
rect 11477 16970 11545 17016
rect 11591 16970 11659 17016
rect 11705 16970 11773 17016
rect 11819 16970 11927 17016
rect 11973 16970 12041 17016
rect 12087 16970 12098 17016
rect 1576 16902 12098 16970
rect 1576 16856 1587 16902
rect 1633 16856 1701 16902
rect 1747 16856 1855 16902
rect 1901 16856 1969 16902
rect 2015 16856 2083 16902
rect 2129 16856 2197 16902
rect 2243 16856 2311 16902
rect 2357 16856 2425 16902
rect 2471 16856 2539 16902
rect 2585 16856 2653 16902
rect 2699 16856 2767 16902
rect 2813 16856 2881 16902
rect 2927 16856 2995 16902
rect 3041 16856 3109 16902
rect 3155 16856 3223 16902
rect 3269 16856 3337 16902
rect 3383 16856 3451 16902
rect 3497 16856 3565 16902
rect 3611 16856 3679 16902
rect 3725 16856 3793 16902
rect 3839 16856 3907 16902
rect 3953 16856 4021 16902
rect 4067 16856 4135 16902
rect 4181 16856 4249 16902
rect 4295 16856 4363 16902
rect 4409 16856 4477 16902
rect 4523 16856 4591 16902
rect 4637 16856 4705 16902
rect 4751 16856 4819 16902
rect 4865 16856 4933 16902
rect 4979 16856 5047 16902
rect 5093 16856 5161 16902
rect 5207 16856 5275 16902
rect 5321 16856 5389 16902
rect 5435 16856 5503 16902
rect 5549 16856 5617 16902
rect 5663 16856 5731 16902
rect 5777 16856 5845 16902
rect 5891 16856 5959 16902
rect 6005 16856 6073 16902
rect 6119 16856 6187 16902
rect 6233 16856 6301 16902
rect 6347 16856 6415 16902
rect 6461 16856 6529 16902
rect 6575 16856 6643 16902
rect 6689 16856 6757 16902
rect 6803 16856 6871 16902
rect 6917 16856 6985 16902
rect 7031 16856 7099 16902
rect 7145 16856 7213 16902
rect 7259 16856 7327 16902
rect 7373 16856 7441 16902
rect 7487 16856 7555 16902
rect 7601 16856 7669 16902
rect 7715 16856 7783 16902
rect 7829 16856 7897 16902
rect 7943 16856 8011 16902
rect 8057 16856 8125 16902
rect 8171 16856 8239 16902
rect 8285 16856 8353 16902
rect 8399 16856 8467 16902
rect 8513 16856 8581 16902
rect 8627 16856 8695 16902
rect 8741 16856 8809 16902
rect 8855 16856 8923 16902
rect 8969 16856 9037 16902
rect 9083 16856 9151 16902
rect 9197 16856 9265 16902
rect 9311 16856 9379 16902
rect 9425 16856 9493 16902
rect 9539 16856 9607 16902
rect 9653 16856 9721 16902
rect 9767 16856 9835 16902
rect 9881 16856 9949 16902
rect 9995 16856 10063 16902
rect 10109 16856 10177 16902
rect 10223 16856 10291 16902
rect 10337 16856 10405 16902
rect 10451 16856 10519 16902
rect 10565 16856 10633 16902
rect 10679 16856 10747 16902
rect 10793 16856 10861 16902
rect 10907 16856 10975 16902
rect 11021 16856 11089 16902
rect 11135 16856 11203 16902
rect 11249 16856 11317 16902
rect 11363 16856 11431 16902
rect 11477 16856 11545 16902
rect 11591 16856 11659 16902
rect 11705 16856 11773 16902
rect 11819 16856 11927 16902
rect 11973 16856 12041 16902
rect 12087 16856 12098 16902
rect 1576 16844 12098 16856
rect 1576 16788 1758 16844
rect 1576 16742 1587 16788
rect 1633 16742 1701 16788
rect 1747 16742 1758 16788
rect 1576 16681 1758 16742
rect 11916 16788 12098 16844
rect 11916 16742 11927 16788
rect 11973 16742 12041 16788
rect 12087 16742 12098 16788
rect 11916 16674 12098 16742
rect 11916 16628 11927 16674
rect 11973 16628 12041 16674
rect 12087 16628 12098 16674
rect 306 16441 11446 16573
rect 306 16430 4138 16441
rect 306 16411 2233 16430
rect 306 5279 466 16411
rect 2222 16384 2233 16411
rect 4127 16384 4138 16430
rect 2222 16373 4138 16384
rect 4658 16430 6574 16441
rect 4658 16384 4669 16430
rect 6563 16384 6574 16430
rect 4658 16373 6574 16384
rect 7094 16430 9010 16441
rect 7094 16384 7105 16430
rect 8999 16384 9010 16430
rect 7094 16373 9010 16384
rect 9530 16430 11446 16441
rect 9530 16384 9541 16430
rect 11435 16384 11446 16430
rect 9530 16373 11446 16384
rect 11916 16560 12098 16628
rect 11916 16514 11927 16560
rect 11973 16514 12041 16560
rect 12087 16514 12098 16560
rect 11916 16446 12098 16514
rect 11916 16400 11927 16446
rect 11973 16400 12041 16446
rect 12087 16400 12098 16446
rect 1576 16314 2162 16351
rect 1576 16218 2105 16314
rect 1576 16172 1587 16218
rect 1633 16172 1701 16218
rect 1747 16172 2105 16218
rect 1576 16104 2105 16172
rect 1576 16058 1587 16104
rect 1633 16058 1701 16104
rect 1747 16058 2105 16104
rect 1576 15990 2105 16058
rect 1576 15944 1587 15990
rect 1633 15944 1701 15990
rect 1747 15944 2105 15990
rect 1576 15876 2105 15944
rect 1576 15830 1587 15876
rect 1633 15830 1701 15876
rect 1747 15830 2105 15876
rect 1576 15762 2105 15830
rect 1576 15716 1587 15762
rect 1633 15716 1701 15762
rect 1747 15716 2105 15762
rect 1576 15648 2105 15716
rect 1576 15602 1587 15648
rect 1633 15602 1701 15648
rect 1747 15602 2105 15648
rect 1576 15534 2105 15602
rect 1576 15488 1587 15534
rect 1633 15488 1701 15534
rect 1747 15488 2105 15534
rect 1576 15420 2105 15488
rect 1576 15374 1587 15420
rect 1633 15374 1701 15420
rect 1747 15374 2105 15420
rect 1576 15306 2105 15374
rect 1576 15260 1587 15306
rect 1633 15260 1701 15306
rect 1747 15260 2105 15306
rect 1576 15192 2105 15260
rect 1576 15146 1587 15192
rect 1633 15146 1701 15192
rect 1747 15146 2105 15192
rect 1576 15078 2105 15146
rect 1576 15032 1587 15078
rect 1633 15032 1701 15078
rect 1747 15032 2105 15078
rect 1576 14964 2105 15032
rect 1576 14918 1587 14964
rect 1633 14918 1701 14964
rect 1747 14918 2105 14964
rect 1576 14850 2105 14918
rect 1576 14804 1587 14850
rect 1633 14804 1701 14850
rect 1747 14804 2105 14850
rect 1576 14736 2105 14804
rect 1576 14690 1587 14736
rect 1633 14690 1701 14736
rect 1747 14690 2105 14736
rect 1576 14622 2105 14690
rect 1576 14576 1587 14622
rect 1633 14576 1701 14622
rect 1747 14576 2105 14622
rect 1576 14508 2105 14576
rect 1576 14462 1587 14508
rect 1633 14462 1701 14508
rect 1747 14462 2105 14508
rect 1576 14394 2105 14462
rect 1576 14348 1587 14394
rect 1633 14348 1701 14394
rect 1747 14348 2105 14394
rect 1576 14280 2105 14348
rect 1576 14234 1587 14280
rect 1633 14234 1701 14280
rect 1747 14234 2105 14280
rect 1576 14166 2105 14234
rect 1576 14120 1587 14166
rect 1633 14120 1701 14166
rect 1747 14120 2105 14166
rect 1576 14052 2105 14120
rect 1576 14006 1587 14052
rect 1633 14006 1701 14052
rect 1747 14006 2105 14052
rect 1576 13938 2105 14006
rect 1576 13892 1587 13938
rect 1633 13892 1701 13938
rect 1747 13892 2105 13938
rect 1576 13824 2105 13892
rect 1576 13778 1587 13824
rect 1633 13778 1701 13824
rect 1747 13778 2105 13824
rect 1576 13710 2105 13778
rect 1576 13664 1587 13710
rect 1633 13664 1701 13710
rect 1747 13664 2105 13710
rect 1576 13596 2105 13664
rect 1576 13550 1587 13596
rect 1633 13550 1701 13596
rect 1747 13550 2105 13596
rect 1576 13482 2105 13550
rect 1576 13436 1587 13482
rect 1633 13436 1701 13482
rect 1747 13436 2105 13482
rect 1576 13368 2105 13436
rect 1576 13322 1587 13368
rect 1633 13322 1701 13368
rect 1747 13322 2105 13368
rect 1576 13254 2105 13322
rect 1576 13208 1587 13254
rect 1633 13208 1701 13254
rect 1747 13208 2105 13254
rect 1576 13140 2105 13208
rect 1576 13094 1587 13140
rect 1633 13094 1701 13140
rect 1747 13094 2105 13140
rect 1576 13026 2105 13094
rect 1576 12980 1587 13026
rect 1633 12980 1701 13026
rect 1747 12980 2105 13026
rect 1576 12912 2105 12980
rect 1576 12866 1587 12912
rect 1633 12866 1701 12912
rect 1747 12866 2105 12912
rect 1576 12798 2105 12866
rect 1576 12752 1587 12798
rect 1633 12752 1701 12798
rect 1747 12752 2105 12798
rect 1576 12684 2105 12752
rect 1576 12638 1587 12684
rect 1633 12638 1701 12684
rect 1747 12638 2105 12684
rect 1576 12570 2105 12638
rect 1576 12524 1587 12570
rect 1633 12524 1701 12570
rect 1747 12524 2105 12570
rect 1576 12456 2105 12524
rect 1576 12410 1587 12456
rect 1633 12410 1701 12456
rect 1747 12410 2105 12456
rect 1576 12342 2105 12410
rect 1576 12296 1587 12342
rect 1633 12296 1701 12342
rect 1747 12296 2105 12342
rect 1576 12228 2105 12296
rect 1576 12182 1587 12228
rect 1633 12182 1701 12228
rect 1747 12182 2105 12228
rect 1576 12114 2105 12182
rect 1576 12068 1587 12114
rect 1633 12068 1701 12114
rect 1747 12068 2105 12114
rect 1576 12000 2105 12068
rect 1576 11954 1587 12000
rect 1633 11954 1701 12000
rect 1747 11954 2105 12000
rect 1576 11886 2105 11954
rect 1576 11840 1587 11886
rect 1633 11840 1701 11886
rect 1747 11840 2105 11886
rect 1576 11772 2105 11840
rect 1576 11726 1587 11772
rect 1633 11726 1701 11772
rect 1747 11726 2105 11772
rect 1576 11658 2105 11726
rect 1576 11612 1587 11658
rect 1633 11612 1701 11658
rect 1747 11612 2105 11658
rect 1576 11544 2105 11612
rect 1576 11498 1587 11544
rect 1633 11498 1701 11544
rect 1747 11498 2105 11544
rect 1576 11430 2105 11498
rect 1576 11384 1587 11430
rect 1633 11384 1701 11430
rect 1747 11388 2105 11430
rect 2151 11388 2162 16314
rect 1747 11384 2162 11388
rect 1576 11316 2162 11384
rect 2680 11329 3680 16373
rect 4198 16314 4598 16351
rect 4198 11388 4209 16314
rect 4255 11388 4541 16314
rect 4587 11388 4598 16314
rect 1576 11270 1587 11316
rect 1633 11270 1701 11316
rect 1747 11270 2162 11316
rect 1576 11202 2162 11270
rect 2222 11318 4138 11329
rect 2222 11272 2233 11318
rect 4127 11272 4138 11318
rect 2222 11261 4138 11272
rect 1576 11156 1587 11202
rect 1633 11156 1701 11202
rect 1747 11201 2162 11202
rect 4198 11201 4598 11388
rect 5116 11329 6116 16373
rect 6634 16314 7034 16351
rect 6634 11388 6645 16314
rect 6691 11388 6977 16314
rect 7023 11388 7034 16314
rect 4658 11318 6574 11329
rect 4658 11272 4669 11318
rect 6563 11272 6574 11318
rect 4658 11261 6574 11272
rect 6634 11201 7034 11388
rect 7552 11329 8552 16373
rect 9070 16314 9470 16351
rect 9070 11388 9081 16314
rect 9127 11388 9413 16314
rect 9459 11388 9470 16314
rect 7094 11318 9010 11329
rect 7094 11272 7105 11318
rect 8999 11272 9010 11318
rect 7094 11261 9010 11272
rect 9070 11201 9470 11388
rect 9988 11329 10988 16373
rect 11916 16351 12098 16400
rect 11506 16332 12098 16351
rect 11506 16314 11927 16332
rect 11506 11388 11517 16314
rect 11563 16286 11927 16314
rect 11973 16286 12041 16332
rect 12087 16286 12098 16332
rect 11563 16218 12098 16286
rect 11563 16172 11927 16218
rect 11973 16172 12041 16218
rect 12087 16172 12098 16218
rect 11563 16104 12098 16172
rect 11563 16058 11927 16104
rect 11973 16058 12041 16104
rect 12087 16058 12098 16104
rect 11563 15990 12098 16058
rect 11563 15944 11927 15990
rect 11973 15944 12041 15990
rect 12087 15944 12098 15990
rect 11563 15876 12098 15944
rect 11563 15830 11927 15876
rect 11973 15830 12041 15876
rect 12087 15830 12098 15876
rect 11563 15762 12098 15830
rect 11563 15716 11927 15762
rect 11973 15716 12041 15762
rect 12087 15716 12098 15762
rect 11563 15648 12098 15716
rect 11563 15602 11927 15648
rect 11973 15602 12041 15648
rect 12087 15602 12098 15648
rect 11563 15534 12098 15602
rect 11563 15488 11927 15534
rect 11973 15488 12041 15534
rect 12087 15488 12098 15534
rect 11563 15420 12098 15488
rect 11563 15374 11927 15420
rect 11973 15374 12041 15420
rect 12087 15374 12098 15420
rect 11563 15306 12098 15374
rect 11563 15260 11927 15306
rect 11973 15260 12041 15306
rect 12087 15260 12098 15306
rect 11563 15192 12098 15260
rect 11563 15146 11927 15192
rect 11973 15146 12041 15192
rect 12087 15146 12098 15192
rect 11563 15078 12098 15146
rect 11563 15032 11927 15078
rect 11973 15032 12041 15078
rect 12087 15032 12098 15078
rect 11563 14964 12098 15032
rect 11563 14918 11927 14964
rect 11973 14918 12041 14964
rect 12087 14918 12098 14964
rect 11563 14850 12098 14918
rect 11563 14804 11927 14850
rect 11973 14804 12041 14850
rect 12087 14804 12098 14850
rect 11563 14736 12098 14804
rect 11563 14690 11927 14736
rect 11973 14690 12041 14736
rect 12087 14690 12098 14736
rect 11563 14622 12098 14690
rect 11563 14576 11927 14622
rect 11973 14576 12041 14622
rect 12087 14576 12098 14622
rect 11563 14508 12098 14576
rect 11563 14462 11927 14508
rect 11973 14462 12041 14508
rect 12087 14462 12098 14508
rect 11563 14394 12098 14462
rect 11563 14348 11927 14394
rect 11973 14348 12041 14394
rect 12087 14348 12098 14394
rect 11563 14280 12098 14348
rect 11563 14234 11927 14280
rect 11973 14234 12041 14280
rect 12087 14234 12098 14280
rect 11563 14166 12098 14234
rect 11563 14120 11927 14166
rect 11973 14120 12041 14166
rect 12087 14120 12098 14166
rect 11563 14052 12098 14120
rect 11563 14006 11927 14052
rect 11973 14006 12041 14052
rect 12087 14006 12098 14052
rect 11563 13938 12098 14006
rect 11563 13892 11927 13938
rect 11973 13892 12041 13938
rect 12087 13892 12098 13938
rect 11563 13824 12098 13892
rect 11563 13778 11927 13824
rect 11973 13778 12041 13824
rect 12087 13778 12098 13824
rect 11563 13710 12098 13778
rect 11563 13664 11927 13710
rect 11973 13664 12041 13710
rect 12087 13664 12098 13710
rect 11563 13596 12098 13664
rect 11563 13550 11927 13596
rect 11973 13550 12041 13596
rect 12087 13550 12098 13596
rect 11563 13482 12098 13550
rect 11563 13436 11927 13482
rect 11973 13436 12041 13482
rect 12087 13436 12098 13482
rect 11563 13368 12098 13436
rect 11563 13322 11927 13368
rect 11973 13322 12041 13368
rect 12087 13322 12098 13368
rect 11563 13254 12098 13322
rect 11563 13208 11927 13254
rect 11973 13208 12041 13254
rect 12087 13208 12098 13254
rect 11563 13140 12098 13208
rect 11563 13094 11927 13140
rect 11973 13094 12041 13140
rect 12087 13094 12098 13140
rect 11563 13026 12098 13094
rect 11563 12980 11927 13026
rect 11973 12980 12041 13026
rect 12087 12980 12098 13026
rect 11563 12912 12098 12980
rect 11563 12866 11927 12912
rect 11973 12866 12041 12912
rect 12087 12866 12098 12912
rect 11563 12798 12098 12866
rect 11563 12752 11927 12798
rect 11973 12752 12041 12798
rect 12087 12752 12098 12798
rect 11563 12684 12098 12752
rect 11563 12638 11927 12684
rect 11973 12638 12041 12684
rect 12087 12638 12098 12684
rect 11563 12570 12098 12638
rect 11563 12524 11927 12570
rect 11973 12524 12041 12570
rect 12087 12524 12098 12570
rect 11563 12456 12098 12524
rect 11563 12410 11927 12456
rect 11973 12410 12041 12456
rect 12087 12410 12098 12456
rect 11563 12342 12098 12410
rect 11563 12296 11927 12342
rect 11973 12296 12041 12342
rect 12087 12296 12098 12342
rect 11563 12228 12098 12296
rect 11563 12182 11927 12228
rect 11973 12182 12041 12228
rect 12087 12182 12098 12228
rect 11563 12114 12098 12182
rect 11563 12068 11927 12114
rect 11973 12068 12041 12114
rect 12087 12068 12098 12114
rect 11563 12000 12098 12068
rect 11563 11954 11927 12000
rect 11973 11954 12041 12000
rect 12087 11954 12098 12000
rect 11563 11886 12098 11954
rect 11563 11840 11927 11886
rect 11973 11840 12041 11886
rect 12087 11840 12098 11886
rect 11563 11772 12098 11840
rect 11563 11726 11927 11772
rect 11973 11726 12041 11772
rect 12087 11726 12098 11772
rect 11563 11658 12098 11726
rect 11563 11612 11927 11658
rect 11973 11612 12041 11658
rect 12087 11612 12098 11658
rect 11563 11544 12098 11612
rect 11563 11498 11927 11544
rect 11973 11498 12041 11544
rect 12087 11498 12098 11544
rect 11563 11430 12098 11498
rect 11563 11388 11927 11430
rect 11506 11384 11927 11388
rect 11973 11384 12041 11430
rect 12087 11384 12098 11430
rect 9530 11318 11446 11329
rect 9530 11272 9541 11318
rect 11435 11272 11446 11318
rect 9530 11261 11446 11272
rect 11506 11316 12098 11384
rect 11506 11270 11927 11316
rect 11973 11270 12041 11316
rect 12087 11270 12098 11316
rect 11506 11202 12098 11270
rect 11506 11201 11927 11202
rect 1747 11156 11927 11201
rect 11973 11156 12041 11202
rect 12087 11156 12098 11202
rect 1576 11088 12098 11156
rect 1576 11042 1587 11088
rect 1633 11042 1701 11088
rect 1747 11042 11927 11088
rect 11973 11042 12041 11088
rect 12087 11042 12098 11088
rect 1576 10974 12098 11042
rect 1576 10928 1587 10974
rect 1633 10928 1701 10974
rect 1747 10928 11927 10974
rect 11973 10928 12041 10974
rect 12087 10928 12098 10974
rect 1576 10925 12098 10928
rect 1576 10879 1855 10925
rect 1901 10879 1969 10925
rect 2015 10879 2083 10925
rect 2129 10879 2197 10925
rect 2243 10879 2311 10925
rect 2357 10879 2425 10925
rect 2471 10879 2539 10925
rect 2585 10879 2653 10925
rect 2699 10879 2767 10925
rect 2813 10879 2881 10925
rect 2927 10879 2995 10925
rect 3041 10879 3109 10925
rect 3155 10879 3223 10925
rect 3269 10879 3337 10925
rect 3383 10879 3451 10925
rect 3497 10879 3565 10925
rect 3611 10879 3679 10925
rect 3725 10879 3793 10925
rect 3839 10879 3907 10925
rect 3953 10879 4021 10925
rect 4067 10879 4135 10925
rect 4181 10879 4249 10925
rect 4295 10879 4363 10925
rect 4409 10879 4477 10925
rect 4523 10879 4591 10925
rect 4637 10879 4705 10925
rect 4751 10879 4819 10925
rect 4865 10879 4933 10925
rect 4979 10879 5047 10925
rect 5093 10879 5161 10925
rect 5207 10879 5275 10925
rect 5321 10879 5389 10925
rect 5435 10879 5503 10925
rect 5549 10879 5617 10925
rect 5663 10879 5731 10925
rect 5777 10879 5845 10925
rect 5891 10879 5959 10925
rect 6005 10879 6073 10925
rect 6119 10879 6187 10925
rect 6233 10879 6301 10925
rect 6347 10879 6415 10925
rect 6461 10879 6529 10925
rect 6575 10879 6643 10925
rect 6689 10879 6757 10925
rect 6803 10879 6871 10925
rect 6917 10879 6985 10925
rect 7031 10879 7099 10925
rect 7145 10879 7213 10925
rect 7259 10879 7327 10925
rect 7373 10879 7441 10925
rect 7487 10879 7555 10925
rect 7601 10879 7669 10925
rect 7715 10879 7783 10925
rect 7829 10879 7897 10925
rect 7943 10879 8011 10925
rect 8057 10879 8125 10925
rect 8171 10879 8239 10925
rect 8285 10879 8353 10925
rect 8399 10879 8467 10925
rect 8513 10879 8581 10925
rect 8627 10879 8695 10925
rect 8741 10879 8809 10925
rect 8855 10879 8923 10925
rect 8969 10879 9037 10925
rect 9083 10879 9151 10925
rect 9197 10879 9265 10925
rect 9311 10879 9379 10925
rect 9425 10879 9493 10925
rect 9539 10879 9607 10925
rect 9653 10879 9721 10925
rect 9767 10879 9835 10925
rect 9881 10879 9949 10925
rect 9995 10879 10063 10925
rect 10109 10879 10177 10925
rect 10223 10879 10291 10925
rect 10337 10879 10405 10925
rect 10451 10879 10519 10925
rect 10565 10879 10633 10925
rect 10679 10879 10747 10925
rect 10793 10879 10861 10925
rect 10907 10879 10975 10925
rect 11021 10879 11089 10925
rect 11135 10879 11203 10925
rect 11249 10879 11317 10925
rect 11363 10879 11431 10925
rect 11477 10879 11545 10925
rect 11591 10879 11659 10925
rect 11705 10879 11773 10925
rect 11819 10879 12098 10925
rect 1576 10860 12098 10879
rect 1576 10814 1587 10860
rect 1633 10814 1701 10860
rect 1747 10814 11927 10860
rect 11973 10814 12041 10860
rect 12087 10814 12098 10860
rect 1576 10811 12098 10814
rect 1576 10765 1855 10811
rect 1901 10765 1969 10811
rect 2015 10765 2083 10811
rect 2129 10765 2197 10811
rect 2243 10765 2311 10811
rect 2357 10765 2425 10811
rect 2471 10765 2539 10811
rect 2585 10765 2653 10811
rect 2699 10765 2767 10811
rect 2813 10765 2881 10811
rect 2927 10765 2995 10811
rect 3041 10765 3109 10811
rect 3155 10765 3223 10811
rect 3269 10765 3337 10811
rect 3383 10765 3451 10811
rect 3497 10765 3565 10811
rect 3611 10765 3679 10811
rect 3725 10765 3793 10811
rect 3839 10765 3907 10811
rect 3953 10765 4021 10811
rect 4067 10765 4135 10811
rect 4181 10765 4249 10811
rect 4295 10765 4363 10811
rect 4409 10765 4477 10811
rect 4523 10765 4591 10811
rect 4637 10765 4705 10811
rect 4751 10765 4819 10811
rect 4865 10765 4933 10811
rect 4979 10765 5047 10811
rect 5093 10765 5161 10811
rect 5207 10765 5275 10811
rect 5321 10765 5389 10811
rect 5435 10765 5503 10811
rect 5549 10765 5617 10811
rect 5663 10765 5731 10811
rect 5777 10765 5845 10811
rect 5891 10765 5959 10811
rect 6005 10765 6073 10811
rect 6119 10765 6187 10811
rect 6233 10765 6301 10811
rect 6347 10765 6415 10811
rect 6461 10765 6529 10811
rect 6575 10765 6643 10811
rect 6689 10765 6757 10811
rect 6803 10765 6871 10811
rect 6917 10765 6985 10811
rect 7031 10765 7099 10811
rect 7145 10765 7213 10811
rect 7259 10765 7327 10811
rect 7373 10765 7441 10811
rect 7487 10765 7555 10811
rect 7601 10765 7669 10811
rect 7715 10765 7783 10811
rect 7829 10765 7897 10811
rect 7943 10765 8011 10811
rect 8057 10765 8125 10811
rect 8171 10765 8239 10811
rect 8285 10765 8353 10811
rect 8399 10765 8467 10811
rect 8513 10765 8581 10811
rect 8627 10765 8695 10811
rect 8741 10765 8809 10811
rect 8855 10765 8923 10811
rect 8969 10765 9037 10811
rect 9083 10765 9151 10811
rect 9197 10765 9265 10811
rect 9311 10765 9379 10811
rect 9425 10765 9493 10811
rect 9539 10765 9607 10811
rect 9653 10765 9721 10811
rect 9767 10765 9835 10811
rect 9881 10765 9949 10811
rect 9995 10765 10063 10811
rect 10109 10765 10177 10811
rect 10223 10765 10291 10811
rect 10337 10765 10405 10811
rect 10451 10765 10519 10811
rect 10565 10765 10633 10811
rect 10679 10765 10747 10811
rect 10793 10765 10861 10811
rect 10907 10765 10975 10811
rect 11021 10765 11089 10811
rect 11135 10765 11203 10811
rect 11249 10765 11317 10811
rect 11363 10765 11431 10811
rect 11477 10765 11545 10811
rect 11591 10765 11659 10811
rect 11705 10765 11773 10811
rect 11819 10765 12098 10811
rect 1576 10746 12098 10765
rect 1576 10700 1587 10746
rect 1633 10700 1701 10746
rect 1747 10700 11927 10746
rect 11973 10700 12041 10746
rect 12087 10700 12098 10746
rect 1576 10632 12098 10700
rect 1576 10586 1587 10632
rect 1633 10586 1701 10632
rect 1747 10586 11927 10632
rect 11973 10586 12041 10632
rect 12087 10586 12098 10632
rect 1576 10518 12098 10586
rect 1576 10472 1587 10518
rect 1633 10472 1701 10518
rect 1747 10489 11927 10518
rect 1747 10472 2162 10489
rect 1576 10404 2162 10472
rect 1576 10358 1587 10404
rect 1633 10358 1701 10404
rect 1747 10358 2162 10404
rect 2222 10418 4138 10429
rect 2222 10372 2233 10418
rect 4127 10372 4138 10418
rect 2222 10361 4138 10372
rect 1576 10302 2162 10358
rect 1576 10290 2105 10302
rect 1576 10244 1587 10290
rect 1633 10244 1701 10290
rect 1747 10244 2105 10290
rect 1576 10176 2105 10244
rect 1576 10130 1587 10176
rect 1633 10130 1701 10176
rect 1747 10130 2105 10176
rect 1576 10062 2105 10130
rect 1576 10016 1587 10062
rect 1633 10016 1701 10062
rect 1747 10016 2105 10062
rect 1576 9948 2105 10016
rect 1576 9902 1587 9948
rect 1633 9902 1701 9948
rect 1747 9902 2105 9948
rect 1576 9834 2105 9902
rect 1576 9788 1587 9834
rect 1633 9788 1701 9834
rect 1747 9788 2105 9834
rect 1576 9720 2105 9788
rect 1576 9674 1587 9720
rect 1633 9674 1701 9720
rect 1747 9674 2105 9720
rect 1576 9606 2105 9674
rect 1576 9560 1587 9606
rect 1633 9560 1701 9606
rect 1747 9560 2105 9606
rect 1576 9492 2105 9560
rect 1576 9446 1587 9492
rect 1633 9446 1701 9492
rect 1747 9446 2105 9492
rect 1576 9378 2105 9446
rect 1576 9332 1587 9378
rect 1633 9332 1701 9378
rect 1747 9332 2105 9378
rect 1576 9264 2105 9332
rect 1576 9218 1587 9264
rect 1633 9218 1701 9264
rect 1747 9218 2105 9264
rect 1576 9150 2105 9218
rect 1576 9104 1587 9150
rect 1633 9104 1701 9150
rect 1747 9104 2105 9150
rect 1576 9036 2105 9104
rect 1576 8990 1587 9036
rect 1633 8990 1701 9036
rect 1747 8990 2105 9036
rect 1576 8922 2105 8990
rect 1576 8876 1587 8922
rect 1633 8876 1701 8922
rect 1747 8876 2105 8922
rect 1576 8808 2105 8876
rect 1576 8762 1587 8808
rect 1633 8762 1701 8808
rect 1747 8762 2105 8808
rect 1576 8694 2105 8762
rect 1576 8648 1587 8694
rect 1633 8648 1701 8694
rect 1747 8648 2105 8694
rect 1576 8580 2105 8648
rect 1576 8534 1587 8580
rect 1633 8534 1701 8580
rect 1747 8534 2105 8580
rect 1576 8466 2105 8534
rect 1576 8420 1587 8466
rect 1633 8420 1701 8466
rect 1747 8420 2105 8466
rect 1576 8352 2105 8420
rect 1576 8306 1587 8352
rect 1633 8306 1701 8352
rect 1747 8306 2105 8352
rect 1576 8238 2105 8306
rect 1576 8192 1587 8238
rect 1633 8192 1701 8238
rect 1747 8192 2105 8238
rect 1576 8124 2105 8192
rect 1576 8078 1587 8124
rect 1633 8078 1701 8124
rect 1747 8078 2105 8124
rect 1576 8010 2105 8078
rect 1576 7964 1587 8010
rect 1633 7964 1701 8010
rect 1747 7964 2105 8010
rect 1576 7896 2105 7964
rect 1576 7850 1587 7896
rect 1633 7850 1701 7896
rect 1747 7850 2105 7896
rect 1576 7782 2105 7850
rect 1576 7736 1587 7782
rect 1633 7736 1701 7782
rect 1747 7736 2105 7782
rect 1576 7668 2105 7736
rect 1576 7622 1587 7668
rect 1633 7622 1701 7668
rect 1747 7622 2105 7668
rect 1576 7554 2105 7622
rect 1576 7508 1587 7554
rect 1633 7508 1701 7554
rect 1747 7508 2105 7554
rect 1576 7440 2105 7508
rect 1576 7394 1587 7440
rect 1633 7394 1701 7440
rect 1747 7394 2105 7440
rect 1576 7326 2105 7394
rect 1576 7280 1587 7326
rect 1633 7280 1701 7326
rect 1747 7280 2105 7326
rect 1576 7212 2105 7280
rect 1576 7166 1587 7212
rect 1633 7166 1701 7212
rect 1747 7166 2105 7212
rect 1576 7098 2105 7166
rect 1576 7052 1587 7098
rect 1633 7052 1701 7098
rect 1747 7052 2105 7098
rect 1576 6984 2105 7052
rect 1576 6938 1587 6984
rect 1633 6938 1701 6984
rect 1747 6938 2105 6984
rect 1576 6870 2105 6938
rect 1576 6824 1587 6870
rect 1633 6824 1701 6870
rect 1747 6824 2105 6870
rect 1576 6756 2105 6824
rect 1576 6710 1587 6756
rect 1633 6710 1701 6756
rect 1747 6710 2105 6756
rect 1576 6642 2105 6710
rect 1576 6596 1587 6642
rect 1633 6596 1701 6642
rect 1747 6596 2105 6642
rect 1576 6528 2105 6596
rect 1576 6482 1587 6528
rect 1633 6482 1701 6528
rect 1747 6482 2105 6528
rect 1576 6414 2105 6482
rect 1576 6368 1587 6414
rect 1633 6368 1701 6414
rect 1747 6368 2105 6414
rect 1576 6300 2105 6368
rect 1576 6254 1587 6300
rect 1633 6254 1701 6300
rect 1747 6254 2105 6300
rect 1576 6186 2105 6254
rect 1576 6140 1587 6186
rect 1633 6140 1701 6186
rect 1747 6140 2105 6186
rect 1576 6072 2105 6140
rect 1576 6026 1587 6072
rect 1633 6026 1701 6072
rect 1747 6026 2105 6072
rect 1576 5958 2105 6026
rect 1576 5912 1587 5958
rect 1633 5912 1701 5958
rect 1747 5912 2105 5958
rect 1576 5844 2105 5912
rect 1576 5798 1587 5844
rect 1633 5798 1701 5844
rect 1747 5798 2105 5844
rect 1576 5730 2105 5798
rect 1576 5684 1587 5730
rect 1633 5684 1701 5730
rect 1747 5684 2105 5730
rect 1576 5616 2105 5684
rect 1576 5570 1587 5616
rect 1633 5570 1701 5616
rect 1747 5570 2105 5616
rect 1576 5502 2105 5570
rect 1576 5456 1587 5502
rect 1633 5456 1701 5502
rect 1747 5456 2105 5502
rect 1576 5376 2105 5456
rect 2151 5376 2162 10302
rect 1576 5339 2162 5376
rect 2680 5317 3680 10361
rect 4198 10302 4598 10489
rect 4658 10418 6574 10429
rect 4658 10372 4669 10418
rect 6563 10372 6574 10418
rect 4658 10361 6574 10372
rect 4198 5376 4209 10302
rect 4255 5376 4541 10302
rect 4587 5376 4598 10302
rect 4198 5339 4598 5376
rect 5116 5317 6116 10361
rect 6634 10302 7034 10489
rect 7094 10418 9010 10429
rect 7094 10372 7105 10418
rect 8999 10372 9010 10418
rect 7094 10361 9010 10372
rect 6634 5376 6645 10302
rect 6691 5376 6977 10302
rect 7023 5376 7034 10302
rect 6634 5339 7034 5376
rect 7552 5317 8552 10361
rect 9070 10302 9470 10489
rect 11506 10472 11927 10489
rect 11973 10472 12041 10518
rect 12087 10472 12098 10518
rect 9530 10418 11446 10429
rect 9530 10372 9541 10418
rect 11435 10372 11446 10418
rect 9530 10361 11446 10372
rect 11506 10404 12098 10472
rect 9070 5376 9081 10302
rect 9127 5376 9413 10302
rect 9459 5376 9470 10302
rect 9070 5339 9470 5376
rect 9988 5317 10988 10361
rect 11506 10358 11927 10404
rect 11973 10358 12041 10404
rect 12087 10358 12098 10404
rect 11506 10302 12098 10358
rect 11506 5376 11517 10302
rect 11563 10290 12098 10302
rect 11563 10244 11927 10290
rect 11973 10244 12041 10290
rect 12087 10244 12098 10290
rect 11563 10176 12098 10244
rect 11563 10130 11927 10176
rect 11973 10130 12041 10176
rect 12087 10130 12098 10176
rect 11563 10062 12098 10130
rect 11563 10016 11927 10062
rect 11973 10016 12041 10062
rect 12087 10016 12098 10062
rect 11563 9948 12098 10016
rect 11563 9902 11927 9948
rect 11973 9902 12041 9948
rect 12087 9902 12098 9948
rect 11563 9834 12098 9902
rect 11563 9788 11927 9834
rect 11973 9788 12041 9834
rect 12087 9788 12098 9834
rect 11563 9720 12098 9788
rect 11563 9674 11927 9720
rect 11973 9674 12041 9720
rect 12087 9674 12098 9720
rect 11563 9606 12098 9674
rect 11563 9560 11927 9606
rect 11973 9560 12041 9606
rect 12087 9560 12098 9606
rect 11563 9492 12098 9560
rect 11563 9446 11927 9492
rect 11973 9446 12041 9492
rect 12087 9446 12098 9492
rect 11563 9378 12098 9446
rect 11563 9332 11927 9378
rect 11973 9332 12041 9378
rect 12087 9332 12098 9378
rect 11563 9264 12098 9332
rect 11563 9218 11927 9264
rect 11973 9218 12041 9264
rect 12087 9218 12098 9264
rect 11563 9150 12098 9218
rect 11563 9104 11927 9150
rect 11973 9104 12041 9150
rect 12087 9104 12098 9150
rect 11563 9036 12098 9104
rect 11563 8990 11927 9036
rect 11973 8990 12041 9036
rect 12087 8990 12098 9036
rect 11563 8922 12098 8990
rect 11563 8876 11927 8922
rect 11973 8876 12041 8922
rect 12087 8876 12098 8922
rect 11563 8808 12098 8876
rect 11563 8762 11927 8808
rect 11973 8762 12041 8808
rect 12087 8762 12098 8808
rect 11563 8694 12098 8762
rect 11563 8648 11927 8694
rect 11973 8648 12041 8694
rect 12087 8648 12098 8694
rect 11563 8580 12098 8648
rect 11563 8534 11927 8580
rect 11973 8534 12041 8580
rect 12087 8534 12098 8580
rect 11563 8466 12098 8534
rect 11563 8420 11927 8466
rect 11973 8420 12041 8466
rect 12087 8420 12098 8466
rect 11563 8352 12098 8420
rect 11563 8306 11927 8352
rect 11973 8306 12041 8352
rect 12087 8306 12098 8352
rect 11563 8238 12098 8306
rect 11563 8192 11927 8238
rect 11973 8192 12041 8238
rect 12087 8192 12098 8238
rect 11563 8124 12098 8192
rect 11563 8078 11927 8124
rect 11973 8078 12041 8124
rect 12087 8078 12098 8124
rect 11563 8010 12098 8078
rect 11563 7964 11927 8010
rect 11973 7964 12041 8010
rect 12087 7964 12098 8010
rect 11563 7896 12098 7964
rect 11563 7850 11927 7896
rect 11973 7850 12041 7896
rect 12087 7850 12098 7896
rect 11563 7782 12098 7850
rect 11563 7736 11927 7782
rect 11973 7736 12041 7782
rect 12087 7736 12098 7782
rect 11563 7668 12098 7736
rect 11563 7622 11927 7668
rect 11973 7622 12041 7668
rect 12087 7622 12098 7668
rect 11563 7554 12098 7622
rect 11563 7508 11927 7554
rect 11973 7508 12041 7554
rect 12087 7508 12098 7554
rect 11563 7440 12098 7508
rect 11563 7394 11927 7440
rect 11973 7394 12041 7440
rect 12087 7394 12098 7440
rect 11563 7326 12098 7394
rect 11563 7280 11927 7326
rect 11973 7280 12041 7326
rect 12087 7280 12098 7326
rect 11563 7212 12098 7280
rect 11563 7166 11927 7212
rect 11973 7166 12041 7212
rect 12087 7166 12098 7212
rect 11563 7098 12098 7166
rect 11563 7052 11927 7098
rect 11973 7052 12041 7098
rect 12087 7052 12098 7098
rect 11563 6984 12098 7052
rect 11563 6938 11927 6984
rect 11973 6938 12041 6984
rect 12087 6938 12098 6984
rect 11563 6870 12098 6938
rect 11563 6824 11927 6870
rect 11973 6824 12041 6870
rect 12087 6824 12098 6870
rect 11563 6756 12098 6824
rect 11563 6710 11927 6756
rect 11973 6710 12041 6756
rect 12087 6710 12098 6756
rect 11563 6642 12098 6710
rect 11563 6596 11927 6642
rect 11973 6596 12041 6642
rect 12087 6596 12098 6642
rect 11563 6528 12098 6596
rect 11563 6482 11927 6528
rect 11973 6482 12041 6528
rect 12087 6482 12098 6528
rect 11563 6414 12098 6482
rect 11563 6368 11927 6414
rect 11973 6368 12041 6414
rect 12087 6368 12098 6414
rect 11563 6300 12098 6368
rect 11563 6254 11927 6300
rect 11973 6254 12041 6300
rect 12087 6254 12098 6300
rect 11563 6186 12098 6254
rect 11563 6140 11927 6186
rect 11973 6140 12041 6186
rect 12087 6140 12098 6186
rect 11563 6072 12098 6140
rect 11563 6026 11927 6072
rect 11973 6026 12041 6072
rect 12087 6026 12098 6072
rect 11563 5958 12098 6026
rect 11563 5912 11927 5958
rect 11973 5912 12041 5958
rect 12087 5912 12098 5958
rect 11563 5844 12098 5912
rect 11563 5798 11927 5844
rect 11973 5798 12041 5844
rect 12087 5798 12098 5844
rect 11563 5730 12098 5798
rect 11563 5684 11927 5730
rect 11973 5684 12041 5730
rect 12087 5684 12098 5730
rect 11563 5616 12098 5684
rect 11563 5570 11927 5616
rect 11973 5570 12041 5616
rect 12087 5570 12098 5616
rect 11563 5502 12098 5570
rect 11563 5456 11927 5502
rect 11973 5456 12041 5502
rect 12087 5456 12098 5502
rect 11563 5388 12098 5456
rect 11563 5376 11927 5388
rect 11506 5342 11927 5376
rect 11973 5342 12041 5388
rect 12087 5342 12098 5388
rect 11506 5339 12098 5342
rect 2222 5306 4138 5317
rect 2222 5279 2233 5306
rect 306 5260 2233 5279
rect 4127 5260 4138 5306
rect 306 5249 4138 5260
rect 4658 5306 6574 5317
rect 4658 5260 4669 5306
rect 6563 5260 6574 5306
rect 4658 5249 6574 5260
rect 7094 5306 9010 5317
rect 7094 5260 7105 5306
rect 8999 5260 9010 5306
rect 7094 5249 9010 5260
rect 9530 5306 11446 5317
rect 9530 5260 9541 5306
rect 11435 5260 11446 5306
rect 9530 5249 11446 5260
rect 306 5117 11446 5249
rect 11916 5274 12098 5339
rect 11916 5228 11927 5274
rect 11973 5228 12041 5274
rect 12087 5228 12098 5274
rect 11916 5160 12098 5228
rect 43 4382 233 4393
rect 43 4336 54 4382
rect 100 4336 158 4382
rect 204 4336 233 4382
rect 43 4325 233 4336
rect 43 4228 111 4325
rect 43 4182 54 4228
rect 100 4182 111 4228
rect 43 4124 111 4182
rect 43 4078 54 4124
rect 100 4078 111 4124
rect 43 4020 111 4078
rect 43 3974 54 4020
rect 100 3974 111 4020
rect 43 3916 111 3974
rect 306 4052 466 5117
rect 11916 5114 11927 5160
rect 11973 5114 12041 5160
rect 12087 5114 12098 5160
rect 1576 5046 1758 5067
rect 1576 5000 1587 5046
rect 1633 5000 1701 5046
rect 1747 5000 1758 5046
rect 1576 4944 1758 5000
rect 11916 5046 12098 5114
rect 11916 5000 11927 5046
rect 11973 5000 12041 5046
rect 12087 5000 12098 5046
rect 11916 4944 12098 5000
rect 1576 4932 12098 4944
rect 1576 4886 1587 4932
rect 1633 4886 1701 4932
rect 1747 4886 1855 4932
rect 1901 4886 1969 4932
rect 2015 4886 2083 4932
rect 2129 4886 2197 4932
rect 2243 4886 2311 4932
rect 2357 4886 2425 4932
rect 2471 4886 2539 4932
rect 2585 4886 2653 4932
rect 2699 4886 2767 4932
rect 2813 4886 2881 4932
rect 2927 4886 2995 4932
rect 3041 4886 3109 4932
rect 3155 4886 3223 4932
rect 3269 4886 3337 4932
rect 3383 4886 3451 4932
rect 3497 4886 3565 4932
rect 3611 4886 3679 4932
rect 3725 4886 3793 4932
rect 3839 4886 3907 4932
rect 3953 4886 4021 4932
rect 4067 4886 4135 4932
rect 4181 4886 4249 4932
rect 4295 4886 4363 4932
rect 4409 4886 4477 4932
rect 4523 4886 4591 4932
rect 4637 4886 4705 4932
rect 4751 4886 4819 4932
rect 4865 4886 4933 4932
rect 4979 4886 5047 4932
rect 5093 4886 5161 4932
rect 5207 4886 5275 4932
rect 5321 4886 5389 4932
rect 5435 4886 5503 4932
rect 5549 4886 5617 4932
rect 5663 4886 5731 4932
rect 5777 4886 5845 4932
rect 5891 4886 5959 4932
rect 6005 4886 6073 4932
rect 6119 4886 6187 4932
rect 6233 4886 6301 4932
rect 6347 4886 6415 4932
rect 6461 4886 6529 4932
rect 6575 4886 6643 4932
rect 6689 4886 6757 4932
rect 6803 4886 6871 4932
rect 6917 4886 6985 4932
rect 7031 4886 7099 4932
rect 7145 4886 7213 4932
rect 7259 4886 7327 4932
rect 7373 4886 7441 4932
rect 7487 4886 7555 4932
rect 7601 4886 7669 4932
rect 7715 4886 7783 4932
rect 7829 4886 7897 4932
rect 7943 4886 8011 4932
rect 8057 4886 8125 4932
rect 8171 4886 8239 4932
rect 8285 4886 8353 4932
rect 8399 4886 8467 4932
rect 8513 4886 8581 4932
rect 8627 4886 8695 4932
rect 8741 4886 8809 4932
rect 8855 4886 8923 4932
rect 8969 4886 9037 4932
rect 9083 4886 9151 4932
rect 9197 4886 9265 4932
rect 9311 4886 9379 4932
rect 9425 4886 9493 4932
rect 9539 4886 9607 4932
rect 9653 4886 9721 4932
rect 9767 4886 9835 4932
rect 9881 4886 9949 4932
rect 9995 4886 10063 4932
rect 10109 4886 10177 4932
rect 10223 4886 10291 4932
rect 10337 4886 10405 4932
rect 10451 4886 10519 4932
rect 10565 4886 10633 4932
rect 10679 4886 10747 4932
rect 10793 4886 10861 4932
rect 10907 4886 10975 4932
rect 11021 4886 11089 4932
rect 11135 4886 11203 4932
rect 11249 4886 11317 4932
rect 11363 4886 11431 4932
rect 11477 4886 11545 4932
rect 11591 4886 11659 4932
rect 11705 4886 11773 4932
rect 11819 4886 11927 4932
rect 11973 4886 12041 4932
rect 12087 4886 12098 4932
rect 1576 4818 12098 4886
rect 1576 4772 1587 4818
rect 1633 4772 1701 4818
rect 1747 4772 1855 4818
rect 1901 4772 1969 4818
rect 2015 4772 2083 4818
rect 2129 4772 2197 4818
rect 2243 4772 2311 4818
rect 2357 4772 2425 4818
rect 2471 4772 2539 4818
rect 2585 4772 2653 4818
rect 2699 4772 2767 4818
rect 2813 4772 2881 4818
rect 2927 4772 2995 4818
rect 3041 4772 3109 4818
rect 3155 4772 3223 4818
rect 3269 4772 3337 4818
rect 3383 4772 3451 4818
rect 3497 4772 3565 4818
rect 3611 4772 3679 4818
rect 3725 4772 3793 4818
rect 3839 4772 3907 4818
rect 3953 4772 4021 4818
rect 4067 4772 4135 4818
rect 4181 4772 4249 4818
rect 4295 4772 4363 4818
rect 4409 4772 4477 4818
rect 4523 4772 4591 4818
rect 4637 4772 4705 4818
rect 4751 4772 4819 4818
rect 4865 4772 4933 4818
rect 4979 4772 5047 4818
rect 5093 4772 5161 4818
rect 5207 4772 5275 4818
rect 5321 4772 5389 4818
rect 5435 4772 5503 4818
rect 5549 4772 5617 4818
rect 5663 4772 5731 4818
rect 5777 4772 5845 4818
rect 5891 4772 5959 4818
rect 6005 4772 6073 4818
rect 6119 4772 6187 4818
rect 6233 4772 6301 4818
rect 6347 4772 6415 4818
rect 6461 4772 6529 4818
rect 6575 4772 6643 4818
rect 6689 4772 6757 4818
rect 6803 4772 6871 4818
rect 6917 4772 6985 4818
rect 7031 4772 7099 4818
rect 7145 4772 7213 4818
rect 7259 4772 7327 4818
rect 7373 4772 7441 4818
rect 7487 4772 7555 4818
rect 7601 4772 7669 4818
rect 7715 4772 7783 4818
rect 7829 4772 7897 4818
rect 7943 4772 8011 4818
rect 8057 4772 8125 4818
rect 8171 4772 8239 4818
rect 8285 4772 8353 4818
rect 8399 4772 8467 4818
rect 8513 4772 8581 4818
rect 8627 4772 8695 4818
rect 8741 4772 8809 4818
rect 8855 4772 8923 4818
rect 8969 4772 9037 4818
rect 9083 4772 9151 4818
rect 9197 4772 9265 4818
rect 9311 4772 9379 4818
rect 9425 4772 9493 4818
rect 9539 4772 9607 4818
rect 9653 4772 9721 4818
rect 9767 4772 9835 4818
rect 9881 4772 9949 4818
rect 9995 4772 10063 4818
rect 10109 4772 10177 4818
rect 10223 4772 10291 4818
rect 10337 4772 10405 4818
rect 10451 4772 10519 4818
rect 10565 4772 10633 4818
rect 10679 4772 10747 4818
rect 10793 4772 10861 4818
rect 10907 4772 10975 4818
rect 11021 4772 11089 4818
rect 11135 4772 11203 4818
rect 11249 4772 11317 4818
rect 11363 4772 11431 4818
rect 11477 4772 11545 4818
rect 11591 4772 11659 4818
rect 11705 4772 11773 4818
rect 11819 4772 11927 4818
rect 11973 4772 12041 4818
rect 12087 4772 12098 4818
rect 1576 4760 12098 4772
rect 540 4382 13631 4397
rect 540 4336 574 4382
rect 620 4336 678 4382
rect 724 4336 782 4382
rect 828 4336 886 4382
rect 932 4336 990 4382
rect 1036 4336 1094 4382
rect 1140 4336 1198 4382
rect 1244 4336 1302 4382
rect 1348 4336 1406 4382
rect 1452 4336 1510 4382
rect 1556 4336 1614 4382
rect 1660 4336 1718 4382
rect 1764 4336 1822 4382
rect 1868 4336 1926 4382
rect 1972 4336 2030 4382
rect 2076 4336 2134 4382
rect 2180 4336 2238 4382
rect 2284 4336 2342 4382
rect 2388 4336 2446 4382
rect 2492 4336 2550 4382
rect 2596 4336 2654 4382
rect 2700 4336 2758 4382
rect 2804 4336 2862 4382
rect 2908 4336 2966 4382
rect 3012 4336 3070 4382
rect 3116 4336 3174 4382
rect 3220 4336 3278 4382
rect 3324 4336 3382 4382
rect 3428 4336 3486 4382
rect 3532 4336 3590 4382
rect 3636 4336 3694 4382
rect 3740 4336 3798 4382
rect 3844 4336 3902 4382
rect 3948 4336 4006 4382
rect 4052 4336 4110 4382
rect 4156 4336 4214 4382
rect 4260 4336 4318 4382
rect 4364 4336 4422 4382
rect 4468 4336 4526 4382
rect 4572 4336 4630 4382
rect 4676 4336 4734 4382
rect 4780 4336 4838 4382
rect 4884 4336 4942 4382
rect 4988 4336 5046 4382
rect 5092 4336 5150 4382
rect 5196 4336 5254 4382
rect 5300 4336 5358 4382
rect 5404 4336 5462 4382
rect 5508 4336 5566 4382
rect 5612 4336 5670 4382
rect 5716 4336 5774 4382
rect 5820 4336 5878 4382
rect 5924 4336 5982 4382
rect 6028 4336 6086 4382
rect 6132 4336 6190 4382
rect 6236 4336 6294 4382
rect 6340 4336 6398 4382
rect 6444 4336 6502 4382
rect 6548 4336 6606 4382
rect 6652 4336 6710 4382
rect 6756 4336 6814 4382
rect 6860 4336 6918 4382
rect 6964 4336 7022 4382
rect 7068 4336 7126 4382
rect 7172 4336 7230 4382
rect 7276 4336 7334 4382
rect 7380 4336 7438 4382
rect 7484 4336 7542 4382
rect 7588 4336 7646 4382
rect 7692 4336 7750 4382
rect 7796 4336 7854 4382
rect 7900 4336 7958 4382
rect 8004 4336 8062 4382
rect 8108 4336 8166 4382
rect 8212 4336 8270 4382
rect 8316 4336 8374 4382
rect 8420 4336 8478 4382
rect 8524 4336 8582 4382
rect 8628 4336 8686 4382
rect 8732 4336 8790 4382
rect 8836 4336 8894 4382
rect 8940 4336 8998 4382
rect 9044 4336 9102 4382
rect 9148 4336 9206 4382
rect 9252 4336 9310 4382
rect 9356 4336 9414 4382
rect 9460 4336 9518 4382
rect 9564 4336 9622 4382
rect 9668 4336 9726 4382
rect 9772 4336 9830 4382
rect 9876 4336 9934 4382
rect 9980 4336 10038 4382
rect 10084 4336 10142 4382
rect 10188 4336 10246 4382
rect 10292 4336 10350 4382
rect 10396 4336 10454 4382
rect 10500 4336 10558 4382
rect 10604 4336 10662 4382
rect 10708 4336 10766 4382
rect 10812 4336 10870 4382
rect 10916 4336 10974 4382
rect 11020 4336 11078 4382
rect 11124 4336 11182 4382
rect 11228 4336 11286 4382
rect 11332 4336 11390 4382
rect 11436 4336 11494 4382
rect 11540 4336 11598 4382
rect 11644 4336 11702 4382
rect 11748 4336 11806 4382
rect 11852 4336 11910 4382
rect 11956 4336 12014 4382
rect 12060 4336 12118 4382
rect 12164 4336 12222 4382
rect 12268 4336 12326 4382
rect 12372 4336 12430 4382
rect 12476 4336 12534 4382
rect 12580 4336 12638 4382
rect 12684 4336 12742 4382
rect 12788 4336 12846 4382
rect 12892 4336 12950 4382
rect 12996 4336 13054 4382
rect 13100 4336 13158 4382
rect 13204 4336 13262 4382
rect 13308 4336 13366 4382
rect 13412 4336 13470 4382
rect 13516 4336 13574 4382
rect 13620 4336 13631 4382
rect 540 4321 13631 4336
rect 13563 4228 13631 4321
rect 13563 4182 13574 4228
rect 13620 4182 13631 4228
rect 13563 4124 13631 4182
rect 306 4006 366 4052
rect 412 4006 466 4052
rect 306 3951 466 4006
rect 13258 4052 13326 4107
rect 13258 4006 13269 4052
rect 13315 4006 13326 4052
rect 43 3870 54 3916
rect 100 3870 111 3916
rect 43 3812 111 3870
rect 43 3766 54 3812
rect 100 3766 111 3812
rect 43 3708 111 3766
rect 43 3662 54 3708
rect 100 3662 111 3708
rect 43 3604 111 3662
rect 43 3558 54 3604
rect 100 3558 111 3604
rect 43 3500 111 3558
rect 43 3454 54 3500
rect 100 3454 111 3500
rect 43 3396 111 3454
rect 43 3350 54 3396
rect 100 3350 111 3396
rect 355 3772 423 3827
rect 355 3726 366 3772
rect 412 3726 423 3772
rect 355 3492 423 3726
rect 13258 3772 13326 4006
rect 13258 3726 13269 3772
rect 13315 3726 13326 3772
rect 13258 3671 13326 3726
rect 13563 4078 13574 4124
rect 13620 4078 13631 4124
rect 13563 4020 13631 4078
rect 13563 3974 13574 4020
rect 13620 3974 13631 4020
rect 13563 3916 13631 3974
rect 13563 3870 13574 3916
rect 13620 3870 13631 3916
rect 13563 3812 13631 3870
rect 13563 3766 13574 3812
rect 13620 3766 13631 3812
rect 13563 3708 13631 3766
rect 13563 3662 13574 3708
rect 13620 3662 13631 3708
rect 13563 3604 13631 3662
rect 13563 3558 13574 3604
rect 13620 3558 13631 3604
rect 355 3446 366 3492
rect 412 3446 423 3492
rect 355 3391 423 3446
rect 13258 3492 13326 3547
rect 13258 3446 13269 3492
rect 13315 3446 13326 3492
rect 43 3292 111 3350
rect 43 3246 54 3292
rect 100 3246 111 3292
rect 43 3188 111 3246
rect 43 3142 54 3188
rect 100 3142 111 3188
rect 43 3084 111 3142
rect 43 3038 54 3084
rect 100 3038 111 3084
rect 43 2980 111 3038
rect 43 2934 54 2980
rect 100 2934 111 2980
rect 43 2876 111 2934
rect 43 2830 54 2876
rect 100 2830 111 2876
rect 355 3212 423 3267
rect 355 3166 366 3212
rect 412 3166 423 3212
rect 355 2932 423 3166
rect 13258 3212 13326 3446
rect 13258 3166 13269 3212
rect 13315 3166 13326 3212
rect 13258 3111 13326 3166
rect 13563 3500 13631 3558
rect 13563 3454 13574 3500
rect 13620 3454 13631 3500
rect 13563 3396 13631 3454
rect 13563 3350 13574 3396
rect 13620 3350 13631 3396
rect 13563 3292 13631 3350
rect 13563 3246 13574 3292
rect 13620 3246 13631 3292
rect 13563 3188 13631 3246
rect 13563 3142 13574 3188
rect 13620 3142 13631 3188
rect 13563 3084 13631 3142
rect 13563 3038 13574 3084
rect 13620 3038 13631 3084
rect 355 2886 366 2932
rect 412 2886 423 2932
rect 355 2831 423 2886
rect 13258 2932 13326 2987
rect 13258 2886 13269 2932
rect 13315 2886 13326 2932
rect 43 2772 111 2830
rect 43 2726 54 2772
rect 100 2726 111 2772
rect 43 2668 111 2726
rect 43 2622 54 2668
rect 100 2622 111 2668
rect 43 2564 111 2622
rect 43 2518 54 2564
rect 100 2518 111 2564
rect 43 2460 111 2518
rect 43 2414 54 2460
rect 100 2414 111 2460
rect 43 2356 111 2414
rect 43 2310 54 2356
rect 100 2310 111 2356
rect 43 2252 111 2310
rect 355 2652 423 2707
rect 355 2606 366 2652
rect 412 2606 423 2652
rect 355 2372 423 2606
rect 13258 2652 13326 2886
rect 13258 2606 13269 2652
rect 13315 2606 13326 2652
rect 13258 2551 13326 2606
rect 13563 2980 13631 3038
rect 13563 2934 13574 2980
rect 13620 2934 13631 2980
rect 13563 2876 13631 2934
rect 13563 2830 13574 2876
rect 13620 2830 13631 2876
rect 13563 2772 13631 2830
rect 13563 2726 13574 2772
rect 13620 2726 13631 2772
rect 13563 2668 13631 2726
rect 13563 2622 13574 2668
rect 13620 2622 13631 2668
rect 13563 2564 13631 2622
rect 13563 2518 13574 2564
rect 13620 2518 13631 2564
rect 13563 2460 13631 2518
rect 355 2326 366 2372
rect 412 2326 423 2372
rect 355 2271 423 2326
rect 13258 2372 13326 2427
rect 13258 2326 13269 2372
rect 13315 2326 13326 2372
rect 43 2206 54 2252
rect 100 2206 111 2252
rect 43 2148 111 2206
rect 43 2102 54 2148
rect 100 2102 111 2148
rect 43 2044 111 2102
rect 43 1998 54 2044
rect 100 1998 111 2044
rect 43 1940 111 1998
rect 43 1894 54 1940
rect 100 1894 111 1940
rect 43 1836 111 1894
rect 43 1790 54 1836
rect 100 1790 111 1836
rect 43 1732 111 1790
rect 43 1686 54 1732
rect 100 1686 111 1732
rect 355 2092 423 2147
rect 355 2046 366 2092
rect 412 2046 423 2092
rect 355 1812 423 2046
rect 13258 2092 13326 2326
rect 13258 2046 13269 2092
rect 13315 2046 13326 2092
rect 13258 1991 13326 2046
rect 13563 2414 13574 2460
rect 13620 2414 13631 2460
rect 13563 2356 13631 2414
rect 13563 2310 13574 2356
rect 13620 2310 13631 2356
rect 13563 2252 13631 2310
rect 13563 2206 13574 2252
rect 13620 2206 13631 2252
rect 13563 2148 13631 2206
rect 13563 2102 13574 2148
rect 13620 2102 13631 2148
rect 13563 2044 13631 2102
rect 13563 1998 13574 2044
rect 13620 1998 13631 2044
rect 13563 1940 13631 1998
rect 13563 1894 13574 1940
rect 13620 1894 13631 1940
rect 355 1766 366 1812
rect 412 1766 423 1812
rect 355 1711 423 1766
rect 13258 1812 13326 1867
rect 13258 1766 13269 1812
rect 13315 1766 13326 1812
rect 43 1628 111 1686
rect 43 1582 54 1628
rect 100 1582 111 1628
rect 43 1524 111 1582
rect 43 1478 54 1524
rect 100 1478 111 1524
rect 43 1420 111 1478
rect 43 1374 54 1420
rect 100 1374 111 1420
rect 43 1316 111 1374
rect 43 1270 54 1316
rect 100 1270 111 1316
rect 43 1212 111 1270
rect 43 1166 54 1212
rect 100 1166 111 1212
rect 43 1108 111 1166
rect 355 1532 423 1587
rect 355 1486 366 1532
rect 412 1486 423 1532
rect 355 1252 423 1486
rect 13258 1532 13326 1766
rect 13258 1486 13269 1532
rect 13315 1486 13326 1532
rect 13258 1431 13326 1486
rect 13563 1836 13631 1894
rect 13563 1790 13574 1836
rect 13620 1790 13631 1836
rect 13563 1732 13631 1790
rect 13563 1686 13574 1732
rect 13620 1686 13631 1732
rect 13563 1628 13631 1686
rect 13563 1582 13574 1628
rect 13620 1582 13631 1628
rect 13563 1524 13631 1582
rect 13563 1478 13574 1524
rect 13620 1478 13631 1524
rect 13563 1420 13631 1478
rect 13563 1374 13574 1420
rect 13620 1374 13631 1420
rect 13563 1316 13631 1374
rect 355 1206 366 1252
rect 412 1206 423 1252
rect 355 1151 423 1206
rect 13258 1252 13326 1307
rect 13258 1206 13269 1252
rect 13315 1206 13326 1252
rect 43 1062 54 1108
rect 100 1062 111 1108
rect 43 1004 111 1062
rect 43 958 54 1004
rect 100 958 111 1004
rect 43 900 111 958
rect 43 854 54 900
rect 100 854 111 900
rect 43 796 111 854
rect 43 750 54 796
rect 100 750 111 796
rect 43 657 111 750
rect 355 972 423 1027
rect 355 926 366 972
rect 412 926 423 972
rect 355 657 423 926
rect 13258 972 13326 1206
rect 13258 926 13269 972
rect 13315 926 13326 972
rect 13258 871 13326 926
rect 13563 1270 13574 1316
rect 13620 1270 13631 1316
rect 13563 1212 13631 1270
rect 13563 1166 13574 1212
rect 13620 1166 13631 1212
rect 13563 1108 13631 1166
rect 13563 1062 13574 1108
rect 13620 1062 13631 1108
rect 13563 1004 13631 1062
rect 13563 958 13574 1004
rect 13620 958 13631 1004
rect 13563 900 13631 958
rect 13563 854 13574 900
rect 13620 854 13631 900
rect 13563 796 13631 854
rect 13563 750 13574 796
rect 13620 750 13631 796
rect 13563 657 13631 750
rect 43 642 13631 657
rect 43 596 54 642
rect 100 596 158 642
rect 204 596 262 642
rect 308 596 366 642
rect 412 596 470 642
rect 516 596 574 642
rect 620 596 678 642
rect 724 596 782 642
rect 828 596 886 642
rect 932 596 990 642
rect 1036 596 1094 642
rect 1140 596 1198 642
rect 1244 596 1302 642
rect 1348 596 1406 642
rect 1452 596 1510 642
rect 1556 596 1614 642
rect 1660 596 1718 642
rect 1764 596 1822 642
rect 1868 596 1926 642
rect 1972 596 2030 642
rect 2076 596 2134 642
rect 2180 596 2238 642
rect 2284 596 2342 642
rect 2388 596 2446 642
rect 2492 596 2550 642
rect 2596 596 2654 642
rect 2700 596 2758 642
rect 2804 596 2862 642
rect 2908 596 2966 642
rect 3012 596 3070 642
rect 3116 596 3174 642
rect 3220 596 3278 642
rect 3324 596 3382 642
rect 3428 596 3486 642
rect 3532 596 3590 642
rect 3636 596 3694 642
rect 3740 596 3798 642
rect 3844 596 3902 642
rect 3948 596 4006 642
rect 4052 596 4110 642
rect 4156 596 4214 642
rect 4260 596 4318 642
rect 4364 596 4422 642
rect 4468 596 4526 642
rect 4572 596 4630 642
rect 4676 596 4734 642
rect 4780 596 4838 642
rect 4884 596 4942 642
rect 4988 596 5046 642
rect 5092 596 5150 642
rect 5196 596 5254 642
rect 5300 596 5358 642
rect 5404 596 5462 642
rect 5508 596 5566 642
rect 5612 596 5670 642
rect 5716 596 5774 642
rect 5820 596 5878 642
rect 5924 596 5982 642
rect 6028 596 6086 642
rect 6132 596 6190 642
rect 6236 596 6294 642
rect 6340 596 6398 642
rect 6444 596 6502 642
rect 6548 596 6606 642
rect 6652 596 6710 642
rect 6756 596 6814 642
rect 6860 596 6918 642
rect 6964 596 7022 642
rect 7068 596 7126 642
rect 7172 596 7230 642
rect 7276 596 7334 642
rect 7380 596 7438 642
rect 7484 596 7542 642
rect 7588 596 7646 642
rect 7692 596 7750 642
rect 7796 596 7854 642
rect 7900 596 7958 642
rect 8004 596 8062 642
rect 8108 596 8166 642
rect 8212 596 8270 642
rect 8316 596 8374 642
rect 8420 596 8478 642
rect 8524 596 8582 642
rect 8628 596 8686 642
rect 8732 596 8790 642
rect 8836 596 8894 642
rect 8940 596 8998 642
rect 9044 596 9102 642
rect 9148 596 9206 642
rect 9252 596 9310 642
rect 9356 596 9414 642
rect 9460 596 9518 642
rect 9564 596 9622 642
rect 9668 596 9726 642
rect 9772 596 9830 642
rect 9876 596 9934 642
rect 9980 596 10038 642
rect 10084 596 10142 642
rect 10188 596 10246 642
rect 10292 596 10350 642
rect 10396 596 10454 642
rect 10500 596 10558 642
rect 10604 596 10662 642
rect 10708 596 10766 642
rect 10812 596 10870 642
rect 10916 596 10974 642
rect 11020 596 11078 642
rect 11124 596 11182 642
rect 11228 596 11286 642
rect 11332 596 11390 642
rect 11436 596 11494 642
rect 11540 596 11598 642
rect 11644 596 11702 642
rect 11748 596 11806 642
rect 11852 596 11910 642
rect 11956 596 12014 642
rect 12060 596 12118 642
rect 12164 596 12222 642
rect 12268 596 12326 642
rect 12372 596 12430 642
rect 12476 596 12534 642
rect 12580 596 12638 642
rect 12684 596 12742 642
rect 12788 596 12846 642
rect 12892 596 12950 642
rect 12996 596 13054 642
rect 13100 596 13158 642
rect 13204 596 13262 642
rect 13308 596 13366 642
rect 13412 596 13470 642
rect 13516 596 13574 642
rect 13620 596 13631 642
rect 43 581 13631 596
<< labels >>
rlabel metal1 s 984 16493 984 16493 4 VRC
port 1 nsew
rlabel metal1 s 475 619 475 619 4 VPLUS
port 2 nsew
rlabel metal1 s 6835 10844 6835 10844 4 VMINUS
port 3 nsew
<< end >>
