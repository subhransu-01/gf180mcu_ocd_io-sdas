magic
tech gf180mcuD
magscale 1 10
timestamp 1764272961
<< nwell >>
rect 15980 51147 16518 51697
<< nmos >>
rect 16224 50941 16280 51061
<< pmos >>
rect 16224 51233 16280 51473
<< ndiff >>
rect 16135 51048 16224 51061
rect 16135 50956 16149 51048
rect 16195 50956 16224 51048
rect 16135 50941 16224 50956
rect 16280 51047 16368 51061
rect 16280 50955 16309 51047
rect 16355 50955 16368 51047
rect 16280 50941 16368 50955
<< pdiff >>
rect 16131 51459 16224 51473
rect 16131 51246 16144 51459
rect 16190 51246 16224 51459
rect 16131 51233 16224 51246
rect 16280 51459 16368 51473
rect 16280 51246 16309 51459
rect 16355 51246 16368 51459
rect 16280 51233 16368 51246
<< ndiffc >>
rect 16149 50956 16195 51048
rect 16309 50955 16355 51047
<< pdiffc >>
rect 16144 51246 16190 51459
rect 16309 51246 16355 51459
<< psubdiff >>
rect 16066 50862 16432 50875
rect 16066 50816 16079 50862
rect 16125 50816 16373 50862
rect 16419 50816 16432 50862
rect 16066 50803 16432 50816
<< nsubdiff >>
rect 16066 51598 16432 51611
rect 16066 51552 16079 51598
rect 16125 51552 16373 51598
rect 16419 51552 16432 51598
rect 16066 51539 16432 51552
<< psubdiffcont >>
rect 16079 50816 16125 50862
rect 16373 50816 16419 50862
<< nsubdiffcont >>
rect 16079 51552 16125 51598
rect 16373 51552 16419 51598
<< polysilicon >>
rect 16224 51473 16280 51519
rect 16224 51178 16280 51233
rect 16119 51165 16280 51178
rect 16119 51119 16132 51165
rect 16252 51119 16280 51165
rect 16119 51106 16280 51119
rect 16224 51061 16280 51106
rect 16224 50897 16280 50941
<< polycontact >>
rect 16132 51119 16252 51165
<< metal1 >>
rect 16066 51598 16432 51611
rect 16066 51552 16079 51598
rect 16125 51552 16373 51598
rect 16419 51552 16432 51598
rect 16066 51536 16432 51552
rect 16144 51459 16190 51536
rect 16144 51235 16190 51246
rect 16309 51459 16355 51470
rect 16121 51119 16132 51165
rect 16252 51119 16263 51165
rect 16149 51048 16195 51059
rect 16149 50879 16195 50956
rect 16309 51047 16355 51246
rect 16309 50944 16355 50955
rect 16066 50862 16432 50879
rect 16066 50816 16079 50862
rect 16125 50816 16373 50862
rect 16419 50816 16432 50862
rect 16066 50803 16432 50816
<< end >>
