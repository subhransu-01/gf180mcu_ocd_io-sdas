magic
tech gf180mcuD
magscale 1 10
timestamp 1764347740
<< nwell >>
rect 18130 54786 19237 55988
rect 18130 54691 19183 54786
<< hvnmos >>
rect 18491 53764 18631 54064
rect 18735 53764 18875 54064
<< hvpmos >>
rect 18491 55332 18631 55632
rect 18735 55332 18875 55632
<< mvndiff >>
rect 18403 54051 18491 54064
rect 18403 54005 18416 54051
rect 18462 54005 18491 54051
rect 18403 53937 18491 54005
rect 18403 53891 18416 53937
rect 18462 53891 18491 53937
rect 18403 53823 18491 53891
rect 18403 53777 18416 53823
rect 18462 53777 18491 53823
rect 18403 53764 18491 53777
rect 18631 54051 18735 54064
rect 18631 54005 18660 54051
rect 18706 54005 18735 54051
rect 18631 53937 18735 54005
rect 18631 53891 18660 53937
rect 18706 53891 18735 53937
rect 18631 53823 18735 53891
rect 18631 53777 18660 53823
rect 18706 53777 18735 53823
rect 18631 53764 18735 53777
rect 18875 54051 18965 54064
rect 18875 54005 18904 54051
rect 18950 54005 18965 54051
rect 18875 53937 18965 54005
rect 18875 53891 18904 53937
rect 18950 53891 18965 53937
rect 18875 53823 18965 53891
rect 18875 53777 18904 53823
rect 18950 53777 18965 53823
rect 18875 53764 18965 53777
<< mvpdiff >>
rect 18403 55619 18491 55632
rect 18403 55573 18416 55619
rect 18462 55573 18491 55619
rect 18403 55514 18491 55573
rect 18403 55468 18416 55514
rect 18462 55468 18491 55514
rect 18403 55409 18491 55468
rect 18403 55363 18416 55409
rect 18462 55363 18491 55409
rect 18403 55332 18491 55363
rect 18631 55619 18735 55632
rect 18631 55573 18660 55619
rect 18706 55573 18735 55619
rect 18631 55514 18735 55573
rect 18631 55468 18660 55514
rect 18706 55468 18735 55514
rect 18631 55409 18735 55468
rect 18631 55363 18660 55409
rect 18706 55363 18735 55409
rect 18631 55332 18735 55363
rect 18875 55619 18965 55632
rect 18875 55573 18904 55619
rect 18950 55573 18965 55619
rect 18875 55514 18965 55573
rect 18875 55468 18904 55514
rect 18950 55468 18965 55514
rect 18875 55409 18965 55468
rect 18875 55363 18904 55409
rect 18950 55363 18965 55409
rect 18875 55332 18965 55363
<< mvndiffc >>
rect 18416 54005 18462 54051
rect 18416 53891 18462 53937
rect 18416 53777 18462 53823
rect 18660 54005 18706 54051
rect 18660 53891 18706 53937
rect 18660 53777 18706 53823
rect 18904 54005 18950 54051
rect 18904 53891 18950 53937
rect 18904 53777 18950 53823
<< mvpdiffc >>
rect 18416 55573 18462 55619
rect 18416 55468 18462 55514
rect 18416 55363 18462 55409
rect 18660 55573 18706 55619
rect 18660 55468 18706 55514
rect 18660 55363 18706 55409
rect 18904 55573 18950 55619
rect 18904 55468 18950 55514
rect 18904 55363 18950 55409
<< psubdiff >>
rect 18216 54324 18306 54346
rect 18216 53432 18238 54324
rect 18284 53500 18306 54324
rect 19061 54418 19151 54440
rect 19061 53500 19083 54418
rect 18284 53478 19083 53500
rect 18284 53432 18369 53478
rect 18966 53432 19083 53478
rect 19129 53432 19151 54418
rect 18216 53410 19151 53432
<< nsubdiff >>
rect 18216 55880 19151 55902
rect 18216 54894 18238 55880
rect 18284 55834 18378 55880
rect 18977 55834 19083 55880
rect 18284 55812 19083 55834
rect 18284 54894 18306 55812
rect 18216 54872 18306 54894
rect 19061 54894 19083 55812
rect 19129 54894 19151 55880
rect 19061 54872 19151 54894
<< psubdiffcont >>
rect 18238 53432 18284 54324
rect 18369 53432 18966 53478
rect 19083 53432 19129 54418
<< nsubdiffcont >>
rect 18238 54894 18284 55880
rect 18378 55834 18977 55880
rect 19083 54894 19129 55880
<< polysilicon >>
rect 18491 55632 18631 55676
rect 18735 55632 18875 55676
rect 18491 55272 18631 55332
rect 18491 55257 18665 55272
rect 18491 55195 18537 55257
rect 18649 55195 18665 55257
rect 18491 55181 18665 55195
rect 18735 55130 18875 55332
rect 18505 55116 18875 55130
rect 18505 55056 18521 55116
rect 18724 55056 18875 55116
rect 18505 55040 18875 55056
rect 18481 54786 18875 54830
rect 18481 54687 18500 54786
rect 18621 54687 18875 54786
rect 18481 54667 18875 54687
rect 18479 54527 18631 54544
rect 18479 54420 18492 54527
rect 18616 54420 18631 54527
rect 18479 54386 18631 54420
rect 18491 54064 18631 54386
rect 18735 54064 18875 54667
rect 18491 53720 18631 53764
rect 18735 53720 18875 53764
<< polycontact >>
rect 18537 55195 18649 55257
rect 18521 55056 18724 55116
rect 18500 54687 18621 54786
rect 18492 54420 18616 54527
<< metal1 >>
rect 18227 55880 19144 55891
rect 18227 54894 18238 55880
rect 18284 55834 18378 55880
rect 18977 55834 19083 55880
rect 18284 55823 19083 55834
rect 18284 54894 18295 55823
rect 18401 55619 18477 55632
rect 18401 55573 18416 55619
rect 18462 55573 18477 55619
rect 18401 55514 18477 55573
rect 18401 55468 18416 55514
rect 18462 55468 18477 55514
rect 18401 55409 18477 55468
rect 18401 55363 18416 55409
rect 18462 55363 18477 55409
rect 18401 55129 18477 55363
rect 18645 55619 18722 55823
rect 18645 55573 18660 55619
rect 18706 55573 18722 55619
rect 18645 55514 18722 55573
rect 18645 55468 18660 55514
rect 18706 55468 18722 55514
rect 18645 55409 18722 55468
rect 18645 55363 18660 55409
rect 18706 55363 18722 55409
rect 18645 55328 18722 55363
rect 18889 55619 18965 55632
rect 18889 55573 18904 55619
rect 18950 55573 18965 55619
rect 18889 55514 18965 55573
rect 18889 55468 18904 55514
rect 18950 55468 18965 55514
rect 18889 55409 18965 55468
rect 18889 55363 18904 55409
rect 18950 55363 18965 55409
rect 18889 55272 18965 55363
rect 18524 55257 18965 55272
rect 18524 55195 18537 55257
rect 18649 55195 18965 55257
rect 18524 55178 18965 55195
rect 18401 55116 18782 55129
rect 18401 55056 18521 55116
rect 18724 55056 18782 55116
rect 18401 55043 18782 55056
rect 18227 54883 18295 54894
rect 18371 54786 18632 54820
rect 18371 54687 18500 54786
rect 18621 54687 18632 54786
rect 18371 54663 18632 54687
rect 18371 54527 18632 54543
rect 18371 54420 18492 54527
rect 18616 54420 18632 54527
rect 18371 54386 18632 54420
rect 18227 54324 18295 54335
rect 18227 53432 18238 54324
rect 18284 53489 18295 54324
rect 18706 54208 18782 55043
rect 18401 54132 18782 54208
rect 18401 54051 18477 54132
rect 18401 54005 18416 54051
rect 18462 54005 18477 54051
rect 18401 53937 18477 54005
rect 18401 53891 18416 53937
rect 18462 53891 18477 53937
rect 18401 53823 18477 53891
rect 18401 53777 18416 53823
rect 18462 53777 18477 53823
rect 18401 53764 18477 53777
rect 18645 54051 18720 54064
rect 18645 54005 18660 54051
rect 18706 54005 18720 54051
rect 18645 53937 18720 54005
rect 18645 53891 18660 53937
rect 18706 53891 18720 53937
rect 18645 53823 18720 53891
rect 18645 53777 18660 53823
rect 18706 53777 18720 53823
rect 18645 53489 18720 53777
rect 18889 54051 18965 55178
rect 19068 54894 19083 55823
rect 19129 54894 19144 55880
rect 19068 54883 19144 54894
rect 19072 54418 19140 54429
rect 19072 54329 19083 54418
rect 18889 54005 18904 54051
rect 18950 54005 18965 54051
rect 18889 53937 18965 54005
rect 18889 53891 18904 53937
rect 18950 53891 18965 53937
rect 18889 53823 18965 53891
rect 18889 53777 18904 53823
rect 18950 53777 18965 53823
rect 18889 53764 18965 53777
rect 19068 53489 19083 54329
rect 18284 53478 19083 53489
rect 18284 53432 18369 53478
rect 18966 53432 19083 53478
rect 19129 54329 19140 54418
rect 19129 53432 19144 54329
rect 18227 53421 19144 53432
<< end >>
