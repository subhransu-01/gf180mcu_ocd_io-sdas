magic
tech gf180mcuD
magscale 1 10
timestamp 1764272961
<< metal1 >>
rect -44 7953 200 8000
rect -44 7901 0 7953
rect 156 7901 200 7953
rect -44 7829 200 7901
rect -44 7777 0 7829
rect 156 7777 200 7829
rect -44 7705 200 7777
rect -44 7653 0 7705
rect 156 7653 200 7705
rect -44 7581 200 7653
rect -44 7529 0 7581
rect 156 7529 200 7581
rect -44 7457 200 7529
rect -44 7405 0 7457
rect 156 7405 200 7457
rect -44 7333 200 7405
rect -44 7281 0 7333
rect 156 7281 200 7333
rect -44 7209 200 7281
rect -44 7157 0 7209
rect 156 7157 200 7209
rect -44 7085 200 7157
rect -44 7033 0 7085
rect 156 7033 200 7085
rect -44 6961 200 7033
rect -44 6909 0 6961
rect 156 6909 200 6961
rect -44 6837 200 6909
rect -44 6785 0 6837
rect 156 6785 200 6837
rect -44 6713 200 6785
rect -44 6661 0 6713
rect 156 6661 200 6713
rect -44 6589 200 6661
rect -44 6537 0 6589
rect 156 6537 200 6589
rect -44 6465 200 6537
rect -44 6413 0 6465
rect 156 6413 200 6465
rect -44 6341 200 6413
rect -44 6289 0 6341
rect 156 6289 200 6341
rect -44 6217 200 6289
rect -44 6165 0 6217
rect 156 6165 200 6217
rect -44 6093 200 6165
rect -44 6041 0 6093
rect 156 6041 200 6093
rect -44 5969 200 6041
rect -44 5917 0 5969
rect 156 5917 200 5969
rect -44 5845 200 5917
rect -44 5793 0 5845
rect 156 5793 200 5845
rect -44 5721 200 5793
rect -44 5669 0 5721
rect 156 5669 200 5721
rect -44 5597 200 5669
rect -44 5545 0 5597
rect 156 5545 200 5597
rect -44 5473 200 5545
rect -44 5421 0 5473
rect 156 5421 200 5473
rect -44 5349 200 5421
rect -44 5297 0 5349
rect 156 5297 200 5349
rect -44 5225 200 5297
rect -44 5173 0 5225
rect 156 5173 200 5225
rect -44 5101 200 5173
rect -44 5049 0 5101
rect 156 5049 200 5101
rect -44 4977 200 5049
rect -44 4925 0 4977
rect 156 4925 200 4977
rect -44 4853 200 4925
rect -44 4801 0 4853
rect 156 4801 200 4853
rect -44 4729 200 4801
rect -44 4677 0 4729
rect 156 4677 200 4729
rect -44 4605 200 4677
rect -44 4553 0 4605
rect 156 4553 200 4605
rect -44 4481 200 4553
rect -44 4429 0 4481
rect 156 4429 200 4481
rect -44 4357 200 4429
rect -44 4305 0 4357
rect 156 4305 200 4357
rect -44 4233 200 4305
rect -44 4181 0 4233
rect 156 4181 200 4233
rect -44 4109 200 4181
rect -44 4057 0 4109
rect 156 4057 200 4109
rect -44 3985 200 4057
rect -44 3933 0 3985
rect 156 3933 200 3985
rect -44 3861 200 3933
rect -44 3809 0 3861
rect 156 3809 200 3861
rect -44 3737 200 3809
rect -44 3685 0 3737
rect 156 3685 200 3737
rect -44 3613 200 3685
rect -44 3561 0 3613
rect 156 3561 200 3613
rect -44 3489 200 3561
rect -44 3437 0 3489
rect 156 3437 200 3489
rect -44 3365 200 3437
rect -44 3313 0 3365
rect 156 3313 200 3365
rect -44 3241 200 3313
rect -44 3189 0 3241
rect 156 3189 200 3241
rect -44 3117 200 3189
rect -44 3065 0 3117
rect 156 3065 200 3117
rect -44 2993 200 3065
rect -44 2941 0 2993
rect 156 2941 200 2993
rect -44 2869 200 2941
rect -44 2817 0 2869
rect 156 2817 200 2869
rect -44 2745 200 2817
rect -44 2693 0 2745
rect 156 2693 200 2745
rect -44 2621 200 2693
rect -44 2569 0 2621
rect 156 2569 200 2621
rect -44 2497 200 2569
rect -44 2445 0 2497
rect 156 2445 200 2497
rect -44 2373 200 2445
rect -44 2321 0 2373
rect 156 2321 200 2373
rect -44 2249 200 2321
rect -44 2197 0 2249
rect 156 2197 200 2249
rect -44 2125 200 2197
rect -44 2073 0 2125
rect 156 2073 200 2125
rect -44 2001 200 2073
rect -44 1949 0 2001
rect 156 1949 200 2001
rect -44 1877 200 1949
rect -44 1825 0 1877
rect 156 1825 200 1877
rect -44 1753 200 1825
rect -44 1701 0 1753
rect 156 1701 200 1753
rect -44 1629 200 1701
rect -44 1577 0 1629
rect 156 1577 200 1629
rect -44 1505 200 1577
rect -44 1453 0 1505
rect 156 1453 200 1505
rect -44 1381 200 1453
rect -44 1329 0 1381
rect 156 1329 200 1381
rect -44 1257 200 1329
rect -44 1205 0 1257
rect 156 1205 200 1257
rect -44 1133 200 1205
rect -44 1081 0 1133
rect 156 1081 200 1133
rect -44 1009 200 1081
rect -44 957 0 1009
rect 156 957 200 1009
rect -44 885 200 957
rect -44 833 0 885
rect 156 833 200 885
rect -44 761 200 833
rect -44 709 0 761
rect 156 709 200 761
rect -44 637 200 709
rect -44 585 0 637
rect 156 585 200 637
rect -44 513 200 585
rect -44 461 0 513
rect 156 461 200 513
rect -44 400 200 461
rect 430 7945 2074 8000
rect 430 7893 482 7945
rect 534 7893 606 7945
rect 658 7893 730 7945
rect 782 7893 854 7945
rect 906 7893 978 7945
rect 1030 7893 1102 7945
rect 1154 7893 1226 7945
rect 1278 7893 1350 7945
rect 1402 7893 1474 7945
rect 1526 7893 1598 7945
rect 1650 7893 1722 7945
rect 1774 7893 1846 7945
rect 1898 7893 1970 7945
rect 2022 7893 2074 7945
rect 430 7821 2074 7893
rect 430 7769 482 7821
rect 534 7769 606 7821
rect 658 7769 730 7821
rect 782 7769 854 7821
rect 906 7769 978 7821
rect 1030 7769 1102 7821
rect 1154 7769 1226 7821
rect 1278 7769 1350 7821
rect 1402 7769 1474 7821
rect 1526 7769 1598 7821
rect 1650 7769 1722 7821
rect 1774 7769 1846 7821
rect 1898 7769 1970 7821
rect 2022 7769 2074 7821
rect 430 7697 2074 7769
rect 430 7645 482 7697
rect 534 7645 606 7697
rect 658 7645 730 7697
rect 782 7645 854 7697
rect 906 7645 978 7697
rect 1030 7645 1102 7697
rect 1154 7645 1226 7697
rect 1278 7645 1350 7697
rect 1402 7645 1474 7697
rect 1526 7645 1598 7697
rect 1650 7645 1722 7697
rect 1774 7645 1846 7697
rect 1898 7645 1970 7697
rect 2022 7645 2074 7697
rect 430 7573 2074 7645
rect 430 7521 482 7573
rect 534 7521 606 7573
rect 658 7521 730 7573
rect 782 7521 854 7573
rect 906 7521 978 7573
rect 1030 7521 1102 7573
rect 1154 7521 1226 7573
rect 1278 7521 1350 7573
rect 1402 7521 1474 7573
rect 1526 7521 1598 7573
rect 1650 7521 1722 7573
rect 1774 7521 1846 7573
rect 1898 7521 1970 7573
rect 2022 7521 2074 7573
rect 430 7449 2074 7521
rect 430 7397 482 7449
rect 534 7397 606 7449
rect 658 7397 730 7449
rect 782 7397 854 7449
rect 906 7397 978 7449
rect 1030 7397 1102 7449
rect 1154 7397 1226 7449
rect 1278 7397 1350 7449
rect 1402 7397 1474 7449
rect 1526 7397 1598 7449
rect 1650 7397 1722 7449
rect 1774 7397 1846 7449
rect 1898 7397 1970 7449
rect 2022 7397 2074 7449
rect 430 7325 2074 7397
rect 430 7273 482 7325
rect 534 7273 606 7325
rect 658 7273 730 7325
rect 782 7273 854 7325
rect 906 7273 978 7325
rect 1030 7273 1102 7325
rect 1154 7273 1226 7325
rect 1278 7273 1350 7325
rect 1402 7273 1474 7325
rect 1526 7273 1598 7325
rect 1650 7273 1722 7325
rect 1774 7273 1846 7325
rect 1898 7273 1970 7325
rect 2022 7273 2074 7325
rect 430 7201 2074 7273
rect 430 7149 482 7201
rect 534 7149 606 7201
rect 658 7149 730 7201
rect 782 7149 854 7201
rect 906 7149 978 7201
rect 1030 7149 1102 7201
rect 1154 7149 1226 7201
rect 1278 7149 1350 7201
rect 1402 7149 1474 7201
rect 1526 7149 1598 7201
rect 1650 7149 1722 7201
rect 1774 7149 1846 7201
rect 1898 7149 1970 7201
rect 2022 7149 2074 7201
rect 430 7077 2074 7149
rect 430 7025 482 7077
rect 534 7025 606 7077
rect 658 7025 730 7077
rect 782 7025 854 7077
rect 906 7025 978 7077
rect 1030 7025 1102 7077
rect 1154 7025 1226 7077
rect 1278 7025 1350 7077
rect 1402 7025 1474 7077
rect 1526 7025 1598 7077
rect 1650 7025 1722 7077
rect 1774 7025 1846 7077
rect 1898 7025 1970 7077
rect 2022 7025 2074 7077
rect 430 6953 2074 7025
rect 430 6901 482 6953
rect 534 6901 606 6953
rect 658 6901 730 6953
rect 782 6901 854 6953
rect 906 6901 978 6953
rect 1030 6901 1102 6953
rect 1154 6901 1226 6953
rect 1278 6901 1350 6953
rect 1402 6901 1474 6953
rect 1526 6901 1598 6953
rect 1650 6901 1722 6953
rect 1774 6901 1846 6953
rect 1898 6901 1970 6953
rect 2022 6901 2074 6953
rect 430 6829 2074 6901
rect 430 6777 482 6829
rect 534 6777 606 6829
rect 658 6777 730 6829
rect 782 6777 854 6829
rect 906 6777 978 6829
rect 1030 6777 1102 6829
rect 1154 6777 1226 6829
rect 1278 6777 1350 6829
rect 1402 6777 1474 6829
rect 1526 6777 1598 6829
rect 1650 6777 1722 6829
rect 1774 6777 1846 6829
rect 1898 6777 1970 6829
rect 2022 6777 2074 6829
rect 430 6705 2074 6777
rect 430 6653 482 6705
rect 534 6653 606 6705
rect 658 6653 730 6705
rect 782 6653 854 6705
rect 906 6653 978 6705
rect 1030 6653 1102 6705
rect 1154 6653 1226 6705
rect 1278 6653 1350 6705
rect 1402 6653 1474 6705
rect 1526 6653 1598 6705
rect 1650 6653 1722 6705
rect 1774 6653 1846 6705
rect 1898 6653 1970 6705
rect 2022 6653 2074 6705
rect 430 6581 2074 6653
rect 430 6529 482 6581
rect 534 6529 606 6581
rect 658 6529 730 6581
rect 782 6529 854 6581
rect 906 6529 978 6581
rect 1030 6529 1102 6581
rect 1154 6529 1226 6581
rect 1278 6529 1350 6581
rect 1402 6529 1474 6581
rect 1526 6529 1598 6581
rect 1650 6529 1722 6581
rect 1774 6529 1846 6581
rect 1898 6529 1970 6581
rect 2022 6529 2074 6581
rect 430 6457 2074 6529
rect 430 6405 482 6457
rect 534 6405 606 6457
rect 658 6405 730 6457
rect 782 6405 854 6457
rect 906 6405 978 6457
rect 1030 6405 1102 6457
rect 1154 6405 1226 6457
rect 1278 6405 1350 6457
rect 1402 6405 1474 6457
rect 1526 6405 1598 6457
rect 1650 6405 1722 6457
rect 1774 6405 1846 6457
rect 1898 6405 1970 6457
rect 2022 6405 2074 6457
rect 430 6333 2074 6405
rect 430 6281 482 6333
rect 534 6281 606 6333
rect 658 6281 730 6333
rect 782 6281 854 6333
rect 906 6281 978 6333
rect 1030 6281 1102 6333
rect 1154 6281 1226 6333
rect 1278 6281 1350 6333
rect 1402 6281 1474 6333
rect 1526 6281 1598 6333
rect 1650 6281 1722 6333
rect 1774 6281 1846 6333
rect 1898 6281 1970 6333
rect 2022 6281 2074 6333
rect 430 6209 2074 6281
rect 430 6157 482 6209
rect 534 6157 606 6209
rect 658 6157 730 6209
rect 782 6157 854 6209
rect 906 6157 978 6209
rect 1030 6157 1102 6209
rect 1154 6157 1226 6209
rect 1278 6157 1350 6209
rect 1402 6157 1474 6209
rect 1526 6157 1598 6209
rect 1650 6157 1722 6209
rect 1774 6157 1846 6209
rect 1898 6157 1970 6209
rect 2022 6157 2074 6209
rect 430 6085 2074 6157
rect 430 6033 482 6085
rect 534 6033 606 6085
rect 658 6033 730 6085
rect 782 6033 854 6085
rect 906 6033 978 6085
rect 1030 6033 1102 6085
rect 1154 6033 1226 6085
rect 1278 6033 1350 6085
rect 1402 6033 1474 6085
rect 1526 6033 1598 6085
rect 1650 6033 1722 6085
rect 1774 6033 1846 6085
rect 1898 6033 1970 6085
rect 2022 6033 2074 6085
rect 430 5961 2074 6033
rect 430 5909 482 5961
rect 534 5909 606 5961
rect 658 5909 730 5961
rect 782 5909 854 5961
rect 906 5909 978 5961
rect 1030 5909 1102 5961
rect 1154 5909 1226 5961
rect 1278 5909 1350 5961
rect 1402 5909 1474 5961
rect 1526 5909 1598 5961
rect 1650 5909 1722 5961
rect 1774 5909 1846 5961
rect 1898 5909 1970 5961
rect 2022 5909 2074 5961
rect 430 5837 2074 5909
rect 430 5785 482 5837
rect 534 5785 606 5837
rect 658 5785 730 5837
rect 782 5785 854 5837
rect 906 5785 978 5837
rect 1030 5785 1102 5837
rect 1154 5785 1226 5837
rect 1278 5785 1350 5837
rect 1402 5785 1474 5837
rect 1526 5785 1598 5837
rect 1650 5785 1722 5837
rect 1774 5785 1846 5837
rect 1898 5785 1970 5837
rect 2022 5785 2074 5837
rect 430 5713 2074 5785
rect 430 5661 482 5713
rect 534 5661 606 5713
rect 658 5661 730 5713
rect 782 5661 854 5713
rect 906 5661 978 5713
rect 1030 5661 1102 5713
rect 1154 5661 1226 5713
rect 1278 5661 1350 5713
rect 1402 5661 1474 5713
rect 1526 5661 1598 5713
rect 1650 5661 1722 5713
rect 1774 5661 1846 5713
rect 1898 5661 1970 5713
rect 2022 5661 2074 5713
rect 430 5589 2074 5661
rect 430 5537 482 5589
rect 534 5537 606 5589
rect 658 5537 730 5589
rect 782 5537 854 5589
rect 906 5537 978 5589
rect 1030 5537 1102 5589
rect 1154 5537 1226 5589
rect 1278 5537 1350 5589
rect 1402 5537 1474 5589
rect 1526 5537 1598 5589
rect 1650 5537 1722 5589
rect 1774 5537 1846 5589
rect 1898 5537 1970 5589
rect 2022 5537 2074 5589
rect 430 5465 2074 5537
rect 430 5413 482 5465
rect 534 5413 606 5465
rect 658 5413 730 5465
rect 782 5413 854 5465
rect 906 5413 978 5465
rect 1030 5413 1102 5465
rect 1154 5413 1226 5465
rect 1278 5413 1350 5465
rect 1402 5413 1474 5465
rect 1526 5413 1598 5465
rect 1650 5413 1722 5465
rect 1774 5413 1846 5465
rect 1898 5413 1970 5465
rect 2022 5413 2074 5465
rect 430 5341 2074 5413
rect 430 5289 482 5341
rect 534 5289 606 5341
rect 658 5289 730 5341
rect 782 5289 854 5341
rect 906 5289 978 5341
rect 1030 5289 1102 5341
rect 1154 5289 1226 5341
rect 1278 5289 1350 5341
rect 1402 5289 1474 5341
rect 1526 5289 1598 5341
rect 1650 5289 1722 5341
rect 1774 5289 1846 5341
rect 1898 5289 1970 5341
rect 2022 5289 2074 5341
rect 430 5217 2074 5289
rect 430 5165 482 5217
rect 534 5165 606 5217
rect 658 5165 730 5217
rect 782 5165 854 5217
rect 906 5165 978 5217
rect 1030 5165 1102 5217
rect 1154 5165 1226 5217
rect 1278 5165 1350 5217
rect 1402 5165 1474 5217
rect 1526 5165 1598 5217
rect 1650 5165 1722 5217
rect 1774 5165 1846 5217
rect 1898 5165 1970 5217
rect 2022 5165 2074 5217
rect 430 5093 2074 5165
rect 430 5041 482 5093
rect 534 5041 606 5093
rect 658 5041 730 5093
rect 782 5041 854 5093
rect 906 5041 978 5093
rect 1030 5041 1102 5093
rect 1154 5041 1226 5093
rect 1278 5041 1350 5093
rect 1402 5041 1474 5093
rect 1526 5041 1598 5093
rect 1650 5041 1722 5093
rect 1774 5041 1846 5093
rect 1898 5041 1970 5093
rect 2022 5041 2074 5093
rect 430 4969 2074 5041
rect 430 4917 482 4969
rect 534 4917 606 4969
rect 658 4917 730 4969
rect 782 4917 854 4969
rect 906 4917 978 4969
rect 1030 4917 1102 4969
rect 1154 4917 1226 4969
rect 1278 4917 1350 4969
rect 1402 4917 1474 4969
rect 1526 4917 1598 4969
rect 1650 4917 1722 4969
rect 1774 4917 1846 4969
rect 1898 4917 1970 4969
rect 2022 4917 2074 4969
rect 430 4845 2074 4917
rect 430 4793 482 4845
rect 534 4793 606 4845
rect 658 4793 730 4845
rect 782 4793 854 4845
rect 906 4793 978 4845
rect 1030 4793 1102 4845
rect 1154 4793 1226 4845
rect 1278 4793 1350 4845
rect 1402 4793 1474 4845
rect 1526 4793 1598 4845
rect 1650 4793 1722 4845
rect 1774 4793 1846 4845
rect 1898 4793 1970 4845
rect 2022 4793 2074 4845
rect 430 4721 2074 4793
rect 430 4669 482 4721
rect 534 4669 606 4721
rect 658 4669 730 4721
rect 782 4669 854 4721
rect 906 4669 978 4721
rect 1030 4669 1102 4721
rect 1154 4669 1226 4721
rect 1278 4669 1350 4721
rect 1402 4669 1474 4721
rect 1526 4669 1598 4721
rect 1650 4669 1722 4721
rect 1774 4669 1846 4721
rect 1898 4669 1970 4721
rect 2022 4669 2074 4721
rect 430 4597 2074 4669
rect 430 4545 482 4597
rect 534 4545 606 4597
rect 658 4545 730 4597
rect 782 4545 854 4597
rect 906 4545 978 4597
rect 1030 4545 1102 4597
rect 1154 4545 1226 4597
rect 1278 4545 1350 4597
rect 1402 4545 1474 4597
rect 1526 4545 1598 4597
rect 1650 4545 1722 4597
rect 1774 4545 1846 4597
rect 1898 4545 1970 4597
rect 2022 4545 2074 4597
rect 430 4473 2074 4545
rect 430 4421 482 4473
rect 534 4421 606 4473
rect 658 4421 730 4473
rect 782 4421 854 4473
rect 906 4421 978 4473
rect 1030 4421 1102 4473
rect 1154 4421 1226 4473
rect 1278 4421 1350 4473
rect 1402 4421 1474 4473
rect 1526 4421 1598 4473
rect 1650 4421 1722 4473
rect 1774 4421 1846 4473
rect 1898 4421 1970 4473
rect 2022 4421 2074 4473
rect 430 4349 2074 4421
rect 430 4297 482 4349
rect 534 4297 606 4349
rect 658 4297 730 4349
rect 782 4297 854 4349
rect 906 4297 978 4349
rect 1030 4297 1102 4349
rect 1154 4297 1226 4349
rect 1278 4297 1350 4349
rect 1402 4297 1474 4349
rect 1526 4297 1598 4349
rect 1650 4297 1722 4349
rect 1774 4297 1846 4349
rect 1898 4297 1970 4349
rect 2022 4297 2074 4349
rect 430 4225 2074 4297
rect 430 4173 482 4225
rect 534 4173 606 4225
rect 658 4173 730 4225
rect 782 4173 854 4225
rect 906 4173 978 4225
rect 1030 4173 1102 4225
rect 1154 4173 1226 4225
rect 1278 4173 1350 4225
rect 1402 4173 1474 4225
rect 1526 4173 1598 4225
rect 1650 4173 1722 4225
rect 1774 4173 1846 4225
rect 1898 4173 1970 4225
rect 2022 4173 2074 4225
rect 430 4101 2074 4173
rect 430 4049 482 4101
rect 534 4049 606 4101
rect 658 4049 730 4101
rect 782 4049 854 4101
rect 906 4049 978 4101
rect 1030 4049 1102 4101
rect 1154 4049 1226 4101
rect 1278 4049 1350 4101
rect 1402 4049 1474 4101
rect 1526 4049 1598 4101
rect 1650 4049 1722 4101
rect 1774 4049 1846 4101
rect 1898 4049 1970 4101
rect 2022 4049 2074 4101
rect 430 3977 2074 4049
rect 430 3925 482 3977
rect 534 3925 606 3977
rect 658 3925 730 3977
rect 782 3925 854 3977
rect 906 3925 978 3977
rect 1030 3925 1102 3977
rect 1154 3925 1226 3977
rect 1278 3925 1350 3977
rect 1402 3925 1474 3977
rect 1526 3925 1598 3977
rect 1650 3925 1722 3977
rect 1774 3925 1846 3977
rect 1898 3925 1970 3977
rect 2022 3925 2074 3977
rect 430 3853 2074 3925
rect 430 3801 482 3853
rect 534 3801 606 3853
rect 658 3801 730 3853
rect 782 3801 854 3853
rect 906 3801 978 3853
rect 1030 3801 1102 3853
rect 1154 3801 1226 3853
rect 1278 3801 1350 3853
rect 1402 3801 1474 3853
rect 1526 3801 1598 3853
rect 1650 3801 1722 3853
rect 1774 3801 1846 3853
rect 1898 3801 1970 3853
rect 2022 3801 2074 3853
rect 430 3729 2074 3801
rect 430 3677 482 3729
rect 534 3677 606 3729
rect 658 3677 730 3729
rect 782 3677 854 3729
rect 906 3677 978 3729
rect 1030 3677 1102 3729
rect 1154 3677 1226 3729
rect 1278 3677 1350 3729
rect 1402 3677 1474 3729
rect 1526 3677 1598 3729
rect 1650 3677 1722 3729
rect 1774 3677 1846 3729
rect 1898 3677 1970 3729
rect 2022 3677 2074 3729
rect 430 3605 2074 3677
rect 430 3553 482 3605
rect 534 3553 606 3605
rect 658 3553 730 3605
rect 782 3553 854 3605
rect 906 3553 978 3605
rect 1030 3553 1102 3605
rect 1154 3553 1226 3605
rect 1278 3553 1350 3605
rect 1402 3553 1474 3605
rect 1526 3553 1598 3605
rect 1650 3553 1722 3605
rect 1774 3553 1846 3605
rect 1898 3553 1970 3605
rect 2022 3553 2074 3605
rect 430 3481 2074 3553
rect 430 3429 482 3481
rect 534 3429 606 3481
rect 658 3429 730 3481
rect 782 3429 854 3481
rect 906 3429 978 3481
rect 1030 3429 1102 3481
rect 1154 3429 1226 3481
rect 1278 3429 1350 3481
rect 1402 3429 1474 3481
rect 1526 3429 1598 3481
rect 1650 3429 1722 3481
rect 1774 3429 1846 3481
rect 1898 3429 1970 3481
rect 2022 3429 2074 3481
rect 430 3357 2074 3429
rect 430 3305 482 3357
rect 534 3305 606 3357
rect 658 3305 730 3357
rect 782 3305 854 3357
rect 906 3305 978 3357
rect 1030 3305 1102 3357
rect 1154 3305 1226 3357
rect 1278 3305 1350 3357
rect 1402 3305 1474 3357
rect 1526 3305 1598 3357
rect 1650 3305 1722 3357
rect 1774 3305 1846 3357
rect 1898 3305 1970 3357
rect 2022 3305 2074 3357
rect 430 3233 2074 3305
rect 430 3181 482 3233
rect 534 3181 606 3233
rect 658 3181 730 3233
rect 782 3181 854 3233
rect 906 3181 978 3233
rect 1030 3181 1102 3233
rect 1154 3181 1226 3233
rect 1278 3181 1350 3233
rect 1402 3181 1474 3233
rect 1526 3181 1598 3233
rect 1650 3181 1722 3233
rect 1774 3181 1846 3233
rect 1898 3181 1970 3233
rect 2022 3181 2074 3233
rect 430 3109 2074 3181
rect 430 3057 482 3109
rect 534 3057 606 3109
rect 658 3057 730 3109
rect 782 3057 854 3109
rect 906 3057 978 3109
rect 1030 3057 1102 3109
rect 1154 3057 1226 3109
rect 1278 3057 1350 3109
rect 1402 3057 1474 3109
rect 1526 3057 1598 3109
rect 1650 3057 1722 3109
rect 1774 3057 1846 3109
rect 1898 3057 1970 3109
rect 2022 3057 2074 3109
rect 430 2985 2074 3057
rect 430 2933 482 2985
rect 534 2933 606 2985
rect 658 2933 730 2985
rect 782 2933 854 2985
rect 906 2933 978 2985
rect 1030 2933 1102 2985
rect 1154 2933 1226 2985
rect 1278 2933 1350 2985
rect 1402 2933 1474 2985
rect 1526 2933 1598 2985
rect 1650 2933 1722 2985
rect 1774 2933 1846 2985
rect 1898 2933 1970 2985
rect 2022 2933 2074 2985
rect 430 2861 2074 2933
rect 430 2809 482 2861
rect 534 2809 606 2861
rect 658 2809 730 2861
rect 782 2809 854 2861
rect 906 2809 978 2861
rect 1030 2809 1102 2861
rect 1154 2809 1226 2861
rect 1278 2809 1350 2861
rect 1402 2809 1474 2861
rect 1526 2809 1598 2861
rect 1650 2809 1722 2861
rect 1774 2809 1846 2861
rect 1898 2809 1970 2861
rect 2022 2809 2074 2861
rect 430 2737 2074 2809
rect 430 2685 482 2737
rect 534 2685 606 2737
rect 658 2685 730 2737
rect 782 2685 854 2737
rect 906 2685 978 2737
rect 1030 2685 1102 2737
rect 1154 2685 1226 2737
rect 1278 2685 1350 2737
rect 1402 2685 1474 2737
rect 1526 2685 1598 2737
rect 1650 2685 1722 2737
rect 1774 2685 1846 2737
rect 1898 2685 1970 2737
rect 2022 2685 2074 2737
rect 430 2613 2074 2685
rect 430 2561 482 2613
rect 534 2561 606 2613
rect 658 2561 730 2613
rect 782 2561 854 2613
rect 906 2561 978 2613
rect 1030 2561 1102 2613
rect 1154 2561 1226 2613
rect 1278 2561 1350 2613
rect 1402 2561 1474 2613
rect 1526 2561 1598 2613
rect 1650 2561 1722 2613
rect 1774 2561 1846 2613
rect 1898 2561 1970 2613
rect 2022 2561 2074 2613
rect 430 2489 2074 2561
rect 430 2437 482 2489
rect 534 2437 606 2489
rect 658 2437 730 2489
rect 782 2437 854 2489
rect 906 2437 978 2489
rect 1030 2437 1102 2489
rect 1154 2437 1226 2489
rect 1278 2437 1350 2489
rect 1402 2437 1474 2489
rect 1526 2437 1598 2489
rect 1650 2437 1722 2489
rect 1774 2437 1846 2489
rect 1898 2437 1970 2489
rect 2022 2437 2074 2489
rect 430 2365 2074 2437
rect 430 2313 482 2365
rect 534 2313 606 2365
rect 658 2313 730 2365
rect 782 2313 854 2365
rect 906 2313 978 2365
rect 1030 2313 1102 2365
rect 1154 2313 1226 2365
rect 1278 2313 1350 2365
rect 1402 2313 1474 2365
rect 1526 2313 1598 2365
rect 1650 2313 1722 2365
rect 1774 2313 1846 2365
rect 1898 2313 1970 2365
rect 2022 2313 2074 2365
rect 430 2241 2074 2313
rect 430 2189 482 2241
rect 534 2189 606 2241
rect 658 2189 730 2241
rect 782 2189 854 2241
rect 906 2189 978 2241
rect 1030 2189 1102 2241
rect 1154 2189 1226 2241
rect 1278 2189 1350 2241
rect 1402 2189 1474 2241
rect 1526 2189 1598 2241
rect 1650 2189 1722 2241
rect 1774 2189 1846 2241
rect 1898 2189 1970 2241
rect 2022 2189 2074 2241
rect 430 2117 2074 2189
rect 430 2065 482 2117
rect 534 2065 606 2117
rect 658 2065 730 2117
rect 782 2065 854 2117
rect 906 2065 978 2117
rect 1030 2065 1102 2117
rect 1154 2065 1226 2117
rect 1278 2065 1350 2117
rect 1402 2065 1474 2117
rect 1526 2065 1598 2117
rect 1650 2065 1722 2117
rect 1774 2065 1846 2117
rect 1898 2065 1970 2117
rect 2022 2065 2074 2117
rect 430 1993 2074 2065
rect 430 1941 482 1993
rect 534 1941 606 1993
rect 658 1941 730 1993
rect 782 1941 854 1993
rect 906 1941 978 1993
rect 1030 1941 1102 1993
rect 1154 1941 1226 1993
rect 1278 1941 1350 1993
rect 1402 1941 1474 1993
rect 1526 1941 1598 1993
rect 1650 1941 1722 1993
rect 1774 1941 1846 1993
rect 1898 1941 1970 1993
rect 2022 1941 2074 1993
rect 430 1869 2074 1941
rect 430 1817 482 1869
rect 534 1817 606 1869
rect 658 1817 730 1869
rect 782 1817 854 1869
rect 906 1817 978 1869
rect 1030 1817 1102 1869
rect 1154 1817 1226 1869
rect 1278 1817 1350 1869
rect 1402 1817 1474 1869
rect 1526 1817 1598 1869
rect 1650 1817 1722 1869
rect 1774 1817 1846 1869
rect 1898 1817 1970 1869
rect 2022 1817 2074 1869
rect 430 1745 2074 1817
rect 430 1693 482 1745
rect 534 1693 606 1745
rect 658 1693 730 1745
rect 782 1693 854 1745
rect 906 1693 978 1745
rect 1030 1693 1102 1745
rect 1154 1693 1226 1745
rect 1278 1693 1350 1745
rect 1402 1693 1474 1745
rect 1526 1693 1598 1745
rect 1650 1693 1722 1745
rect 1774 1693 1846 1745
rect 1898 1693 1970 1745
rect 2022 1693 2074 1745
rect 430 1621 2074 1693
rect 430 1569 482 1621
rect 534 1569 606 1621
rect 658 1569 730 1621
rect 782 1569 854 1621
rect 906 1569 978 1621
rect 1030 1569 1102 1621
rect 1154 1569 1226 1621
rect 1278 1569 1350 1621
rect 1402 1569 1474 1621
rect 1526 1569 1598 1621
rect 1650 1569 1722 1621
rect 1774 1569 1846 1621
rect 1898 1569 1970 1621
rect 2022 1569 2074 1621
rect 430 1497 2074 1569
rect 430 1445 482 1497
rect 534 1445 606 1497
rect 658 1445 730 1497
rect 782 1445 854 1497
rect 906 1445 978 1497
rect 1030 1445 1102 1497
rect 1154 1445 1226 1497
rect 1278 1445 1350 1497
rect 1402 1445 1474 1497
rect 1526 1445 1598 1497
rect 1650 1445 1722 1497
rect 1774 1445 1846 1497
rect 1898 1445 1970 1497
rect 2022 1445 2074 1497
rect 430 1373 2074 1445
rect 430 1321 482 1373
rect 534 1321 606 1373
rect 658 1321 730 1373
rect 782 1321 854 1373
rect 906 1321 978 1373
rect 1030 1321 1102 1373
rect 1154 1321 1226 1373
rect 1278 1321 1350 1373
rect 1402 1321 1474 1373
rect 1526 1321 1598 1373
rect 1650 1321 1722 1373
rect 1774 1321 1846 1373
rect 1898 1321 1970 1373
rect 2022 1321 2074 1373
rect 430 1249 2074 1321
rect 430 1197 482 1249
rect 534 1197 606 1249
rect 658 1197 730 1249
rect 782 1197 854 1249
rect 906 1197 978 1249
rect 1030 1197 1102 1249
rect 1154 1197 1226 1249
rect 1278 1197 1350 1249
rect 1402 1197 1474 1249
rect 1526 1197 1598 1249
rect 1650 1197 1722 1249
rect 1774 1197 1846 1249
rect 1898 1197 1970 1249
rect 2022 1197 2074 1249
rect 430 1125 2074 1197
rect 430 1073 482 1125
rect 534 1073 606 1125
rect 658 1073 730 1125
rect 782 1073 854 1125
rect 906 1073 978 1125
rect 1030 1073 1102 1125
rect 1154 1073 1226 1125
rect 1278 1073 1350 1125
rect 1402 1073 1474 1125
rect 1526 1073 1598 1125
rect 1650 1073 1722 1125
rect 1774 1073 1846 1125
rect 1898 1073 1970 1125
rect 2022 1073 2074 1125
rect 430 1001 2074 1073
rect 430 949 482 1001
rect 534 949 606 1001
rect 658 949 730 1001
rect 782 949 854 1001
rect 906 949 978 1001
rect 1030 949 1102 1001
rect 1154 949 1226 1001
rect 1278 949 1350 1001
rect 1402 949 1474 1001
rect 1526 949 1598 1001
rect 1650 949 1722 1001
rect 1774 949 1846 1001
rect 1898 949 1970 1001
rect 2022 949 2074 1001
rect 430 877 2074 949
rect 430 825 482 877
rect 534 825 606 877
rect 658 825 730 877
rect 782 825 854 877
rect 906 825 978 877
rect 1030 825 1102 877
rect 1154 825 1226 877
rect 1278 825 1350 877
rect 1402 825 1474 877
rect 1526 825 1598 877
rect 1650 825 1722 877
rect 1774 825 1846 877
rect 1898 825 1970 877
rect 2022 825 2074 877
rect 430 753 2074 825
rect 430 701 482 753
rect 534 701 606 753
rect 658 701 730 753
rect 782 701 854 753
rect 906 701 978 753
rect 1030 701 1102 753
rect 1154 701 1226 753
rect 1278 701 1350 753
rect 1402 701 1474 753
rect 1526 701 1598 753
rect 1650 701 1722 753
rect 1774 701 1846 753
rect 1898 701 1970 753
rect 2022 701 2074 753
rect 430 629 2074 701
rect 430 577 482 629
rect 534 577 606 629
rect 658 577 730 629
rect 782 577 854 629
rect 906 577 978 629
rect 1030 577 1102 629
rect 1154 577 1226 629
rect 1278 577 1350 629
rect 1402 577 1474 629
rect 1526 577 1598 629
rect 1650 577 1722 629
rect 1774 577 1846 629
rect 1898 577 1970 629
rect 2022 577 2074 629
rect 430 505 2074 577
rect 430 453 482 505
rect 534 453 606 505
rect 658 453 730 505
rect 782 453 854 505
rect 906 453 978 505
rect 1030 453 1102 505
rect 1154 453 1226 505
rect 1278 453 1350 505
rect 1402 453 1474 505
rect 1526 453 1598 505
rect 1650 453 1722 505
rect 1774 453 1846 505
rect 1898 453 1970 505
rect 2022 453 2074 505
rect 430 401 2074 453
<< via1 >>
rect 0 7901 156 7953
rect 0 7777 156 7829
rect 0 7653 156 7705
rect 0 7529 156 7581
rect 0 7405 156 7457
rect 0 7281 156 7333
rect 0 7157 156 7209
rect 0 7033 156 7085
rect 0 6909 156 6961
rect 0 6785 156 6837
rect 0 6661 156 6713
rect 0 6537 156 6589
rect 0 6413 156 6465
rect 0 6289 156 6341
rect 0 6165 156 6217
rect 0 6041 156 6093
rect 0 5917 156 5969
rect 0 5793 156 5845
rect 0 5669 156 5721
rect 0 5545 156 5597
rect 0 5421 156 5473
rect 0 5297 156 5349
rect 0 5173 156 5225
rect 0 5049 156 5101
rect 0 4925 156 4977
rect 0 4801 156 4853
rect 0 4677 156 4729
rect 0 4553 156 4605
rect 0 4429 156 4481
rect 0 4305 156 4357
rect 0 4181 156 4233
rect 0 4057 156 4109
rect 0 3933 156 3985
rect 0 3809 156 3861
rect 0 3685 156 3737
rect 0 3561 156 3613
rect 0 3437 156 3489
rect 0 3313 156 3365
rect 0 3189 156 3241
rect 0 3065 156 3117
rect 0 2941 156 2993
rect 0 2817 156 2869
rect 0 2693 156 2745
rect 0 2569 156 2621
rect 0 2445 156 2497
rect 0 2321 156 2373
rect 0 2197 156 2249
rect 0 2073 156 2125
rect 0 1949 156 2001
rect 0 1825 156 1877
rect 0 1701 156 1753
rect 0 1577 156 1629
rect 0 1453 156 1505
rect 0 1329 156 1381
rect 0 1205 156 1257
rect 0 1081 156 1133
rect 0 957 156 1009
rect 0 833 156 885
rect 0 709 156 761
rect 0 585 156 637
rect 0 461 156 513
rect 482 7893 534 7945
rect 606 7893 658 7945
rect 730 7893 782 7945
rect 854 7893 906 7945
rect 978 7893 1030 7945
rect 1102 7893 1154 7945
rect 1226 7893 1278 7945
rect 1350 7893 1402 7945
rect 1474 7893 1526 7945
rect 1598 7893 1650 7945
rect 1722 7893 1774 7945
rect 1846 7893 1898 7945
rect 1970 7893 2022 7945
rect 482 7769 534 7821
rect 606 7769 658 7821
rect 730 7769 782 7821
rect 854 7769 906 7821
rect 978 7769 1030 7821
rect 1102 7769 1154 7821
rect 1226 7769 1278 7821
rect 1350 7769 1402 7821
rect 1474 7769 1526 7821
rect 1598 7769 1650 7821
rect 1722 7769 1774 7821
rect 1846 7769 1898 7821
rect 1970 7769 2022 7821
rect 482 7645 534 7697
rect 606 7645 658 7697
rect 730 7645 782 7697
rect 854 7645 906 7697
rect 978 7645 1030 7697
rect 1102 7645 1154 7697
rect 1226 7645 1278 7697
rect 1350 7645 1402 7697
rect 1474 7645 1526 7697
rect 1598 7645 1650 7697
rect 1722 7645 1774 7697
rect 1846 7645 1898 7697
rect 1970 7645 2022 7697
rect 482 7521 534 7573
rect 606 7521 658 7573
rect 730 7521 782 7573
rect 854 7521 906 7573
rect 978 7521 1030 7573
rect 1102 7521 1154 7573
rect 1226 7521 1278 7573
rect 1350 7521 1402 7573
rect 1474 7521 1526 7573
rect 1598 7521 1650 7573
rect 1722 7521 1774 7573
rect 1846 7521 1898 7573
rect 1970 7521 2022 7573
rect 482 7397 534 7449
rect 606 7397 658 7449
rect 730 7397 782 7449
rect 854 7397 906 7449
rect 978 7397 1030 7449
rect 1102 7397 1154 7449
rect 1226 7397 1278 7449
rect 1350 7397 1402 7449
rect 1474 7397 1526 7449
rect 1598 7397 1650 7449
rect 1722 7397 1774 7449
rect 1846 7397 1898 7449
rect 1970 7397 2022 7449
rect 482 7273 534 7325
rect 606 7273 658 7325
rect 730 7273 782 7325
rect 854 7273 906 7325
rect 978 7273 1030 7325
rect 1102 7273 1154 7325
rect 1226 7273 1278 7325
rect 1350 7273 1402 7325
rect 1474 7273 1526 7325
rect 1598 7273 1650 7325
rect 1722 7273 1774 7325
rect 1846 7273 1898 7325
rect 1970 7273 2022 7325
rect 482 7149 534 7201
rect 606 7149 658 7201
rect 730 7149 782 7201
rect 854 7149 906 7201
rect 978 7149 1030 7201
rect 1102 7149 1154 7201
rect 1226 7149 1278 7201
rect 1350 7149 1402 7201
rect 1474 7149 1526 7201
rect 1598 7149 1650 7201
rect 1722 7149 1774 7201
rect 1846 7149 1898 7201
rect 1970 7149 2022 7201
rect 482 7025 534 7077
rect 606 7025 658 7077
rect 730 7025 782 7077
rect 854 7025 906 7077
rect 978 7025 1030 7077
rect 1102 7025 1154 7077
rect 1226 7025 1278 7077
rect 1350 7025 1402 7077
rect 1474 7025 1526 7077
rect 1598 7025 1650 7077
rect 1722 7025 1774 7077
rect 1846 7025 1898 7077
rect 1970 7025 2022 7077
rect 482 6901 534 6953
rect 606 6901 658 6953
rect 730 6901 782 6953
rect 854 6901 906 6953
rect 978 6901 1030 6953
rect 1102 6901 1154 6953
rect 1226 6901 1278 6953
rect 1350 6901 1402 6953
rect 1474 6901 1526 6953
rect 1598 6901 1650 6953
rect 1722 6901 1774 6953
rect 1846 6901 1898 6953
rect 1970 6901 2022 6953
rect 482 6777 534 6829
rect 606 6777 658 6829
rect 730 6777 782 6829
rect 854 6777 906 6829
rect 978 6777 1030 6829
rect 1102 6777 1154 6829
rect 1226 6777 1278 6829
rect 1350 6777 1402 6829
rect 1474 6777 1526 6829
rect 1598 6777 1650 6829
rect 1722 6777 1774 6829
rect 1846 6777 1898 6829
rect 1970 6777 2022 6829
rect 482 6653 534 6705
rect 606 6653 658 6705
rect 730 6653 782 6705
rect 854 6653 906 6705
rect 978 6653 1030 6705
rect 1102 6653 1154 6705
rect 1226 6653 1278 6705
rect 1350 6653 1402 6705
rect 1474 6653 1526 6705
rect 1598 6653 1650 6705
rect 1722 6653 1774 6705
rect 1846 6653 1898 6705
rect 1970 6653 2022 6705
rect 482 6529 534 6581
rect 606 6529 658 6581
rect 730 6529 782 6581
rect 854 6529 906 6581
rect 978 6529 1030 6581
rect 1102 6529 1154 6581
rect 1226 6529 1278 6581
rect 1350 6529 1402 6581
rect 1474 6529 1526 6581
rect 1598 6529 1650 6581
rect 1722 6529 1774 6581
rect 1846 6529 1898 6581
rect 1970 6529 2022 6581
rect 482 6405 534 6457
rect 606 6405 658 6457
rect 730 6405 782 6457
rect 854 6405 906 6457
rect 978 6405 1030 6457
rect 1102 6405 1154 6457
rect 1226 6405 1278 6457
rect 1350 6405 1402 6457
rect 1474 6405 1526 6457
rect 1598 6405 1650 6457
rect 1722 6405 1774 6457
rect 1846 6405 1898 6457
rect 1970 6405 2022 6457
rect 482 6281 534 6333
rect 606 6281 658 6333
rect 730 6281 782 6333
rect 854 6281 906 6333
rect 978 6281 1030 6333
rect 1102 6281 1154 6333
rect 1226 6281 1278 6333
rect 1350 6281 1402 6333
rect 1474 6281 1526 6333
rect 1598 6281 1650 6333
rect 1722 6281 1774 6333
rect 1846 6281 1898 6333
rect 1970 6281 2022 6333
rect 482 6157 534 6209
rect 606 6157 658 6209
rect 730 6157 782 6209
rect 854 6157 906 6209
rect 978 6157 1030 6209
rect 1102 6157 1154 6209
rect 1226 6157 1278 6209
rect 1350 6157 1402 6209
rect 1474 6157 1526 6209
rect 1598 6157 1650 6209
rect 1722 6157 1774 6209
rect 1846 6157 1898 6209
rect 1970 6157 2022 6209
rect 482 6033 534 6085
rect 606 6033 658 6085
rect 730 6033 782 6085
rect 854 6033 906 6085
rect 978 6033 1030 6085
rect 1102 6033 1154 6085
rect 1226 6033 1278 6085
rect 1350 6033 1402 6085
rect 1474 6033 1526 6085
rect 1598 6033 1650 6085
rect 1722 6033 1774 6085
rect 1846 6033 1898 6085
rect 1970 6033 2022 6085
rect 482 5909 534 5961
rect 606 5909 658 5961
rect 730 5909 782 5961
rect 854 5909 906 5961
rect 978 5909 1030 5961
rect 1102 5909 1154 5961
rect 1226 5909 1278 5961
rect 1350 5909 1402 5961
rect 1474 5909 1526 5961
rect 1598 5909 1650 5961
rect 1722 5909 1774 5961
rect 1846 5909 1898 5961
rect 1970 5909 2022 5961
rect 482 5785 534 5837
rect 606 5785 658 5837
rect 730 5785 782 5837
rect 854 5785 906 5837
rect 978 5785 1030 5837
rect 1102 5785 1154 5837
rect 1226 5785 1278 5837
rect 1350 5785 1402 5837
rect 1474 5785 1526 5837
rect 1598 5785 1650 5837
rect 1722 5785 1774 5837
rect 1846 5785 1898 5837
rect 1970 5785 2022 5837
rect 482 5661 534 5713
rect 606 5661 658 5713
rect 730 5661 782 5713
rect 854 5661 906 5713
rect 978 5661 1030 5713
rect 1102 5661 1154 5713
rect 1226 5661 1278 5713
rect 1350 5661 1402 5713
rect 1474 5661 1526 5713
rect 1598 5661 1650 5713
rect 1722 5661 1774 5713
rect 1846 5661 1898 5713
rect 1970 5661 2022 5713
rect 482 5537 534 5589
rect 606 5537 658 5589
rect 730 5537 782 5589
rect 854 5537 906 5589
rect 978 5537 1030 5589
rect 1102 5537 1154 5589
rect 1226 5537 1278 5589
rect 1350 5537 1402 5589
rect 1474 5537 1526 5589
rect 1598 5537 1650 5589
rect 1722 5537 1774 5589
rect 1846 5537 1898 5589
rect 1970 5537 2022 5589
rect 482 5413 534 5465
rect 606 5413 658 5465
rect 730 5413 782 5465
rect 854 5413 906 5465
rect 978 5413 1030 5465
rect 1102 5413 1154 5465
rect 1226 5413 1278 5465
rect 1350 5413 1402 5465
rect 1474 5413 1526 5465
rect 1598 5413 1650 5465
rect 1722 5413 1774 5465
rect 1846 5413 1898 5465
rect 1970 5413 2022 5465
rect 482 5289 534 5341
rect 606 5289 658 5341
rect 730 5289 782 5341
rect 854 5289 906 5341
rect 978 5289 1030 5341
rect 1102 5289 1154 5341
rect 1226 5289 1278 5341
rect 1350 5289 1402 5341
rect 1474 5289 1526 5341
rect 1598 5289 1650 5341
rect 1722 5289 1774 5341
rect 1846 5289 1898 5341
rect 1970 5289 2022 5341
rect 482 5165 534 5217
rect 606 5165 658 5217
rect 730 5165 782 5217
rect 854 5165 906 5217
rect 978 5165 1030 5217
rect 1102 5165 1154 5217
rect 1226 5165 1278 5217
rect 1350 5165 1402 5217
rect 1474 5165 1526 5217
rect 1598 5165 1650 5217
rect 1722 5165 1774 5217
rect 1846 5165 1898 5217
rect 1970 5165 2022 5217
rect 482 5041 534 5093
rect 606 5041 658 5093
rect 730 5041 782 5093
rect 854 5041 906 5093
rect 978 5041 1030 5093
rect 1102 5041 1154 5093
rect 1226 5041 1278 5093
rect 1350 5041 1402 5093
rect 1474 5041 1526 5093
rect 1598 5041 1650 5093
rect 1722 5041 1774 5093
rect 1846 5041 1898 5093
rect 1970 5041 2022 5093
rect 482 4917 534 4969
rect 606 4917 658 4969
rect 730 4917 782 4969
rect 854 4917 906 4969
rect 978 4917 1030 4969
rect 1102 4917 1154 4969
rect 1226 4917 1278 4969
rect 1350 4917 1402 4969
rect 1474 4917 1526 4969
rect 1598 4917 1650 4969
rect 1722 4917 1774 4969
rect 1846 4917 1898 4969
rect 1970 4917 2022 4969
rect 482 4793 534 4845
rect 606 4793 658 4845
rect 730 4793 782 4845
rect 854 4793 906 4845
rect 978 4793 1030 4845
rect 1102 4793 1154 4845
rect 1226 4793 1278 4845
rect 1350 4793 1402 4845
rect 1474 4793 1526 4845
rect 1598 4793 1650 4845
rect 1722 4793 1774 4845
rect 1846 4793 1898 4845
rect 1970 4793 2022 4845
rect 482 4669 534 4721
rect 606 4669 658 4721
rect 730 4669 782 4721
rect 854 4669 906 4721
rect 978 4669 1030 4721
rect 1102 4669 1154 4721
rect 1226 4669 1278 4721
rect 1350 4669 1402 4721
rect 1474 4669 1526 4721
rect 1598 4669 1650 4721
rect 1722 4669 1774 4721
rect 1846 4669 1898 4721
rect 1970 4669 2022 4721
rect 482 4545 534 4597
rect 606 4545 658 4597
rect 730 4545 782 4597
rect 854 4545 906 4597
rect 978 4545 1030 4597
rect 1102 4545 1154 4597
rect 1226 4545 1278 4597
rect 1350 4545 1402 4597
rect 1474 4545 1526 4597
rect 1598 4545 1650 4597
rect 1722 4545 1774 4597
rect 1846 4545 1898 4597
rect 1970 4545 2022 4597
rect 482 4421 534 4473
rect 606 4421 658 4473
rect 730 4421 782 4473
rect 854 4421 906 4473
rect 978 4421 1030 4473
rect 1102 4421 1154 4473
rect 1226 4421 1278 4473
rect 1350 4421 1402 4473
rect 1474 4421 1526 4473
rect 1598 4421 1650 4473
rect 1722 4421 1774 4473
rect 1846 4421 1898 4473
rect 1970 4421 2022 4473
rect 482 4297 534 4349
rect 606 4297 658 4349
rect 730 4297 782 4349
rect 854 4297 906 4349
rect 978 4297 1030 4349
rect 1102 4297 1154 4349
rect 1226 4297 1278 4349
rect 1350 4297 1402 4349
rect 1474 4297 1526 4349
rect 1598 4297 1650 4349
rect 1722 4297 1774 4349
rect 1846 4297 1898 4349
rect 1970 4297 2022 4349
rect 482 4173 534 4225
rect 606 4173 658 4225
rect 730 4173 782 4225
rect 854 4173 906 4225
rect 978 4173 1030 4225
rect 1102 4173 1154 4225
rect 1226 4173 1278 4225
rect 1350 4173 1402 4225
rect 1474 4173 1526 4225
rect 1598 4173 1650 4225
rect 1722 4173 1774 4225
rect 1846 4173 1898 4225
rect 1970 4173 2022 4225
rect 482 4049 534 4101
rect 606 4049 658 4101
rect 730 4049 782 4101
rect 854 4049 906 4101
rect 978 4049 1030 4101
rect 1102 4049 1154 4101
rect 1226 4049 1278 4101
rect 1350 4049 1402 4101
rect 1474 4049 1526 4101
rect 1598 4049 1650 4101
rect 1722 4049 1774 4101
rect 1846 4049 1898 4101
rect 1970 4049 2022 4101
rect 482 3925 534 3977
rect 606 3925 658 3977
rect 730 3925 782 3977
rect 854 3925 906 3977
rect 978 3925 1030 3977
rect 1102 3925 1154 3977
rect 1226 3925 1278 3977
rect 1350 3925 1402 3977
rect 1474 3925 1526 3977
rect 1598 3925 1650 3977
rect 1722 3925 1774 3977
rect 1846 3925 1898 3977
rect 1970 3925 2022 3977
rect 482 3801 534 3853
rect 606 3801 658 3853
rect 730 3801 782 3853
rect 854 3801 906 3853
rect 978 3801 1030 3853
rect 1102 3801 1154 3853
rect 1226 3801 1278 3853
rect 1350 3801 1402 3853
rect 1474 3801 1526 3853
rect 1598 3801 1650 3853
rect 1722 3801 1774 3853
rect 1846 3801 1898 3853
rect 1970 3801 2022 3853
rect 482 3677 534 3729
rect 606 3677 658 3729
rect 730 3677 782 3729
rect 854 3677 906 3729
rect 978 3677 1030 3729
rect 1102 3677 1154 3729
rect 1226 3677 1278 3729
rect 1350 3677 1402 3729
rect 1474 3677 1526 3729
rect 1598 3677 1650 3729
rect 1722 3677 1774 3729
rect 1846 3677 1898 3729
rect 1970 3677 2022 3729
rect 482 3553 534 3605
rect 606 3553 658 3605
rect 730 3553 782 3605
rect 854 3553 906 3605
rect 978 3553 1030 3605
rect 1102 3553 1154 3605
rect 1226 3553 1278 3605
rect 1350 3553 1402 3605
rect 1474 3553 1526 3605
rect 1598 3553 1650 3605
rect 1722 3553 1774 3605
rect 1846 3553 1898 3605
rect 1970 3553 2022 3605
rect 482 3429 534 3481
rect 606 3429 658 3481
rect 730 3429 782 3481
rect 854 3429 906 3481
rect 978 3429 1030 3481
rect 1102 3429 1154 3481
rect 1226 3429 1278 3481
rect 1350 3429 1402 3481
rect 1474 3429 1526 3481
rect 1598 3429 1650 3481
rect 1722 3429 1774 3481
rect 1846 3429 1898 3481
rect 1970 3429 2022 3481
rect 482 3305 534 3357
rect 606 3305 658 3357
rect 730 3305 782 3357
rect 854 3305 906 3357
rect 978 3305 1030 3357
rect 1102 3305 1154 3357
rect 1226 3305 1278 3357
rect 1350 3305 1402 3357
rect 1474 3305 1526 3357
rect 1598 3305 1650 3357
rect 1722 3305 1774 3357
rect 1846 3305 1898 3357
rect 1970 3305 2022 3357
rect 482 3181 534 3233
rect 606 3181 658 3233
rect 730 3181 782 3233
rect 854 3181 906 3233
rect 978 3181 1030 3233
rect 1102 3181 1154 3233
rect 1226 3181 1278 3233
rect 1350 3181 1402 3233
rect 1474 3181 1526 3233
rect 1598 3181 1650 3233
rect 1722 3181 1774 3233
rect 1846 3181 1898 3233
rect 1970 3181 2022 3233
rect 482 3057 534 3109
rect 606 3057 658 3109
rect 730 3057 782 3109
rect 854 3057 906 3109
rect 978 3057 1030 3109
rect 1102 3057 1154 3109
rect 1226 3057 1278 3109
rect 1350 3057 1402 3109
rect 1474 3057 1526 3109
rect 1598 3057 1650 3109
rect 1722 3057 1774 3109
rect 1846 3057 1898 3109
rect 1970 3057 2022 3109
rect 482 2933 534 2985
rect 606 2933 658 2985
rect 730 2933 782 2985
rect 854 2933 906 2985
rect 978 2933 1030 2985
rect 1102 2933 1154 2985
rect 1226 2933 1278 2985
rect 1350 2933 1402 2985
rect 1474 2933 1526 2985
rect 1598 2933 1650 2985
rect 1722 2933 1774 2985
rect 1846 2933 1898 2985
rect 1970 2933 2022 2985
rect 482 2809 534 2861
rect 606 2809 658 2861
rect 730 2809 782 2861
rect 854 2809 906 2861
rect 978 2809 1030 2861
rect 1102 2809 1154 2861
rect 1226 2809 1278 2861
rect 1350 2809 1402 2861
rect 1474 2809 1526 2861
rect 1598 2809 1650 2861
rect 1722 2809 1774 2861
rect 1846 2809 1898 2861
rect 1970 2809 2022 2861
rect 482 2685 534 2737
rect 606 2685 658 2737
rect 730 2685 782 2737
rect 854 2685 906 2737
rect 978 2685 1030 2737
rect 1102 2685 1154 2737
rect 1226 2685 1278 2737
rect 1350 2685 1402 2737
rect 1474 2685 1526 2737
rect 1598 2685 1650 2737
rect 1722 2685 1774 2737
rect 1846 2685 1898 2737
rect 1970 2685 2022 2737
rect 482 2561 534 2613
rect 606 2561 658 2613
rect 730 2561 782 2613
rect 854 2561 906 2613
rect 978 2561 1030 2613
rect 1102 2561 1154 2613
rect 1226 2561 1278 2613
rect 1350 2561 1402 2613
rect 1474 2561 1526 2613
rect 1598 2561 1650 2613
rect 1722 2561 1774 2613
rect 1846 2561 1898 2613
rect 1970 2561 2022 2613
rect 482 2437 534 2489
rect 606 2437 658 2489
rect 730 2437 782 2489
rect 854 2437 906 2489
rect 978 2437 1030 2489
rect 1102 2437 1154 2489
rect 1226 2437 1278 2489
rect 1350 2437 1402 2489
rect 1474 2437 1526 2489
rect 1598 2437 1650 2489
rect 1722 2437 1774 2489
rect 1846 2437 1898 2489
rect 1970 2437 2022 2489
rect 482 2313 534 2365
rect 606 2313 658 2365
rect 730 2313 782 2365
rect 854 2313 906 2365
rect 978 2313 1030 2365
rect 1102 2313 1154 2365
rect 1226 2313 1278 2365
rect 1350 2313 1402 2365
rect 1474 2313 1526 2365
rect 1598 2313 1650 2365
rect 1722 2313 1774 2365
rect 1846 2313 1898 2365
rect 1970 2313 2022 2365
rect 482 2189 534 2241
rect 606 2189 658 2241
rect 730 2189 782 2241
rect 854 2189 906 2241
rect 978 2189 1030 2241
rect 1102 2189 1154 2241
rect 1226 2189 1278 2241
rect 1350 2189 1402 2241
rect 1474 2189 1526 2241
rect 1598 2189 1650 2241
rect 1722 2189 1774 2241
rect 1846 2189 1898 2241
rect 1970 2189 2022 2241
rect 482 2065 534 2117
rect 606 2065 658 2117
rect 730 2065 782 2117
rect 854 2065 906 2117
rect 978 2065 1030 2117
rect 1102 2065 1154 2117
rect 1226 2065 1278 2117
rect 1350 2065 1402 2117
rect 1474 2065 1526 2117
rect 1598 2065 1650 2117
rect 1722 2065 1774 2117
rect 1846 2065 1898 2117
rect 1970 2065 2022 2117
rect 482 1941 534 1993
rect 606 1941 658 1993
rect 730 1941 782 1993
rect 854 1941 906 1993
rect 978 1941 1030 1993
rect 1102 1941 1154 1993
rect 1226 1941 1278 1993
rect 1350 1941 1402 1993
rect 1474 1941 1526 1993
rect 1598 1941 1650 1993
rect 1722 1941 1774 1993
rect 1846 1941 1898 1993
rect 1970 1941 2022 1993
rect 482 1817 534 1869
rect 606 1817 658 1869
rect 730 1817 782 1869
rect 854 1817 906 1869
rect 978 1817 1030 1869
rect 1102 1817 1154 1869
rect 1226 1817 1278 1869
rect 1350 1817 1402 1869
rect 1474 1817 1526 1869
rect 1598 1817 1650 1869
rect 1722 1817 1774 1869
rect 1846 1817 1898 1869
rect 1970 1817 2022 1869
rect 482 1693 534 1745
rect 606 1693 658 1745
rect 730 1693 782 1745
rect 854 1693 906 1745
rect 978 1693 1030 1745
rect 1102 1693 1154 1745
rect 1226 1693 1278 1745
rect 1350 1693 1402 1745
rect 1474 1693 1526 1745
rect 1598 1693 1650 1745
rect 1722 1693 1774 1745
rect 1846 1693 1898 1745
rect 1970 1693 2022 1745
rect 482 1569 534 1621
rect 606 1569 658 1621
rect 730 1569 782 1621
rect 854 1569 906 1621
rect 978 1569 1030 1621
rect 1102 1569 1154 1621
rect 1226 1569 1278 1621
rect 1350 1569 1402 1621
rect 1474 1569 1526 1621
rect 1598 1569 1650 1621
rect 1722 1569 1774 1621
rect 1846 1569 1898 1621
rect 1970 1569 2022 1621
rect 482 1445 534 1497
rect 606 1445 658 1497
rect 730 1445 782 1497
rect 854 1445 906 1497
rect 978 1445 1030 1497
rect 1102 1445 1154 1497
rect 1226 1445 1278 1497
rect 1350 1445 1402 1497
rect 1474 1445 1526 1497
rect 1598 1445 1650 1497
rect 1722 1445 1774 1497
rect 1846 1445 1898 1497
rect 1970 1445 2022 1497
rect 482 1321 534 1373
rect 606 1321 658 1373
rect 730 1321 782 1373
rect 854 1321 906 1373
rect 978 1321 1030 1373
rect 1102 1321 1154 1373
rect 1226 1321 1278 1373
rect 1350 1321 1402 1373
rect 1474 1321 1526 1373
rect 1598 1321 1650 1373
rect 1722 1321 1774 1373
rect 1846 1321 1898 1373
rect 1970 1321 2022 1373
rect 482 1197 534 1249
rect 606 1197 658 1249
rect 730 1197 782 1249
rect 854 1197 906 1249
rect 978 1197 1030 1249
rect 1102 1197 1154 1249
rect 1226 1197 1278 1249
rect 1350 1197 1402 1249
rect 1474 1197 1526 1249
rect 1598 1197 1650 1249
rect 1722 1197 1774 1249
rect 1846 1197 1898 1249
rect 1970 1197 2022 1249
rect 482 1073 534 1125
rect 606 1073 658 1125
rect 730 1073 782 1125
rect 854 1073 906 1125
rect 978 1073 1030 1125
rect 1102 1073 1154 1125
rect 1226 1073 1278 1125
rect 1350 1073 1402 1125
rect 1474 1073 1526 1125
rect 1598 1073 1650 1125
rect 1722 1073 1774 1125
rect 1846 1073 1898 1125
rect 1970 1073 2022 1125
rect 482 949 534 1001
rect 606 949 658 1001
rect 730 949 782 1001
rect 854 949 906 1001
rect 978 949 1030 1001
rect 1102 949 1154 1001
rect 1226 949 1278 1001
rect 1350 949 1402 1001
rect 1474 949 1526 1001
rect 1598 949 1650 1001
rect 1722 949 1774 1001
rect 1846 949 1898 1001
rect 1970 949 2022 1001
rect 482 825 534 877
rect 606 825 658 877
rect 730 825 782 877
rect 854 825 906 877
rect 978 825 1030 877
rect 1102 825 1154 877
rect 1226 825 1278 877
rect 1350 825 1402 877
rect 1474 825 1526 877
rect 1598 825 1650 877
rect 1722 825 1774 877
rect 1846 825 1898 877
rect 1970 825 2022 877
rect 482 701 534 753
rect 606 701 658 753
rect 730 701 782 753
rect 854 701 906 753
rect 978 701 1030 753
rect 1102 701 1154 753
rect 1226 701 1278 753
rect 1350 701 1402 753
rect 1474 701 1526 753
rect 1598 701 1650 753
rect 1722 701 1774 753
rect 1846 701 1898 753
rect 1970 701 2022 753
rect 482 577 534 629
rect 606 577 658 629
rect 730 577 782 629
rect 854 577 906 629
rect 978 577 1030 629
rect 1102 577 1154 629
rect 1226 577 1278 629
rect 1350 577 1402 629
rect 1474 577 1526 629
rect 1598 577 1650 629
rect 1722 577 1774 629
rect 1846 577 1898 629
rect 1970 577 2022 629
rect 482 453 534 505
rect 606 453 658 505
rect 730 453 782 505
rect 854 453 906 505
rect 978 453 1030 505
rect 1102 453 1154 505
rect 1226 453 1278 505
rect 1350 453 1402 505
rect 1474 453 1526 505
rect 1598 453 1650 505
rect 1722 453 1774 505
rect 1846 453 1898 505
rect 1970 453 2022 505
<< metal2 >>
rect -44 7953 200 8000
rect -44 7901 0 7953
rect 156 7901 200 7953
rect -44 7829 200 7901
rect -44 7777 0 7829
rect 156 7777 200 7829
rect -44 7705 200 7777
rect -44 7653 0 7705
rect 156 7653 200 7705
rect -44 7648 200 7653
rect -44 6032 0 7648
rect 160 6032 200 7648
rect -44 5969 200 6032
rect -44 5917 0 5969
rect 156 5917 200 5969
rect -44 5845 200 5917
rect -44 5793 0 5845
rect 156 5793 200 5845
rect -44 5721 200 5793
rect -44 5669 0 5721
rect 156 5669 200 5721
rect -44 5597 200 5669
rect -44 5545 0 5597
rect 156 5545 200 5597
rect -44 5473 200 5545
rect -44 5421 0 5473
rect 156 5421 200 5473
rect -44 5349 200 5421
rect -44 5297 0 5349
rect 156 5297 200 5349
rect -44 5225 200 5297
rect -44 5173 0 5225
rect 156 5173 200 5225
rect -44 5101 200 5173
rect -44 5049 0 5101
rect 156 5049 200 5101
rect -44 5047 200 5049
rect -44 2911 0 5047
rect 160 2911 200 5047
rect -44 2869 200 2911
rect -44 2817 0 2869
rect 156 2817 200 2869
rect -44 2745 200 2817
rect -44 2693 0 2745
rect 156 2693 200 2745
rect -44 2621 200 2693
rect -44 2569 0 2621
rect 156 2569 200 2621
rect -44 2497 200 2569
rect -44 2445 0 2497
rect 156 2445 200 2497
rect -44 2373 200 2445
rect -44 2321 0 2373
rect 156 2321 200 2373
rect -44 2249 200 2321
rect -44 2197 0 2249
rect 156 2197 200 2249
rect -44 2125 200 2197
rect -44 2073 0 2125
rect 156 2073 200 2125
rect -44 2001 200 2073
rect -44 688 0 2001
rect 156 1992 200 2001
rect 160 688 200 1992
rect -44 637 200 688
rect -44 585 0 637
rect 156 585 200 637
rect -44 513 200 585
rect -44 461 0 513
rect 156 461 200 513
rect -44 400 200 461
rect 430 7945 2074 8000
rect 430 7893 482 7945
rect 534 7893 606 7945
rect 658 7893 730 7945
rect 782 7893 854 7945
rect 906 7893 978 7945
rect 1030 7893 1102 7945
rect 1154 7893 1226 7945
rect 1278 7893 1350 7945
rect 1402 7893 1474 7945
rect 1526 7893 1598 7945
rect 1650 7893 1722 7945
rect 1774 7893 1846 7945
rect 1898 7893 1970 7945
rect 2022 7893 2074 7945
rect 430 7821 2074 7893
rect 430 7769 482 7821
rect 534 7769 606 7821
rect 658 7769 730 7821
rect 782 7769 854 7821
rect 906 7769 978 7821
rect 1030 7769 1102 7821
rect 1154 7769 1226 7821
rect 1278 7769 1350 7821
rect 1402 7769 1474 7821
rect 1526 7769 1598 7821
rect 1650 7769 1722 7821
rect 1774 7769 1846 7821
rect 1898 7769 1970 7821
rect 2022 7769 2074 7821
rect 430 7697 2074 7769
rect 430 7645 482 7697
rect 534 7645 606 7697
rect 658 7645 730 7697
rect 782 7645 854 7697
rect 906 7645 978 7697
rect 1030 7645 1102 7697
rect 1154 7645 1226 7697
rect 1278 7645 1350 7697
rect 1402 7645 1474 7697
rect 1526 7645 1598 7697
rect 1650 7645 1722 7697
rect 1774 7645 1846 7697
rect 1898 7645 1970 7697
rect 2022 7645 2074 7697
rect 430 7573 2074 7645
rect 430 7521 482 7573
rect 534 7521 606 7573
rect 658 7521 730 7573
rect 782 7521 854 7573
rect 906 7521 978 7573
rect 1030 7521 1102 7573
rect 1154 7521 1226 7573
rect 1278 7521 1350 7573
rect 1402 7521 1474 7573
rect 1526 7521 1598 7573
rect 1650 7521 1722 7573
rect 1774 7521 1846 7573
rect 1898 7521 1970 7573
rect 2022 7521 2074 7573
rect 430 7449 2074 7521
rect 430 7397 482 7449
rect 534 7397 606 7449
rect 658 7397 730 7449
rect 782 7397 854 7449
rect 906 7397 978 7449
rect 1030 7397 1102 7449
rect 1154 7397 1226 7449
rect 1278 7397 1350 7449
rect 1402 7397 1474 7449
rect 1526 7397 1598 7449
rect 1650 7397 1722 7449
rect 1774 7397 1846 7449
rect 1898 7397 1970 7449
rect 2022 7397 2074 7449
rect 430 7325 2074 7397
rect 430 7273 482 7325
rect 534 7273 606 7325
rect 658 7273 730 7325
rect 782 7273 854 7325
rect 906 7273 978 7325
rect 1030 7273 1102 7325
rect 1154 7273 1226 7325
rect 1278 7273 1350 7325
rect 1402 7273 1474 7325
rect 1526 7273 1598 7325
rect 1650 7273 1722 7325
rect 1774 7273 1846 7325
rect 1898 7273 1970 7325
rect 2022 7273 2074 7325
rect 430 7201 2074 7273
rect 430 7149 482 7201
rect 534 7149 606 7201
rect 658 7149 730 7201
rect 782 7149 854 7201
rect 906 7149 978 7201
rect 1030 7149 1102 7201
rect 1154 7149 1226 7201
rect 1278 7149 1350 7201
rect 1402 7149 1474 7201
rect 1526 7149 1598 7201
rect 1650 7149 1722 7201
rect 1774 7149 1846 7201
rect 1898 7149 1970 7201
rect 2022 7149 2074 7201
rect 430 7077 2074 7149
rect 430 7025 482 7077
rect 534 7025 606 7077
rect 658 7025 730 7077
rect 782 7025 854 7077
rect 906 7025 978 7077
rect 1030 7025 1102 7077
rect 1154 7025 1226 7077
rect 1278 7025 1350 7077
rect 1402 7025 1474 7077
rect 1526 7025 1598 7077
rect 1650 7025 1722 7077
rect 1774 7025 1846 7077
rect 1898 7025 1970 7077
rect 2022 7025 2074 7077
rect 430 6953 2074 7025
rect 430 6901 482 6953
rect 534 6901 606 6953
rect 658 6901 730 6953
rect 782 6901 854 6953
rect 906 6901 978 6953
rect 1030 6901 1102 6953
rect 1154 6901 1226 6953
rect 1278 6901 1350 6953
rect 1402 6901 1474 6953
rect 1526 6901 1598 6953
rect 1650 6901 1722 6953
rect 1774 6901 1846 6953
rect 1898 6901 1970 6953
rect 2022 6901 2074 6953
rect 430 6829 2074 6901
rect 430 6777 482 6829
rect 534 6777 606 6829
rect 658 6777 730 6829
rect 782 6777 854 6829
rect 906 6777 978 6829
rect 1030 6777 1102 6829
rect 1154 6777 1226 6829
rect 1278 6777 1350 6829
rect 1402 6777 1474 6829
rect 1526 6777 1598 6829
rect 1650 6777 1722 6829
rect 1774 6777 1846 6829
rect 1898 6777 1970 6829
rect 2022 6777 2074 6829
rect 430 6705 2074 6777
rect 430 6653 482 6705
rect 534 6653 606 6705
rect 658 6653 730 6705
rect 782 6653 854 6705
rect 906 6653 978 6705
rect 1030 6653 1102 6705
rect 1154 6653 1226 6705
rect 1278 6653 1350 6705
rect 1402 6653 1474 6705
rect 1526 6653 1598 6705
rect 1650 6653 1722 6705
rect 1774 6653 1846 6705
rect 1898 6653 1970 6705
rect 2022 6653 2074 6705
rect 430 6581 2074 6653
rect 430 6529 482 6581
rect 534 6529 606 6581
rect 658 6529 730 6581
rect 782 6529 854 6581
rect 906 6529 978 6581
rect 1030 6529 1102 6581
rect 1154 6529 1226 6581
rect 1278 6529 1350 6581
rect 1402 6529 1474 6581
rect 1526 6529 1598 6581
rect 1650 6529 1722 6581
rect 1774 6529 1846 6581
rect 1898 6529 1970 6581
rect 2022 6529 2074 6581
rect 430 6457 2074 6529
rect 430 6405 482 6457
rect 534 6405 606 6457
rect 658 6405 730 6457
rect 782 6405 854 6457
rect 906 6405 978 6457
rect 1030 6405 1102 6457
rect 1154 6405 1226 6457
rect 1278 6405 1350 6457
rect 1402 6405 1474 6457
rect 1526 6405 1598 6457
rect 1650 6405 1722 6457
rect 1774 6405 1846 6457
rect 1898 6405 1970 6457
rect 2022 6405 2074 6457
rect 430 6333 2074 6405
rect 430 6281 482 6333
rect 534 6281 606 6333
rect 658 6281 730 6333
rect 782 6281 854 6333
rect 906 6281 978 6333
rect 1030 6281 1102 6333
rect 1154 6281 1226 6333
rect 1278 6281 1350 6333
rect 1402 6281 1474 6333
rect 1526 6281 1598 6333
rect 1650 6281 1722 6333
rect 1774 6281 1846 6333
rect 1898 6281 1970 6333
rect 2022 6281 2074 6333
rect 430 6209 2074 6281
rect 430 6157 482 6209
rect 534 6157 606 6209
rect 658 6157 730 6209
rect 782 6157 854 6209
rect 906 6157 978 6209
rect 1030 6157 1102 6209
rect 1154 6157 1226 6209
rect 1278 6157 1350 6209
rect 1402 6157 1474 6209
rect 1526 6157 1598 6209
rect 1650 6157 1722 6209
rect 1774 6157 1846 6209
rect 1898 6157 1970 6209
rect 2022 6157 2074 6209
rect 430 6085 2074 6157
rect 430 6033 482 6085
rect 534 6033 606 6085
rect 658 6033 730 6085
rect 782 6033 854 6085
rect 906 6033 978 6085
rect 1030 6033 1102 6085
rect 1154 6033 1226 6085
rect 1278 6033 1350 6085
rect 1402 6033 1474 6085
rect 1526 6033 1598 6085
rect 1650 6033 1722 6085
rect 1774 6033 1846 6085
rect 1898 6033 1970 6085
rect 2022 6033 2074 6085
rect 430 5961 2074 6033
rect 430 5909 482 5961
rect 534 5909 606 5961
rect 658 5909 730 5961
rect 782 5909 854 5961
rect 906 5909 978 5961
rect 1030 5909 1102 5961
rect 1154 5909 1226 5961
rect 1278 5909 1350 5961
rect 1402 5909 1474 5961
rect 1526 5909 1598 5961
rect 1650 5909 1722 5961
rect 1774 5909 1846 5961
rect 1898 5909 1970 5961
rect 2022 5909 2074 5961
rect 430 5837 2074 5909
rect 430 5785 482 5837
rect 534 5785 606 5837
rect 658 5785 730 5837
rect 782 5785 854 5837
rect 906 5785 978 5837
rect 1030 5785 1102 5837
rect 1154 5785 1226 5837
rect 1278 5785 1350 5837
rect 1402 5785 1474 5837
rect 1526 5785 1598 5837
rect 1650 5785 1722 5837
rect 1774 5785 1846 5837
rect 1898 5785 1970 5837
rect 2022 5785 2074 5837
rect 430 5713 2074 5785
rect 430 5661 482 5713
rect 534 5661 606 5713
rect 658 5661 730 5713
rect 782 5661 854 5713
rect 906 5661 978 5713
rect 1030 5661 1102 5713
rect 1154 5661 1226 5713
rect 1278 5661 1350 5713
rect 1402 5661 1474 5713
rect 1526 5661 1598 5713
rect 1650 5661 1722 5713
rect 1774 5661 1846 5713
rect 1898 5661 1970 5713
rect 2022 5661 2074 5713
rect 430 5589 2074 5661
rect 430 5537 482 5589
rect 534 5537 606 5589
rect 658 5537 730 5589
rect 782 5537 854 5589
rect 906 5537 978 5589
rect 1030 5537 1102 5589
rect 1154 5537 1226 5589
rect 1278 5537 1350 5589
rect 1402 5537 1474 5589
rect 1526 5537 1598 5589
rect 1650 5537 1722 5589
rect 1774 5537 1846 5589
rect 1898 5537 1970 5589
rect 2022 5537 2074 5589
rect 430 5465 2074 5537
rect 430 5413 482 5465
rect 534 5413 606 5465
rect 658 5413 730 5465
rect 782 5413 854 5465
rect 906 5413 978 5465
rect 1030 5413 1102 5465
rect 1154 5413 1226 5465
rect 1278 5413 1350 5465
rect 1402 5413 1474 5465
rect 1526 5413 1598 5465
rect 1650 5413 1722 5465
rect 1774 5413 1846 5465
rect 1898 5413 1970 5465
rect 2022 5413 2074 5465
rect 430 5341 2074 5413
rect 430 5289 482 5341
rect 534 5289 606 5341
rect 658 5289 730 5341
rect 782 5289 854 5341
rect 906 5289 978 5341
rect 1030 5289 1102 5341
rect 1154 5289 1226 5341
rect 1278 5289 1350 5341
rect 1402 5289 1474 5341
rect 1526 5289 1598 5341
rect 1650 5289 1722 5341
rect 1774 5289 1846 5341
rect 1898 5289 1970 5341
rect 2022 5289 2074 5341
rect 430 5217 2074 5289
rect 430 5165 482 5217
rect 534 5165 606 5217
rect 658 5165 730 5217
rect 782 5165 854 5217
rect 906 5165 978 5217
rect 1030 5165 1102 5217
rect 1154 5165 1226 5217
rect 1278 5165 1350 5217
rect 1402 5165 1474 5217
rect 1526 5165 1598 5217
rect 1650 5165 1722 5217
rect 1774 5165 1846 5217
rect 1898 5165 1970 5217
rect 2022 5165 2074 5217
rect 430 5093 2074 5165
rect 430 5041 482 5093
rect 534 5041 606 5093
rect 658 5041 730 5093
rect 782 5041 854 5093
rect 906 5041 978 5093
rect 1030 5041 1102 5093
rect 1154 5041 1226 5093
rect 1278 5041 1350 5093
rect 1402 5041 1474 5093
rect 1526 5041 1598 5093
rect 1650 5041 1722 5093
rect 1774 5041 1846 5093
rect 1898 5041 1970 5093
rect 2022 5041 2074 5093
rect 430 4969 2074 5041
rect 430 4917 482 4969
rect 534 4917 606 4969
rect 658 4917 730 4969
rect 782 4917 854 4969
rect 906 4917 978 4969
rect 1030 4917 1102 4969
rect 1154 4917 1226 4969
rect 1278 4917 1350 4969
rect 1402 4917 1474 4969
rect 1526 4917 1598 4969
rect 1650 4917 1722 4969
rect 1774 4917 1846 4969
rect 1898 4917 1970 4969
rect 2022 4917 2074 4969
rect 430 4845 2074 4917
rect 430 4793 482 4845
rect 534 4793 606 4845
rect 658 4793 730 4845
rect 782 4793 854 4845
rect 906 4793 978 4845
rect 1030 4793 1102 4845
rect 1154 4793 1226 4845
rect 1278 4793 1350 4845
rect 1402 4793 1474 4845
rect 1526 4793 1598 4845
rect 1650 4793 1722 4845
rect 1774 4793 1846 4845
rect 1898 4793 1970 4845
rect 2022 4793 2074 4845
rect 430 4721 2074 4793
rect 430 4669 482 4721
rect 534 4669 606 4721
rect 658 4669 730 4721
rect 782 4669 854 4721
rect 906 4669 978 4721
rect 1030 4669 1102 4721
rect 1154 4669 1226 4721
rect 1278 4669 1350 4721
rect 1402 4669 1474 4721
rect 1526 4669 1598 4721
rect 1650 4669 1722 4721
rect 1774 4669 1846 4721
rect 1898 4669 1970 4721
rect 2022 4669 2074 4721
rect 430 4597 2074 4669
rect 430 4545 482 4597
rect 534 4545 606 4597
rect 658 4545 730 4597
rect 782 4545 854 4597
rect 906 4545 978 4597
rect 1030 4545 1102 4597
rect 1154 4545 1226 4597
rect 1278 4545 1350 4597
rect 1402 4545 1474 4597
rect 1526 4545 1598 4597
rect 1650 4545 1722 4597
rect 1774 4545 1846 4597
rect 1898 4545 1970 4597
rect 2022 4545 2074 4597
rect 430 4473 2074 4545
rect 430 4421 482 4473
rect 534 4421 606 4473
rect 658 4421 730 4473
rect 782 4421 854 4473
rect 906 4421 978 4473
rect 1030 4421 1102 4473
rect 1154 4421 1226 4473
rect 1278 4421 1350 4473
rect 1402 4421 1474 4473
rect 1526 4421 1598 4473
rect 1650 4421 1722 4473
rect 1774 4421 1846 4473
rect 1898 4421 1970 4473
rect 2022 4421 2074 4473
rect 430 4349 2074 4421
rect 430 4297 482 4349
rect 534 4297 606 4349
rect 658 4297 730 4349
rect 782 4297 854 4349
rect 906 4297 978 4349
rect 1030 4297 1102 4349
rect 1154 4297 1226 4349
rect 1278 4297 1350 4349
rect 1402 4297 1474 4349
rect 1526 4297 1598 4349
rect 1650 4297 1722 4349
rect 1774 4297 1846 4349
rect 1898 4297 1970 4349
rect 2022 4297 2074 4349
rect 430 4225 2074 4297
rect 430 4173 482 4225
rect 534 4173 606 4225
rect 658 4173 730 4225
rect 782 4173 854 4225
rect 906 4173 978 4225
rect 1030 4173 1102 4225
rect 1154 4173 1226 4225
rect 1278 4173 1350 4225
rect 1402 4173 1474 4225
rect 1526 4173 1598 4225
rect 1650 4173 1722 4225
rect 1774 4173 1846 4225
rect 1898 4173 1970 4225
rect 2022 4173 2074 4225
rect 430 4101 2074 4173
rect 430 4049 482 4101
rect 534 4049 606 4101
rect 658 4049 730 4101
rect 782 4049 854 4101
rect 906 4049 978 4101
rect 1030 4049 1102 4101
rect 1154 4049 1226 4101
rect 1278 4049 1350 4101
rect 1402 4049 1474 4101
rect 1526 4049 1598 4101
rect 1650 4049 1722 4101
rect 1774 4049 1846 4101
rect 1898 4049 1970 4101
rect 2022 4049 2074 4101
rect 430 3977 2074 4049
rect 430 3925 482 3977
rect 534 3925 606 3977
rect 658 3925 730 3977
rect 782 3925 854 3977
rect 906 3925 978 3977
rect 1030 3925 1102 3977
rect 1154 3925 1226 3977
rect 1278 3925 1350 3977
rect 1402 3925 1474 3977
rect 1526 3925 1598 3977
rect 1650 3925 1722 3977
rect 1774 3925 1846 3977
rect 1898 3925 1970 3977
rect 2022 3925 2074 3977
rect 430 3853 2074 3925
rect 430 3801 482 3853
rect 534 3801 606 3853
rect 658 3801 730 3853
rect 782 3801 854 3853
rect 906 3801 978 3853
rect 1030 3801 1102 3853
rect 1154 3801 1226 3853
rect 1278 3801 1350 3853
rect 1402 3801 1474 3853
rect 1526 3801 1598 3853
rect 1650 3801 1722 3853
rect 1774 3801 1846 3853
rect 1898 3801 1970 3853
rect 2022 3801 2074 3853
rect 430 3729 2074 3801
rect 430 3677 482 3729
rect 534 3677 606 3729
rect 658 3677 730 3729
rect 782 3677 854 3729
rect 906 3677 978 3729
rect 1030 3677 1102 3729
rect 1154 3677 1226 3729
rect 1278 3677 1350 3729
rect 1402 3677 1474 3729
rect 1526 3677 1598 3729
rect 1650 3677 1722 3729
rect 1774 3677 1846 3729
rect 1898 3677 1970 3729
rect 2022 3677 2074 3729
rect 430 3605 2074 3677
rect 430 3553 482 3605
rect 534 3553 606 3605
rect 658 3553 730 3605
rect 782 3553 854 3605
rect 906 3553 978 3605
rect 1030 3553 1102 3605
rect 1154 3553 1226 3605
rect 1278 3553 1350 3605
rect 1402 3553 1474 3605
rect 1526 3553 1598 3605
rect 1650 3553 1722 3605
rect 1774 3553 1846 3605
rect 1898 3553 1970 3605
rect 2022 3553 2074 3605
rect 430 3481 2074 3553
rect 430 3429 482 3481
rect 534 3429 606 3481
rect 658 3429 730 3481
rect 782 3429 854 3481
rect 906 3429 978 3481
rect 1030 3429 1102 3481
rect 1154 3429 1226 3481
rect 1278 3429 1350 3481
rect 1402 3429 1474 3481
rect 1526 3429 1598 3481
rect 1650 3429 1722 3481
rect 1774 3429 1846 3481
rect 1898 3429 1970 3481
rect 2022 3429 2074 3481
rect 430 3357 2074 3429
rect 430 3305 482 3357
rect 534 3305 606 3357
rect 658 3305 730 3357
rect 782 3305 854 3357
rect 906 3305 978 3357
rect 1030 3305 1102 3357
rect 1154 3305 1226 3357
rect 1278 3305 1350 3357
rect 1402 3305 1474 3357
rect 1526 3305 1598 3357
rect 1650 3305 1722 3357
rect 1774 3305 1846 3357
rect 1898 3305 1970 3357
rect 2022 3305 2074 3357
rect 430 3233 2074 3305
rect 430 3181 482 3233
rect 534 3181 606 3233
rect 658 3181 730 3233
rect 782 3181 854 3233
rect 906 3181 978 3233
rect 1030 3181 1102 3233
rect 1154 3181 1226 3233
rect 1278 3181 1350 3233
rect 1402 3181 1474 3233
rect 1526 3181 1598 3233
rect 1650 3181 1722 3233
rect 1774 3181 1846 3233
rect 1898 3181 1970 3233
rect 2022 3181 2074 3233
rect 430 3109 2074 3181
rect 430 3057 482 3109
rect 534 3057 606 3109
rect 658 3057 730 3109
rect 782 3057 854 3109
rect 906 3057 978 3109
rect 1030 3057 1102 3109
rect 1154 3057 1226 3109
rect 1278 3057 1350 3109
rect 1402 3057 1474 3109
rect 1526 3057 1598 3109
rect 1650 3057 1722 3109
rect 1774 3057 1846 3109
rect 1898 3057 1970 3109
rect 2022 3057 2074 3109
rect 430 2985 2074 3057
rect 430 2933 482 2985
rect 534 2933 606 2985
rect 658 2933 730 2985
rect 782 2933 854 2985
rect 906 2933 978 2985
rect 1030 2933 1102 2985
rect 1154 2933 1226 2985
rect 1278 2933 1350 2985
rect 1402 2933 1474 2985
rect 1526 2933 1598 2985
rect 1650 2933 1722 2985
rect 1774 2933 1846 2985
rect 1898 2933 1970 2985
rect 2022 2933 2074 2985
rect 430 2861 2074 2933
rect 430 2809 482 2861
rect 534 2809 606 2861
rect 658 2809 730 2861
rect 782 2809 854 2861
rect 906 2809 978 2861
rect 1030 2809 1102 2861
rect 1154 2809 1226 2861
rect 1278 2809 1350 2861
rect 1402 2809 1474 2861
rect 1526 2809 1598 2861
rect 1650 2809 1722 2861
rect 1774 2809 1846 2861
rect 1898 2809 1970 2861
rect 2022 2809 2074 2861
rect 430 2737 2074 2809
rect 430 2685 482 2737
rect 534 2685 606 2737
rect 658 2685 730 2737
rect 782 2685 854 2737
rect 906 2685 978 2737
rect 1030 2685 1102 2737
rect 1154 2685 1226 2737
rect 1278 2685 1350 2737
rect 1402 2685 1474 2737
rect 1526 2685 1598 2737
rect 1650 2685 1722 2737
rect 1774 2685 1846 2737
rect 1898 2685 1970 2737
rect 2022 2685 2074 2737
rect 430 2613 2074 2685
rect 430 2561 482 2613
rect 534 2561 606 2613
rect 658 2561 730 2613
rect 782 2561 854 2613
rect 906 2561 978 2613
rect 1030 2561 1102 2613
rect 1154 2561 1226 2613
rect 1278 2561 1350 2613
rect 1402 2561 1474 2613
rect 1526 2561 1598 2613
rect 1650 2561 1722 2613
rect 1774 2561 1846 2613
rect 1898 2561 1970 2613
rect 2022 2561 2074 2613
rect 430 2489 2074 2561
rect 430 2437 482 2489
rect 534 2437 606 2489
rect 658 2437 730 2489
rect 782 2437 854 2489
rect 906 2437 978 2489
rect 1030 2437 1102 2489
rect 1154 2437 1226 2489
rect 1278 2437 1350 2489
rect 1402 2437 1474 2489
rect 1526 2437 1598 2489
rect 1650 2437 1722 2489
rect 1774 2437 1846 2489
rect 1898 2437 1970 2489
rect 2022 2437 2074 2489
rect 430 2365 2074 2437
rect 430 2313 482 2365
rect 534 2313 606 2365
rect 658 2313 730 2365
rect 782 2313 854 2365
rect 906 2313 978 2365
rect 1030 2313 1102 2365
rect 1154 2313 1226 2365
rect 1278 2313 1350 2365
rect 1402 2313 1474 2365
rect 1526 2313 1598 2365
rect 1650 2313 1722 2365
rect 1774 2313 1846 2365
rect 1898 2313 1970 2365
rect 2022 2313 2074 2365
rect 430 2241 2074 2313
rect 430 2189 482 2241
rect 534 2189 606 2241
rect 658 2189 730 2241
rect 782 2189 854 2241
rect 906 2189 978 2241
rect 1030 2189 1102 2241
rect 1154 2189 1226 2241
rect 1278 2189 1350 2241
rect 1402 2189 1474 2241
rect 1526 2189 1598 2241
rect 1650 2189 1722 2241
rect 1774 2189 1846 2241
rect 1898 2189 1970 2241
rect 2022 2189 2074 2241
rect 430 2117 2074 2189
rect 430 2065 482 2117
rect 534 2065 606 2117
rect 658 2065 730 2117
rect 782 2065 854 2117
rect 906 2065 978 2117
rect 1030 2065 1102 2117
rect 1154 2065 1226 2117
rect 1278 2065 1350 2117
rect 1402 2065 1474 2117
rect 1526 2065 1598 2117
rect 1650 2065 1722 2117
rect 1774 2065 1846 2117
rect 1898 2065 1970 2117
rect 2022 2065 2074 2117
rect 430 1993 2074 2065
rect 430 1941 482 1993
rect 534 1941 606 1993
rect 658 1941 730 1993
rect 782 1941 854 1993
rect 906 1941 978 1993
rect 1030 1941 1102 1993
rect 1154 1941 1226 1993
rect 1278 1941 1350 1993
rect 1402 1941 1474 1993
rect 1526 1941 1598 1993
rect 1650 1941 1722 1993
rect 1774 1941 1846 1993
rect 1898 1941 1970 1993
rect 2022 1941 2074 1993
rect 430 1869 2074 1941
rect 430 1817 482 1869
rect 534 1817 606 1869
rect 658 1817 730 1869
rect 782 1817 854 1869
rect 906 1817 978 1869
rect 1030 1817 1102 1869
rect 1154 1817 1226 1869
rect 1278 1817 1350 1869
rect 1402 1817 1474 1869
rect 1526 1817 1598 1869
rect 1650 1817 1722 1869
rect 1774 1817 1846 1869
rect 1898 1817 1970 1869
rect 2022 1817 2074 1869
rect 430 1745 2074 1817
rect 430 1693 482 1745
rect 534 1693 606 1745
rect 658 1693 730 1745
rect 782 1693 854 1745
rect 906 1693 978 1745
rect 1030 1693 1102 1745
rect 1154 1693 1226 1745
rect 1278 1693 1350 1745
rect 1402 1693 1474 1745
rect 1526 1693 1598 1745
rect 1650 1693 1722 1745
rect 1774 1693 1846 1745
rect 1898 1693 1970 1745
rect 2022 1693 2074 1745
rect 430 1621 2074 1693
rect 430 1569 482 1621
rect 534 1569 606 1621
rect 658 1569 730 1621
rect 782 1569 854 1621
rect 906 1569 978 1621
rect 1030 1569 1102 1621
rect 1154 1569 1226 1621
rect 1278 1569 1350 1621
rect 1402 1569 1474 1621
rect 1526 1569 1598 1621
rect 1650 1569 1722 1621
rect 1774 1569 1846 1621
rect 1898 1569 1970 1621
rect 2022 1569 2074 1621
rect 430 1497 2074 1569
rect 430 1445 482 1497
rect 534 1445 606 1497
rect 658 1445 730 1497
rect 782 1445 854 1497
rect 906 1445 978 1497
rect 1030 1445 1102 1497
rect 1154 1445 1226 1497
rect 1278 1445 1350 1497
rect 1402 1445 1474 1497
rect 1526 1445 1598 1497
rect 1650 1445 1722 1497
rect 1774 1445 1846 1497
rect 1898 1445 1970 1497
rect 2022 1445 2074 1497
rect 430 1373 2074 1445
rect 430 1321 482 1373
rect 534 1321 606 1373
rect 658 1321 730 1373
rect 782 1321 854 1373
rect 906 1321 978 1373
rect 1030 1321 1102 1373
rect 1154 1321 1226 1373
rect 1278 1321 1350 1373
rect 1402 1321 1474 1373
rect 1526 1321 1598 1373
rect 1650 1321 1722 1373
rect 1774 1321 1846 1373
rect 1898 1321 1970 1373
rect 2022 1321 2074 1373
rect 430 1249 2074 1321
rect 430 1197 482 1249
rect 534 1197 606 1249
rect 658 1197 730 1249
rect 782 1197 854 1249
rect 906 1197 978 1249
rect 1030 1197 1102 1249
rect 1154 1197 1226 1249
rect 1278 1197 1350 1249
rect 1402 1197 1474 1249
rect 1526 1197 1598 1249
rect 1650 1197 1722 1249
rect 1774 1197 1846 1249
rect 1898 1197 1970 1249
rect 2022 1197 2074 1249
rect 430 1125 2074 1197
rect 430 1073 482 1125
rect 534 1073 606 1125
rect 658 1073 730 1125
rect 782 1073 854 1125
rect 906 1073 978 1125
rect 1030 1073 1102 1125
rect 1154 1073 1226 1125
rect 1278 1073 1350 1125
rect 1402 1073 1474 1125
rect 1526 1073 1598 1125
rect 1650 1073 1722 1125
rect 1774 1073 1846 1125
rect 1898 1073 1970 1125
rect 2022 1073 2074 1125
rect 430 1001 2074 1073
rect 430 949 482 1001
rect 534 949 606 1001
rect 658 949 730 1001
rect 782 949 854 1001
rect 906 949 978 1001
rect 1030 949 1102 1001
rect 1154 949 1226 1001
rect 1278 949 1350 1001
rect 1402 949 1474 1001
rect 1526 949 1598 1001
rect 1650 949 1722 1001
rect 1774 949 1846 1001
rect 1898 949 1970 1001
rect 2022 949 2074 1001
rect 430 877 2074 949
rect 430 825 482 877
rect 534 825 606 877
rect 658 825 730 877
rect 782 825 854 877
rect 906 825 978 877
rect 1030 825 1102 877
rect 1154 825 1226 877
rect 1278 825 1350 877
rect 1402 825 1474 877
rect 1526 825 1598 877
rect 1650 825 1722 877
rect 1774 825 1846 877
rect 1898 825 1970 877
rect 2022 825 2074 877
rect 430 753 2074 825
rect 430 701 482 753
rect 534 701 606 753
rect 658 701 730 753
rect 782 701 854 753
rect 906 701 978 753
rect 1030 701 1102 753
rect 1154 701 1226 753
rect 1278 701 1350 753
rect 1402 701 1474 753
rect 1526 701 1598 753
rect 1650 701 1722 753
rect 1774 701 1846 753
rect 1898 701 1970 753
rect 2022 701 2074 753
rect 430 629 2074 701
rect 430 577 482 629
rect 534 577 606 629
rect 658 577 730 629
rect 782 577 854 629
rect 906 577 978 629
rect 1030 577 1102 629
rect 1154 577 1226 629
rect 1278 577 1350 629
rect 1402 577 1474 629
rect 1526 577 1598 629
rect 1650 577 1722 629
rect 1774 577 1846 629
rect 1898 577 1970 629
rect 2022 577 2074 629
rect 430 505 2074 577
rect 430 453 482 505
rect 534 453 606 505
rect 658 453 730 505
rect 782 453 854 505
rect 906 453 978 505
rect 1030 453 1102 505
rect 1154 453 1226 505
rect 1278 453 1350 505
rect 1402 453 1474 505
rect 1526 453 1598 505
rect 1650 453 1722 505
rect 1774 453 1846 505
rect 1898 453 1970 505
rect 2022 453 2074 505
rect 430 401 2074 453
<< via2 >>
rect 0 7581 160 7648
rect 0 7529 156 7581
rect 156 7529 160 7581
rect 0 7457 160 7529
rect 0 7405 156 7457
rect 156 7405 160 7457
rect 0 7333 160 7405
rect 0 7281 156 7333
rect 156 7281 160 7333
rect 0 7209 160 7281
rect 0 7157 156 7209
rect 156 7157 160 7209
rect 0 7085 160 7157
rect 0 7033 156 7085
rect 156 7033 160 7085
rect 0 6961 160 7033
rect 0 6909 156 6961
rect 156 6909 160 6961
rect 0 6837 160 6909
rect 0 6785 156 6837
rect 156 6785 160 6837
rect 0 6713 160 6785
rect 0 6661 156 6713
rect 156 6661 160 6713
rect 0 6589 160 6661
rect 0 6537 156 6589
rect 156 6537 160 6589
rect 0 6465 160 6537
rect 0 6413 156 6465
rect 156 6413 160 6465
rect 0 6341 160 6413
rect 0 6289 156 6341
rect 156 6289 160 6341
rect 0 6217 160 6289
rect 0 6165 156 6217
rect 156 6165 160 6217
rect 0 6093 160 6165
rect 0 6041 156 6093
rect 156 6041 160 6093
rect 0 6032 160 6041
rect 0 4977 160 5047
rect 0 4925 156 4977
rect 156 4925 160 4977
rect 0 4853 160 4925
rect 0 4801 156 4853
rect 156 4801 160 4853
rect 0 4729 160 4801
rect 0 4677 156 4729
rect 156 4677 160 4729
rect 0 4605 160 4677
rect 0 4553 156 4605
rect 156 4553 160 4605
rect 0 4481 160 4553
rect 0 4429 156 4481
rect 156 4429 160 4481
rect 0 4357 160 4429
rect 0 4305 156 4357
rect 156 4305 160 4357
rect 0 4233 160 4305
rect 0 4181 156 4233
rect 156 4181 160 4233
rect 0 4109 160 4181
rect 0 4057 156 4109
rect 156 4057 160 4109
rect 0 3985 160 4057
rect 0 3933 156 3985
rect 156 3933 160 3985
rect 0 3861 160 3933
rect 0 3809 156 3861
rect 156 3809 160 3861
rect 0 3737 160 3809
rect 0 3685 156 3737
rect 156 3685 160 3737
rect 0 3613 160 3685
rect 0 3561 156 3613
rect 156 3561 160 3613
rect 0 3489 160 3561
rect 0 3437 156 3489
rect 156 3437 160 3489
rect 0 3365 160 3437
rect 0 3313 156 3365
rect 156 3313 160 3365
rect 0 3241 160 3313
rect 0 3189 156 3241
rect 156 3189 160 3241
rect 0 3117 160 3189
rect 0 3065 156 3117
rect 156 3065 160 3117
rect 0 2993 160 3065
rect 0 2941 156 2993
rect 156 2941 160 2993
rect 0 2911 160 2941
rect 0 1949 156 1992
rect 156 1949 160 1992
rect 0 1877 160 1949
rect 0 1825 156 1877
rect 156 1825 160 1877
rect 0 1753 160 1825
rect 0 1701 156 1753
rect 156 1701 160 1753
rect 0 1629 160 1701
rect 0 1577 156 1629
rect 156 1577 160 1629
rect 0 1505 160 1577
rect 0 1453 156 1505
rect 156 1453 160 1505
rect 0 1381 160 1453
rect 0 1329 156 1381
rect 156 1329 160 1381
rect 0 1257 160 1329
rect 0 1205 156 1257
rect 156 1205 160 1257
rect 0 1133 160 1205
rect 0 1081 156 1133
rect 156 1081 160 1133
rect 0 1009 160 1081
rect 0 957 156 1009
rect 156 957 160 1009
rect 0 885 160 957
rect 0 833 156 885
rect 156 833 160 885
rect 0 761 160 833
rect 0 709 156 761
rect 156 709 160 761
rect 0 688 160 709
<< metal3 >>
rect -10 7648 170 7658
rect -10 6032 0 7648
rect 160 6032 170 7648
rect -10 6022 170 6032
rect -10 5047 170 5057
rect -10 2911 0 5047
rect 160 2911 170 5047
rect -10 2901 170 2911
rect -10 1992 170 2002
rect -10 688 0 1992
rect 160 688 170 1992
rect -10 678 170 688
<< end >>
