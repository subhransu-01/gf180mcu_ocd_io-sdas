magic
tech gf180mcuD
magscale 1 10
timestamp 1764349902
<< isosubstrate >>
rect 251 53100 14727 57210
rect 2457 47106 12521 53100
rect 601 43110 14377 47106
rect 957 26495 12844 43110
rect 957 1096 14021 26495
<< nwell >>
rect 2457 52160 12521 52716
rect 2457 48116 3008 52160
rect 11970 48116 12521 52160
rect 2457 47560 12521 48116
<< pwell >>
rect 747 53655 3923 56655
rect 4183 53655 7359 56655
rect 7619 53655 10795 56655
rect 11055 53655 14231 56655
<< mvndiff >>
rect 747 56618 835 56655
rect 747 53692 760 56618
rect 806 53692 835 56618
rect 747 53655 835 53692
rect 3835 56618 3923 56655
rect 3835 53692 3864 56618
rect 3910 53692 3923 56618
rect 3835 53655 3923 53692
rect 4183 56618 4271 56655
rect 4183 53692 4196 56618
rect 4242 53692 4271 56618
rect 4183 53655 4271 53692
rect 7271 56618 7359 56655
rect 7271 53692 7300 56618
rect 7346 53692 7359 56618
rect 7271 53655 7359 53692
rect 7619 56618 7707 56655
rect 7619 53692 7632 56618
rect 7678 53692 7707 56618
rect 7619 53655 7707 53692
rect 10707 56618 10795 56655
rect 10707 53692 10736 56618
rect 10782 53692 10795 56618
rect 10707 53655 10795 53692
rect 11055 56618 11143 56655
rect 11055 53692 11068 56618
rect 11114 53692 11143 56618
rect 11055 53655 11143 53692
rect 14143 56618 14231 56655
rect 14143 53692 14172 56618
rect 14218 53692 14231 56618
rect 14143 53655 14231 53692
<< mvndiffc >>
rect 760 53692 806 56618
rect 3864 53692 3910 56618
rect 4196 53692 4242 56618
rect 7300 53692 7346 56618
rect 7632 53692 7678 56618
rect 10736 53692 10782 56618
rect 11068 53692 11114 56618
rect 14172 53692 14218 56618
<< psubdiff >>
rect 334 57105 14644 57127
rect 334 53205 356 57105
rect 402 57059 510 57105
rect 14468 57059 14576 57105
rect 402 57037 14576 57059
rect 402 53273 424 57037
rect 14554 53273 14576 57037
rect 402 53251 14576 53273
rect 402 53205 510 53251
rect 14468 53205 14576 53251
rect 14622 53205 14644 57105
rect 334 53183 14644 53205
rect 246 52611 2236 52633
rect 246 47665 268 52611
rect 2214 47665 2236 52611
rect 246 47643 2236 47665
rect 3094 52029 11884 52051
rect 3094 51983 3142 52029
rect 11836 51983 11884 52029
rect 3094 51900 11884 51983
rect 3094 48376 3116 51900
rect 3162 51875 11816 51900
rect 3162 51844 3424 51875
rect 3162 51234 3270 51844
rect 3316 51829 3424 51844
rect 11554 51844 11816 51875
rect 11554 51829 11662 51844
rect 3316 51807 11662 51829
rect 3316 51271 3338 51807
rect 11640 51271 11662 51807
rect 3316 51249 11662 51271
rect 3316 51234 3424 51249
rect 3162 51203 3424 51234
rect 11554 51234 11662 51249
rect 11708 51234 11816 51844
rect 11554 51203 11816 51234
rect 3162 51095 11816 51203
rect 3162 51049 3330 51095
rect 11648 51049 11816 51095
rect 3162 50941 11816 51049
rect 3162 50910 3424 50941
rect 3162 50300 3270 50910
rect 3316 50895 3424 50910
rect 11554 50910 11816 50941
rect 11554 50895 11662 50910
rect 3316 50873 11662 50895
rect 3316 50337 3338 50873
rect 11640 50337 11662 50873
rect 3316 50315 11662 50337
rect 3316 50300 3424 50315
rect 3162 50269 3424 50300
rect 11554 50300 11662 50315
rect 11708 50300 11816 50910
rect 11554 50269 11816 50300
rect 3162 50161 11816 50269
rect 3162 50115 3330 50161
rect 11648 50115 11816 50161
rect 3162 50007 11816 50115
rect 3162 49976 3424 50007
rect 3162 49366 3270 49976
rect 3316 49961 3424 49976
rect 11554 49976 11816 50007
rect 11554 49961 11662 49976
rect 3316 49939 11662 49961
rect 3316 49403 3338 49939
rect 11640 49403 11662 49939
rect 3316 49381 11662 49403
rect 3316 49366 3424 49381
rect 3162 49335 3424 49366
rect 11554 49366 11662 49381
rect 11708 49366 11816 49976
rect 11554 49335 11816 49366
rect 3162 49227 11816 49335
rect 3162 49181 3330 49227
rect 11648 49181 11816 49227
rect 3162 49073 11816 49181
rect 3162 49042 3424 49073
rect 3162 48432 3270 49042
rect 3316 49027 3424 49042
rect 11554 49042 11816 49073
rect 11554 49027 11662 49042
rect 3316 49005 11662 49027
rect 3316 48469 3338 49005
rect 11640 48469 11662 49005
rect 3316 48447 11662 48469
rect 3316 48432 3424 48447
rect 3162 48401 3424 48432
rect 11554 48432 11662 48447
rect 11708 48432 11816 49042
rect 11554 48401 11816 48432
rect 3162 48376 11816 48401
rect 11862 48376 11884 51900
rect 3094 48293 11884 48376
rect 3094 48247 3142 48293
rect 11836 48247 11884 48293
rect 3094 48225 11884 48247
rect 12742 52611 14732 52633
rect 12742 47665 12764 52611
rect 14710 47665 14732 52611
rect 12742 47643 14732 47665
rect 246 42647 736 42669
rect 246 1201 268 42647
rect 714 1201 736 42647
rect 13001 42647 13991 42669
rect 13001 27201 13023 42647
rect 13969 27201 13991 42647
rect 13001 27179 13991 27201
rect 14242 42647 14732 42669
rect 246 1179 736 1201
rect 14242 1201 14264 42647
rect 14710 1201 14732 42647
rect 14242 1179 14732 1201
<< nsubdiff >>
rect 2540 52611 12438 52633
rect 2540 47665 2562 52611
rect 2908 52265 3016 52611
rect 11962 52265 12070 52611
rect 2908 52243 12070 52265
rect 2908 48033 2930 52243
rect 12048 48033 12070 52243
rect 2908 48011 12070 48033
rect 2908 47665 3016 48011
rect 11962 47665 12070 48011
rect 12416 47665 12438 52611
rect 2540 47643 12438 47665
<< psubdiffcont >>
rect 356 53205 402 57105
rect 510 57059 14468 57105
rect 510 53205 14468 53251
rect 14576 53205 14622 57105
rect 268 47665 2214 52611
rect 3142 51983 11836 52029
rect 3116 48376 3162 51900
rect 3270 51234 3316 51844
rect 3424 51829 11554 51875
rect 3424 51203 11554 51249
rect 11662 51234 11708 51844
rect 3330 51049 11648 51095
rect 3270 50300 3316 50910
rect 3424 50895 11554 50941
rect 3424 50269 11554 50315
rect 11662 50300 11708 50910
rect 3330 50115 11648 50161
rect 3270 49366 3316 49976
rect 3424 49961 11554 50007
rect 3424 49335 11554 49381
rect 11662 49366 11708 49976
rect 3330 49181 11648 49227
rect 3270 48432 3316 49042
rect 3424 49027 11554 49073
rect 3424 48401 11554 48447
rect 11662 48432 11708 49042
rect 11816 48376 11862 51900
rect 3142 48247 11836 48293
rect 12764 47665 14710 52611
rect 268 1201 714 42647
rect 13023 27201 13969 42647
rect 14264 1201 14710 42647
<< nsubdiffcont >>
rect 2562 47665 2908 52611
rect 3016 52265 11962 52611
rect 3016 47665 11962 48011
rect 12070 47665 12416 52611
<< mvnmoscap >>
rect 835 53655 3835 56655
rect 4271 53655 7271 56655
rect 7707 53655 10707 56655
rect 11143 53655 14143 56655
<< polysilicon >>
rect 835 56734 3835 56747
rect 835 56688 888 56734
rect 3782 56688 3835 56734
rect 835 56655 3835 56688
rect 4271 56734 7271 56747
rect 4271 56688 4324 56734
rect 7218 56688 7271 56734
rect 4271 56655 7271 56688
rect 7707 56734 10707 56747
rect 7707 56688 7760 56734
rect 10654 56688 10707 56734
rect 7707 56655 10707 56688
rect 11143 56734 14143 56747
rect 11143 56688 11196 56734
rect 14090 56688 14143 56734
rect 11143 56655 14143 56688
rect 835 53622 3835 53655
rect 835 53576 888 53622
rect 3782 53576 3835 53622
rect 835 53563 3835 53576
rect 4271 53622 7271 53655
rect 4271 53576 4324 53622
rect 7218 53576 7271 53622
rect 4271 53563 7271 53576
rect 7707 53622 10707 53655
rect 7707 53576 7760 53622
rect 10654 53576 10707 53622
rect 7707 53563 10707 53576
rect 11143 53622 14143 53655
rect 11143 53576 11196 53622
rect 14090 53576 14143 53622
rect 11143 53563 14143 53576
<< polycontact >>
rect 888 56688 3782 56734
rect 4324 56688 7218 56734
rect 7760 56688 10654 56734
rect 11196 56688 14090 56734
rect 888 53576 3782 53622
rect 4324 53576 7218 53622
rect 7760 53576 10654 53622
rect 11196 53576 14090 53622
<< mvndiode >>
rect 3489 51626 11489 51639
rect 3489 51580 3502 51626
rect 11476 51580 11489 51626
rect 3489 51498 11489 51580
rect 3489 51452 3502 51498
rect 11476 51452 11489 51498
rect 3489 51439 11489 51452
rect 3489 50692 11489 50705
rect 3489 50646 3502 50692
rect 11476 50646 11489 50692
rect 3489 50564 11489 50646
rect 3489 50518 3502 50564
rect 11476 50518 11489 50564
rect 3489 50505 11489 50518
rect 3489 49758 11489 49771
rect 3489 49712 3502 49758
rect 11476 49712 11489 49758
rect 3489 49630 11489 49712
rect 3489 49584 3502 49630
rect 11476 49584 11489 49630
rect 3489 49571 11489 49584
rect 3489 48824 11489 48837
rect 3489 48778 3502 48824
rect 11476 48778 11489 48824
rect 3489 48696 11489 48778
rect 3489 48650 3502 48696
rect 11476 48650 11489 48696
rect 3489 48637 11489 48650
<< mvndiodec >>
rect 3502 51580 11476 51626
rect 3502 51452 11476 51498
rect 3502 50646 11476 50692
rect 3502 50518 11476 50564
rect 3502 49712 11476 49758
rect 3502 49584 11476 49630
rect 3502 48778 11476 48824
rect 3502 48650 11476 48696
<< metal1 >>
rect 10 57259 86 57271
rect 10 57207 22 57259
rect 74 57207 86 57259
rect 10 57151 86 57207
rect 10 57099 22 57151
rect 74 57099 86 57151
rect 14892 57259 14968 57271
rect 14892 57207 14904 57259
rect 14956 57207 14968 57259
rect 14892 57151 14968 57207
rect 10 57043 86 57099
rect 10 56991 22 57043
rect 74 56991 86 57043
rect 10 56935 86 56991
rect 10 56883 22 56935
rect 74 56883 86 56935
rect 10 56827 86 56883
rect 10 56775 22 56827
rect 74 56775 86 56827
rect 10 56719 86 56775
rect 10 56667 22 56719
rect 74 56667 86 56719
rect 10 56611 86 56667
rect 10 56559 22 56611
rect 74 56559 86 56611
rect 10 56503 86 56559
rect 10 56451 22 56503
rect 74 56451 86 56503
rect 10 56395 86 56451
rect 10 56343 22 56395
rect 74 56343 86 56395
rect 10 56287 86 56343
rect 10 56235 22 56287
rect 74 56235 86 56287
rect 10 56179 86 56235
rect 10 56127 22 56179
rect 74 56127 86 56179
rect 10 56071 86 56127
rect 10 56019 22 56071
rect 74 56019 86 56071
rect 10 56007 86 56019
rect 345 57105 14633 57116
rect 10 54174 86 54186
rect 10 54122 22 54174
rect 74 54122 86 54174
rect 10 54066 86 54122
rect 10 54014 22 54066
rect 74 54014 86 54066
rect 10 53958 86 54014
rect 10 53906 22 53958
rect 74 53906 86 53958
rect 10 53850 86 53906
rect 10 53798 22 53850
rect 74 53798 86 53850
rect 10 53742 86 53798
rect 10 53690 22 53742
rect 74 53690 86 53742
rect 10 53634 86 53690
rect 10 53582 22 53634
rect 74 53582 86 53634
rect 10 53526 86 53582
rect 10 53474 22 53526
rect 74 53474 86 53526
rect 10 53418 86 53474
rect 10 53366 22 53418
rect 74 53366 86 53418
rect 10 53310 86 53366
rect 10 53258 22 53310
rect 74 53258 86 53310
rect 10 53202 86 53258
rect 10 53150 22 53202
rect 74 53150 86 53202
rect 345 53205 356 57105
rect 402 57104 510 57105
rect 14468 57104 14576 57105
rect 427 57052 483 57104
rect 535 57052 591 57059
rect 643 57052 699 57059
rect 751 57052 807 57059
rect 859 57052 915 57059
rect 967 57052 1023 57059
rect 1075 57052 1131 57059
rect 1183 57052 1239 57059
rect 1291 57052 1347 57059
rect 1399 57052 1455 57059
rect 1507 57052 1563 57059
rect 1615 57052 1671 57059
rect 1723 57052 1779 57059
rect 1831 57052 1887 57059
rect 1939 57052 1995 57059
rect 2047 57052 2768 57059
rect 2820 57052 2876 57059
rect 2928 57052 2984 57059
rect 3036 57052 3092 57059
rect 3144 57052 3200 57059
rect 3252 57052 3308 57059
rect 3360 57052 3416 57059
rect 3468 57052 3524 57059
rect 3576 57052 3632 57059
rect 3684 57052 3740 57059
rect 3792 57052 3848 57059
rect 3900 57052 3956 57059
rect 4008 57052 4064 57059
rect 4116 57052 4172 57059
rect 4224 57052 4280 57059
rect 4332 57052 4388 57059
rect 4440 57052 4496 57059
rect 4548 57052 4604 57059
rect 4656 57052 4712 57059
rect 4764 57052 5138 57059
rect 5190 57052 5246 57059
rect 5298 57052 5354 57059
rect 5406 57052 5462 57059
rect 5514 57052 5570 57059
rect 5622 57052 5678 57059
rect 5730 57052 5786 57059
rect 5838 57052 5894 57059
rect 5946 57052 6002 57059
rect 6054 57052 6110 57059
rect 6162 57052 6218 57059
rect 6270 57052 6326 57059
rect 6378 57052 6434 57059
rect 6486 57052 6542 57059
rect 6594 57052 6650 57059
rect 6702 57052 6758 57059
rect 6810 57052 6866 57059
rect 6918 57052 6974 57059
rect 7026 57052 7082 57059
rect 7134 57052 7844 57059
rect 7896 57052 7952 57059
rect 8004 57052 8060 57059
rect 8112 57052 8168 57059
rect 8220 57052 8276 57059
rect 8328 57052 8384 57059
rect 8436 57052 8492 57059
rect 8544 57052 8600 57059
rect 8652 57052 8708 57059
rect 8760 57052 8816 57059
rect 8868 57052 8924 57059
rect 8976 57052 9032 57059
rect 9084 57052 9140 57059
rect 9192 57052 9248 57059
rect 9300 57052 9356 57059
rect 9408 57052 9464 57059
rect 9516 57052 9572 57059
rect 9624 57052 9680 57059
rect 9732 57052 9788 57059
rect 9840 57052 10214 57059
rect 10266 57052 10322 57059
rect 10374 57052 10430 57059
rect 10482 57052 10538 57059
rect 10590 57052 10646 57059
rect 10698 57052 10754 57059
rect 10806 57052 10862 57059
rect 10914 57052 10970 57059
rect 11022 57052 11078 57059
rect 11130 57052 11186 57059
rect 11238 57052 11294 57059
rect 11346 57052 11402 57059
rect 11454 57052 11510 57059
rect 11562 57052 11618 57059
rect 11670 57052 11726 57059
rect 11778 57052 11834 57059
rect 11886 57052 11942 57059
rect 11994 57052 12050 57059
rect 12102 57052 12158 57059
rect 12210 57052 12931 57059
rect 12983 57052 13039 57059
rect 13091 57052 13147 57059
rect 13199 57052 13255 57059
rect 13307 57052 13363 57059
rect 13415 57052 13471 57059
rect 13523 57052 13579 57059
rect 13631 57052 13687 57059
rect 13739 57052 13795 57059
rect 13847 57052 13903 57059
rect 13955 57052 14011 57059
rect 14063 57052 14119 57059
rect 14171 57052 14227 57059
rect 14279 57052 14335 57059
rect 14387 57052 14443 57059
rect 14495 57052 14551 57104
rect 402 57048 14576 57052
rect 402 57040 2059 57048
rect 2756 57040 4776 57048
rect 5126 57040 7146 57048
rect 7832 57040 9852 57048
rect 10202 57040 12222 57048
rect 12919 57040 14576 57048
rect 402 56655 413 57040
rect 2489 56745 2673 56753
rect 12305 56745 12489 56753
rect 877 56741 3793 56745
rect 877 56734 2501 56741
rect 2553 56734 2609 56741
rect 2661 56734 3793 56741
rect 877 56688 888 56734
rect 3782 56688 3793 56734
rect 877 56677 3793 56688
rect 402 56643 817 56655
rect 421 56591 493 56643
rect 545 56591 617 56643
rect 669 56591 741 56643
rect 793 56618 817 56643
rect 402 56519 760 56591
rect 421 56467 493 56519
rect 545 56467 617 56519
rect 669 56467 741 56519
rect 402 56395 760 56467
rect 421 56343 493 56395
rect 545 56343 617 56395
rect 669 56343 741 56395
rect 402 56271 760 56343
rect 421 56219 493 56271
rect 545 56219 617 56271
rect 669 56219 741 56271
rect 402 56147 760 56219
rect 421 56095 493 56147
rect 545 56095 617 56147
rect 669 56095 741 56147
rect 402 56023 760 56095
rect 421 55971 493 56023
rect 545 55971 617 56023
rect 669 55971 741 56023
rect 402 55899 760 55971
rect 421 55847 493 55899
rect 545 55847 617 55899
rect 669 55847 741 55899
rect 402 55775 760 55847
rect 421 55723 493 55775
rect 545 55723 617 55775
rect 669 55723 741 55775
rect 402 55651 760 55723
rect 421 55599 493 55651
rect 545 55599 617 55651
rect 669 55599 741 55651
rect 402 55527 760 55599
rect 421 55475 493 55527
rect 545 55475 617 55527
rect 669 55475 741 55527
rect 402 55403 760 55475
rect 421 55351 493 55403
rect 545 55351 617 55403
rect 669 55351 741 55403
rect 402 55279 760 55351
rect 421 55227 493 55279
rect 545 55227 617 55279
rect 669 55227 741 55279
rect 402 55155 760 55227
rect 421 55103 493 55155
rect 545 55103 617 55155
rect 669 55103 741 55155
rect 402 55031 760 55103
rect 421 54979 493 55031
rect 545 54979 617 55031
rect 669 54979 741 55031
rect 402 54907 760 54979
rect 421 54855 493 54907
rect 545 54855 617 54907
rect 669 54855 741 54907
rect 402 54783 760 54855
rect 421 54731 493 54783
rect 545 54731 617 54783
rect 669 54731 741 54783
rect 402 54659 760 54731
rect 421 54607 493 54659
rect 545 54607 617 54659
rect 669 54607 741 54659
rect 402 54535 760 54607
rect 421 54483 493 54535
rect 545 54483 617 54535
rect 669 54483 741 54535
rect 402 54411 760 54483
rect 421 54359 493 54411
rect 545 54359 617 54411
rect 669 54359 741 54411
rect 402 54287 760 54359
rect 421 54235 493 54287
rect 545 54235 617 54287
rect 669 54235 741 54287
rect 402 54163 760 54235
rect 421 54111 493 54163
rect 545 54111 617 54163
rect 669 54111 741 54163
rect 402 54039 760 54111
rect 421 53987 493 54039
rect 545 53987 617 54039
rect 669 53987 741 54039
rect 402 53915 760 53987
rect 421 53863 493 53915
rect 545 53863 617 53915
rect 669 53863 741 53915
rect 402 53791 760 53863
rect 421 53739 493 53791
rect 545 53739 617 53791
rect 669 53739 741 53791
rect 402 53692 760 53739
rect 806 53692 817 56618
rect 402 53667 817 53692
rect 421 53615 493 53667
rect 545 53615 617 53667
rect 669 53615 741 53667
rect 793 53615 817 53667
rect 402 53543 817 53615
rect 877 53633 1877 56677
rect 2793 53633 3793 56677
rect 4313 56734 7229 56745
rect 4313 56688 4324 56734
rect 7218 56688 7229 56734
rect 877 53622 3793 53633
rect 877 53576 888 53622
rect 3782 53576 3793 53622
rect 877 53569 2501 53576
rect 2553 53569 2609 53576
rect 2661 53569 3793 53576
rect 877 53565 3793 53569
rect 3853 56643 4253 56655
rect 3853 56618 3903 56643
rect 3853 53692 3864 56618
rect 3955 56591 4027 56643
rect 4079 56591 4151 56643
rect 4203 56618 4253 56643
rect 3910 56519 4196 56591
rect 3955 56467 4027 56519
rect 4079 56467 4151 56519
rect 3910 56395 4196 56467
rect 3955 56343 4027 56395
rect 4079 56343 4151 56395
rect 3910 56271 4196 56343
rect 3955 56219 4027 56271
rect 4079 56219 4151 56271
rect 3910 56147 4196 56219
rect 3955 56095 4027 56147
rect 4079 56095 4151 56147
rect 3910 56023 4196 56095
rect 3955 55971 4027 56023
rect 4079 55971 4151 56023
rect 3910 55899 4196 55971
rect 3955 55847 4027 55899
rect 4079 55847 4151 55899
rect 3910 55775 4196 55847
rect 3955 55723 4027 55775
rect 4079 55723 4151 55775
rect 3910 55651 4196 55723
rect 3955 55599 4027 55651
rect 4079 55599 4151 55651
rect 3910 55527 4196 55599
rect 3955 55475 4027 55527
rect 4079 55475 4151 55527
rect 3910 55403 4196 55475
rect 3955 55351 4027 55403
rect 4079 55351 4151 55403
rect 3910 55279 4196 55351
rect 3955 55227 4027 55279
rect 4079 55227 4151 55279
rect 3910 55155 4196 55227
rect 3955 55103 4027 55155
rect 4079 55103 4151 55155
rect 3910 55031 4196 55103
rect 3955 54979 4027 55031
rect 4079 54979 4151 55031
rect 3910 54907 4196 54979
rect 3955 54855 4027 54907
rect 4079 54855 4151 54907
rect 3910 54783 4196 54855
rect 3955 54731 4027 54783
rect 4079 54731 4151 54783
rect 3910 54659 4196 54731
rect 3955 54607 4027 54659
rect 4079 54607 4151 54659
rect 3910 54535 4196 54607
rect 3955 54483 4027 54535
rect 4079 54483 4151 54535
rect 3910 54411 4196 54483
rect 3955 54359 4027 54411
rect 4079 54359 4151 54411
rect 3910 54287 4196 54359
rect 3955 54235 4027 54287
rect 4079 54235 4151 54287
rect 3910 54163 4196 54235
rect 3955 54111 4027 54163
rect 4079 54111 4151 54163
rect 3910 54039 4196 54111
rect 3955 53987 4027 54039
rect 4079 53987 4151 54039
rect 3910 53915 4196 53987
rect 3955 53863 4027 53915
rect 4079 53863 4151 53915
rect 3910 53791 4196 53863
rect 3955 53739 4027 53791
rect 4079 53739 4151 53791
rect 3910 53692 4196 53739
rect 4242 53692 4253 56618
rect 3853 53667 4253 53692
rect 3853 53615 3903 53667
rect 3955 53615 4027 53667
rect 4079 53615 4151 53667
rect 4203 53615 4253 53667
rect 2489 53557 2673 53565
rect 421 53491 493 53543
rect 545 53491 617 53543
rect 669 53491 741 53543
rect 793 53505 817 53543
rect 3853 53543 4253 53615
rect 4313 56641 4871 56688
rect 4923 56641 4979 56688
rect 5031 56677 7229 56688
rect 5031 56641 5313 56677
rect 4313 56585 5313 56641
rect 4313 56533 4871 56585
rect 4923 56533 4979 56585
rect 5031 56533 5313 56585
rect 4313 56477 5313 56533
rect 4313 56425 4871 56477
rect 4923 56425 4979 56477
rect 5031 56425 5313 56477
rect 4313 56369 5313 56425
rect 4313 56317 4871 56369
rect 4923 56317 4979 56369
rect 5031 56317 5313 56369
rect 4313 56261 5313 56317
rect 4313 56209 4871 56261
rect 4923 56209 4979 56261
rect 5031 56209 5313 56261
rect 4313 56153 5313 56209
rect 4313 56101 4871 56153
rect 4923 56101 4979 56153
rect 5031 56101 5313 56153
rect 4313 56045 5313 56101
rect 4313 55993 4871 56045
rect 4923 55993 4979 56045
rect 5031 55993 5313 56045
rect 4313 55937 5313 55993
rect 4313 55885 4871 55937
rect 4923 55885 4979 55937
rect 5031 55885 5313 55937
rect 4313 55829 5313 55885
rect 4313 55777 4871 55829
rect 4923 55777 4979 55829
rect 5031 55777 5313 55829
rect 4313 55721 5313 55777
rect 4313 55669 4871 55721
rect 4923 55669 4979 55721
rect 5031 55669 5313 55721
rect 4313 55613 5313 55669
rect 4313 55561 4871 55613
rect 4923 55561 4979 55613
rect 5031 55561 5313 55613
rect 4313 55505 5313 55561
rect 4313 55453 4871 55505
rect 4923 55453 4979 55505
rect 5031 55453 5313 55505
rect 4313 55397 5313 55453
rect 4313 55345 4871 55397
rect 4923 55345 4979 55397
rect 5031 55345 5313 55397
rect 4313 55289 5313 55345
rect 4313 55237 4871 55289
rect 4923 55237 4979 55289
rect 5031 55237 5313 55289
rect 4313 55181 5313 55237
rect 4313 55129 4871 55181
rect 4923 55129 4979 55181
rect 5031 55129 5313 55181
rect 4313 55073 5313 55129
rect 4313 55021 4871 55073
rect 4923 55021 4979 55073
rect 5031 55021 5313 55073
rect 4313 54965 5313 55021
rect 4313 54913 4871 54965
rect 4923 54913 4979 54965
rect 5031 54913 5313 54965
rect 4313 54857 5313 54913
rect 4313 54805 4871 54857
rect 4923 54805 4979 54857
rect 5031 54805 5313 54857
rect 4313 54749 5313 54805
rect 4313 54697 4871 54749
rect 4923 54697 4979 54749
rect 5031 54697 5313 54749
rect 4313 54641 5313 54697
rect 4313 54589 4871 54641
rect 4923 54589 4979 54641
rect 5031 54589 5313 54641
rect 4313 54533 5313 54589
rect 4313 54481 4871 54533
rect 4923 54481 4979 54533
rect 5031 54481 5313 54533
rect 4313 54425 5313 54481
rect 4313 54373 4871 54425
rect 4923 54373 4979 54425
rect 5031 54373 5313 54425
rect 4313 54317 5313 54373
rect 4313 54265 4871 54317
rect 4923 54265 4979 54317
rect 5031 54265 5313 54317
rect 4313 54209 5313 54265
rect 4313 54157 4871 54209
rect 4923 54157 4979 54209
rect 5031 54157 5313 54209
rect 4313 54101 5313 54157
rect 4313 54049 4871 54101
rect 4923 54049 4979 54101
rect 5031 54049 5313 54101
rect 4313 53993 5313 54049
rect 4313 53941 4871 53993
rect 4923 53941 4979 53993
rect 5031 53941 5313 53993
rect 4313 53885 5313 53941
rect 4313 53833 4871 53885
rect 4923 53833 4979 53885
rect 5031 53833 5313 53885
rect 4313 53777 5313 53833
rect 4313 53725 4871 53777
rect 4923 53725 4979 53777
rect 5031 53725 5313 53777
rect 4313 53669 5313 53725
rect 4313 53622 4871 53669
rect 4923 53622 4979 53669
rect 5031 53633 5313 53669
rect 6229 53633 7229 56677
rect 7749 56734 10665 56745
rect 7749 56688 7760 56734
rect 10654 56688 10665 56734
rect 7749 56677 9947 56688
rect 5031 53622 7229 53633
rect 4313 53576 4324 53622
rect 7218 53576 7229 53622
rect 4313 53565 7229 53576
rect 7289 56618 7689 56655
rect 7289 53692 7300 56618
rect 7346 53692 7632 56618
rect 7678 53692 7689 56618
rect 3853 53505 3903 53543
rect 793 53491 3903 53505
rect 3955 53491 4027 53543
rect 4079 53491 4151 53543
rect 4203 53505 4253 53543
rect 7289 53505 7689 53692
rect 7749 53633 8749 56677
rect 9665 56641 9947 56677
rect 9999 56641 10055 56688
rect 10107 56641 10665 56688
rect 11185 56741 14101 56745
rect 11185 56734 12317 56741
rect 12369 56734 12425 56741
rect 12477 56734 14101 56741
rect 11185 56688 11196 56734
rect 14090 56688 14101 56734
rect 11185 56677 14101 56688
rect 9665 56585 10665 56641
rect 9665 56533 9947 56585
rect 9999 56533 10055 56585
rect 10107 56533 10665 56585
rect 9665 56477 10665 56533
rect 9665 56425 9947 56477
rect 9999 56425 10055 56477
rect 10107 56425 10665 56477
rect 9665 56369 10665 56425
rect 9665 56317 9947 56369
rect 9999 56317 10055 56369
rect 10107 56317 10665 56369
rect 9665 56261 10665 56317
rect 9665 56209 9947 56261
rect 9999 56209 10055 56261
rect 10107 56209 10665 56261
rect 9665 56153 10665 56209
rect 9665 56101 9947 56153
rect 9999 56101 10055 56153
rect 10107 56101 10665 56153
rect 9665 56045 10665 56101
rect 9665 55993 9947 56045
rect 9999 55993 10055 56045
rect 10107 55993 10665 56045
rect 9665 55937 10665 55993
rect 9665 55885 9947 55937
rect 9999 55885 10055 55937
rect 10107 55885 10665 55937
rect 9665 55829 10665 55885
rect 9665 55777 9947 55829
rect 9999 55777 10055 55829
rect 10107 55777 10665 55829
rect 9665 55721 10665 55777
rect 9665 55669 9947 55721
rect 9999 55669 10055 55721
rect 10107 55669 10665 55721
rect 9665 55613 10665 55669
rect 9665 55561 9947 55613
rect 9999 55561 10055 55613
rect 10107 55561 10665 55613
rect 9665 55505 10665 55561
rect 9665 55453 9947 55505
rect 9999 55453 10055 55505
rect 10107 55453 10665 55505
rect 9665 55397 10665 55453
rect 9665 55345 9947 55397
rect 9999 55345 10055 55397
rect 10107 55345 10665 55397
rect 9665 55289 10665 55345
rect 9665 55237 9947 55289
rect 9999 55237 10055 55289
rect 10107 55237 10665 55289
rect 9665 55181 10665 55237
rect 9665 55129 9947 55181
rect 9999 55129 10055 55181
rect 10107 55129 10665 55181
rect 9665 55073 10665 55129
rect 9665 55021 9947 55073
rect 9999 55021 10055 55073
rect 10107 55021 10665 55073
rect 9665 54965 10665 55021
rect 9665 54913 9947 54965
rect 9999 54913 10055 54965
rect 10107 54913 10665 54965
rect 9665 54857 10665 54913
rect 9665 54805 9947 54857
rect 9999 54805 10055 54857
rect 10107 54805 10665 54857
rect 9665 54749 10665 54805
rect 9665 54697 9947 54749
rect 9999 54697 10055 54749
rect 10107 54697 10665 54749
rect 9665 54641 10665 54697
rect 9665 54589 9947 54641
rect 9999 54589 10055 54641
rect 10107 54589 10665 54641
rect 9665 54533 10665 54589
rect 9665 54481 9947 54533
rect 9999 54481 10055 54533
rect 10107 54481 10665 54533
rect 9665 54425 10665 54481
rect 9665 54373 9947 54425
rect 9999 54373 10055 54425
rect 10107 54373 10665 54425
rect 9665 54317 10665 54373
rect 9665 54265 9947 54317
rect 9999 54265 10055 54317
rect 10107 54265 10665 54317
rect 9665 54209 10665 54265
rect 9665 54157 9947 54209
rect 9999 54157 10055 54209
rect 10107 54157 10665 54209
rect 9665 54101 10665 54157
rect 9665 54049 9947 54101
rect 9999 54049 10055 54101
rect 10107 54049 10665 54101
rect 9665 53993 10665 54049
rect 9665 53941 9947 53993
rect 9999 53941 10055 53993
rect 10107 53941 10665 53993
rect 9665 53885 10665 53941
rect 9665 53833 9947 53885
rect 9999 53833 10055 53885
rect 10107 53833 10665 53885
rect 9665 53777 10665 53833
rect 9665 53725 9947 53777
rect 9999 53725 10055 53777
rect 10107 53725 10665 53777
rect 9665 53669 10665 53725
rect 9665 53633 9947 53669
rect 7749 53622 9947 53633
rect 9999 53622 10055 53669
rect 10107 53622 10665 53669
rect 7749 53576 7760 53622
rect 10654 53576 10665 53622
rect 7749 53565 10665 53576
rect 10725 56643 11125 56655
rect 10725 56618 10775 56643
rect 10725 53692 10736 56618
rect 10827 56591 10899 56643
rect 10951 56591 11023 56643
rect 11075 56618 11125 56643
rect 10782 56519 11068 56591
rect 10827 56467 10899 56519
rect 10951 56467 11023 56519
rect 10782 56395 11068 56467
rect 10827 56343 10899 56395
rect 10951 56343 11023 56395
rect 10782 56271 11068 56343
rect 10827 56219 10899 56271
rect 10951 56219 11023 56271
rect 10782 56147 11068 56219
rect 10827 56095 10899 56147
rect 10951 56095 11023 56147
rect 10782 56023 11068 56095
rect 10827 55971 10899 56023
rect 10951 55971 11023 56023
rect 10782 55899 11068 55971
rect 10827 55847 10899 55899
rect 10951 55847 11023 55899
rect 10782 55775 11068 55847
rect 10827 55723 10899 55775
rect 10951 55723 11023 55775
rect 10782 55651 11068 55723
rect 10827 55599 10899 55651
rect 10951 55599 11023 55651
rect 10782 55527 11068 55599
rect 10827 55475 10899 55527
rect 10951 55475 11023 55527
rect 10782 55403 11068 55475
rect 10827 55351 10899 55403
rect 10951 55351 11023 55403
rect 10782 55279 11068 55351
rect 10827 55227 10899 55279
rect 10951 55227 11023 55279
rect 10782 55155 11068 55227
rect 10827 55103 10899 55155
rect 10951 55103 11023 55155
rect 10782 55031 11068 55103
rect 10827 54979 10899 55031
rect 10951 54979 11023 55031
rect 10782 54907 11068 54979
rect 10827 54855 10899 54907
rect 10951 54855 11023 54907
rect 10782 54783 11068 54855
rect 10827 54731 10899 54783
rect 10951 54731 11023 54783
rect 10782 54659 11068 54731
rect 10827 54607 10899 54659
rect 10951 54607 11023 54659
rect 10782 54535 11068 54607
rect 10827 54483 10899 54535
rect 10951 54483 11023 54535
rect 10782 54411 11068 54483
rect 10827 54359 10899 54411
rect 10951 54359 11023 54411
rect 10782 54287 11068 54359
rect 10827 54235 10899 54287
rect 10951 54235 11023 54287
rect 10782 54163 11068 54235
rect 10827 54111 10899 54163
rect 10951 54111 11023 54163
rect 10782 54039 11068 54111
rect 10827 53987 10899 54039
rect 10951 53987 11023 54039
rect 10782 53915 11068 53987
rect 10827 53863 10899 53915
rect 10951 53863 11023 53915
rect 10782 53791 11068 53863
rect 10827 53739 10899 53791
rect 10951 53739 11023 53791
rect 10782 53692 11068 53739
rect 11114 53692 11125 56618
rect 10725 53667 11125 53692
rect 10725 53615 10775 53667
rect 10827 53615 10899 53667
rect 10951 53615 11023 53667
rect 11075 53615 11125 53667
rect 10725 53543 11125 53615
rect 11185 53633 12185 56677
rect 13101 53633 14101 56677
rect 14565 56655 14576 57040
rect 11185 53622 14101 53633
rect 11185 53576 11196 53622
rect 14090 53576 14101 53622
rect 11185 53569 12317 53576
rect 12369 53569 12425 53576
rect 12477 53569 14101 53576
rect 11185 53565 14101 53569
rect 14161 56643 14576 56655
rect 14161 56618 14185 56643
rect 14161 53692 14172 56618
rect 14237 56591 14309 56643
rect 14361 56591 14433 56643
rect 14485 56591 14557 56643
rect 14218 56519 14576 56591
rect 14237 56467 14309 56519
rect 14361 56467 14433 56519
rect 14485 56467 14557 56519
rect 14218 56395 14576 56467
rect 14237 56343 14309 56395
rect 14361 56343 14433 56395
rect 14485 56343 14557 56395
rect 14218 56271 14576 56343
rect 14237 56219 14309 56271
rect 14361 56219 14433 56271
rect 14485 56219 14557 56271
rect 14218 56147 14576 56219
rect 14237 56095 14309 56147
rect 14361 56095 14433 56147
rect 14485 56095 14557 56147
rect 14218 56023 14576 56095
rect 14237 55971 14309 56023
rect 14361 55971 14433 56023
rect 14485 55971 14557 56023
rect 14218 55899 14576 55971
rect 14237 55847 14309 55899
rect 14361 55847 14433 55899
rect 14485 55847 14557 55899
rect 14218 55775 14576 55847
rect 14237 55723 14309 55775
rect 14361 55723 14433 55775
rect 14485 55723 14557 55775
rect 14218 55651 14576 55723
rect 14237 55599 14309 55651
rect 14361 55599 14433 55651
rect 14485 55599 14557 55651
rect 14218 55527 14576 55599
rect 14237 55475 14309 55527
rect 14361 55475 14433 55527
rect 14485 55475 14557 55527
rect 14218 55403 14576 55475
rect 14237 55351 14309 55403
rect 14361 55351 14433 55403
rect 14485 55351 14557 55403
rect 14218 55279 14576 55351
rect 14237 55227 14309 55279
rect 14361 55227 14433 55279
rect 14485 55227 14557 55279
rect 14218 55155 14576 55227
rect 14237 55103 14309 55155
rect 14361 55103 14433 55155
rect 14485 55103 14557 55155
rect 14218 55031 14576 55103
rect 14237 54979 14309 55031
rect 14361 54979 14433 55031
rect 14485 54979 14557 55031
rect 14218 54907 14576 54979
rect 14237 54855 14309 54907
rect 14361 54855 14433 54907
rect 14485 54855 14557 54907
rect 14218 54783 14576 54855
rect 14237 54731 14309 54783
rect 14361 54731 14433 54783
rect 14485 54731 14557 54783
rect 14218 54659 14576 54731
rect 14237 54607 14309 54659
rect 14361 54607 14433 54659
rect 14485 54607 14557 54659
rect 14218 54535 14576 54607
rect 14237 54483 14309 54535
rect 14361 54483 14433 54535
rect 14485 54483 14557 54535
rect 14218 54411 14576 54483
rect 14237 54359 14309 54411
rect 14361 54359 14433 54411
rect 14485 54359 14557 54411
rect 14218 54287 14576 54359
rect 14237 54235 14309 54287
rect 14361 54235 14433 54287
rect 14485 54235 14557 54287
rect 14218 54163 14576 54235
rect 14237 54111 14309 54163
rect 14361 54111 14433 54163
rect 14485 54111 14557 54163
rect 14218 54039 14576 54111
rect 14237 53987 14309 54039
rect 14361 53987 14433 54039
rect 14485 53987 14557 54039
rect 14218 53915 14576 53987
rect 14237 53863 14309 53915
rect 14361 53863 14433 53915
rect 14485 53863 14557 53915
rect 14218 53791 14576 53863
rect 14237 53739 14309 53791
rect 14361 53739 14433 53791
rect 14485 53739 14557 53791
rect 14218 53692 14576 53739
rect 14161 53667 14576 53692
rect 14161 53615 14185 53667
rect 14237 53615 14309 53667
rect 14361 53615 14433 53667
rect 14485 53615 14557 53667
rect 12305 53557 12489 53565
rect 10725 53505 10775 53543
rect 4203 53491 10775 53505
rect 10827 53491 10899 53543
rect 10951 53491 11023 53543
rect 11075 53505 11125 53543
rect 14161 53543 14576 53615
rect 14161 53505 14185 53543
rect 11075 53491 14185 53505
rect 14237 53491 14309 53543
rect 14361 53491 14433 53543
rect 14485 53491 14557 53543
rect 402 53483 14576 53491
rect 402 53431 869 53483
rect 921 53431 977 53483
rect 1029 53431 1085 53483
rect 1137 53431 1193 53483
rect 1245 53431 1301 53483
rect 1353 53431 1409 53483
rect 1461 53431 1517 53483
rect 1569 53431 1625 53483
rect 1677 53431 1733 53483
rect 1785 53431 1841 53483
rect 1893 53431 1949 53483
rect 2001 53431 2057 53483
rect 2109 53431 2763 53483
rect 2815 53431 2871 53483
rect 2923 53431 2979 53483
rect 3031 53431 3087 53483
rect 3139 53431 3195 53483
rect 3247 53431 3303 53483
rect 3355 53431 3411 53483
rect 3463 53431 3519 53483
rect 3571 53431 3627 53483
rect 3679 53431 3735 53483
rect 3787 53431 5138 53483
rect 5190 53431 5246 53483
rect 5298 53431 5354 53483
rect 5406 53431 5462 53483
rect 5514 53431 5570 53483
rect 5622 53431 5678 53483
rect 5730 53431 5786 53483
rect 5838 53431 5894 53483
rect 5946 53431 6002 53483
rect 6054 53431 6110 53483
rect 6162 53431 6218 53483
rect 6270 53431 6326 53483
rect 6378 53431 6434 53483
rect 6486 53431 6542 53483
rect 6594 53431 6650 53483
rect 6702 53431 6758 53483
rect 6810 53431 6866 53483
rect 6918 53431 6974 53483
rect 7026 53431 7082 53483
rect 7134 53431 7844 53483
rect 7896 53431 7952 53483
rect 8004 53431 8060 53483
rect 8112 53431 8168 53483
rect 8220 53431 8276 53483
rect 8328 53431 8384 53483
rect 8436 53431 8492 53483
rect 8544 53431 8600 53483
rect 8652 53431 8708 53483
rect 8760 53431 8816 53483
rect 8868 53431 8924 53483
rect 8976 53431 9032 53483
rect 9084 53431 9140 53483
rect 9192 53431 9248 53483
rect 9300 53431 9356 53483
rect 9408 53431 9464 53483
rect 9516 53431 9572 53483
rect 9624 53431 9680 53483
rect 9732 53431 9788 53483
rect 9840 53431 11191 53483
rect 11243 53431 11299 53483
rect 11351 53431 11407 53483
rect 11459 53431 11515 53483
rect 11567 53431 11623 53483
rect 11675 53431 11731 53483
rect 11783 53431 11839 53483
rect 11891 53431 11947 53483
rect 11999 53431 12055 53483
rect 12107 53431 12163 53483
rect 12215 53431 12869 53483
rect 12921 53431 12977 53483
rect 13029 53431 13085 53483
rect 13137 53431 13193 53483
rect 13245 53431 13301 53483
rect 13353 53431 13409 53483
rect 13461 53431 13517 53483
rect 13569 53431 13625 53483
rect 13677 53431 13733 53483
rect 13785 53431 13841 53483
rect 13893 53431 13949 53483
rect 14001 53431 14057 53483
rect 14109 53431 14576 53483
rect 402 53419 14576 53431
rect 421 53367 493 53419
rect 545 53367 617 53419
rect 669 53367 741 53419
rect 793 53375 3903 53419
rect 793 53367 869 53375
rect 402 53323 869 53367
rect 921 53323 977 53375
rect 1029 53323 1085 53375
rect 1137 53323 1193 53375
rect 1245 53323 1301 53375
rect 1353 53323 1409 53375
rect 1461 53323 1517 53375
rect 1569 53323 1625 53375
rect 1677 53323 1733 53375
rect 1785 53323 1841 53375
rect 1893 53323 1949 53375
rect 2001 53323 2057 53375
rect 2109 53323 2763 53375
rect 2815 53323 2871 53375
rect 2923 53323 2979 53375
rect 3031 53323 3087 53375
rect 3139 53323 3195 53375
rect 3247 53323 3303 53375
rect 3355 53323 3411 53375
rect 3463 53323 3519 53375
rect 3571 53323 3627 53375
rect 3679 53323 3735 53375
rect 3787 53367 3903 53375
rect 3955 53367 4027 53419
rect 4079 53367 4151 53419
rect 4203 53375 10775 53419
rect 4203 53367 5138 53375
rect 3787 53323 5138 53367
rect 5190 53323 5246 53375
rect 5298 53323 5354 53375
rect 5406 53323 5462 53375
rect 5514 53323 5570 53375
rect 5622 53323 5678 53375
rect 5730 53323 5786 53375
rect 5838 53323 5894 53375
rect 5946 53323 6002 53375
rect 6054 53323 6110 53375
rect 6162 53323 6218 53375
rect 6270 53323 6326 53375
rect 6378 53323 6434 53375
rect 6486 53323 6542 53375
rect 6594 53323 6650 53375
rect 6702 53323 6758 53375
rect 6810 53323 6866 53375
rect 6918 53323 6974 53375
rect 7026 53323 7082 53375
rect 7134 53323 7844 53375
rect 7896 53323 7952 53375
rect 8004 53323 8060 53375
rect 8112 53323 8168 53375
rect 8220 53323 8276 53375
rect 8328 53323 8384 53375
rect 8436 53323 8492 53375
rect 8544 53323 8600 53375
rect 8652 53323 8708 53375
rect 8760 53323 8816 53375
rect 8868 53323 8924 53375
rect 8976 53323 9032 53375
rect 9084 53323 9140 53375
rect 9192 53323 9248 53375
rect 9300 53323 9356 53375
rect 9408 53323 9464 53375
rect 9516 53323 9572 53375
rect 9624 53323 9680 53375
rect 9732 53323 9788 53375
rect 9840 53367 10775 53375
rect 10827 53367 10899 53419
rect 10951 53367 11023 53419
rect 11075 53375 14185 53419
rect 11075 53367 11191 53375
rect 9840 53323 11191 53367
rect 11243 53323 11299 53375
rect 11351 53323 11407 53375
rect 11459 53323 11515 53375
rect 11567 53323 11623 53375
rect 11675 53323 11731 53375
rect 11783 53323 11839 53375
rect 11891 53323 11947 53375
rect 11999 53323 12055 53375
rect 12107 53323 12163 53375
rect 12215 53323 12869 53375
rect 12921 53323 12977 53375
rect 13029 53323 13085 53375
rect 13137 53323 13193 53375
rect 13245 53323 13301 53375
rect 13353 53323 13409 53375
rect 13461 53323 13517 53375
rect 13569 53323 13625 53375
rect 13677 53323 13733 53375
rect 13785 53323 13841 53375
rect 13893 53323 13949 53375
rect 14001 53323 14057 53375
rect 14109 53367 14185 53375
rect 14237 53367 14309 53419
rect 14361 53367 14433 53419
rect 14485 53367 14557 53419
rect 14109 53323 14576 53367
rect 402 53295 14576 53323
rect 421 53243 493 53295
rect 545 53251 617 53295
rect 669 53251 741 53295
rect 793 53267 3903 53295
rect 793 53251 869 53267
rect 921 53251 977 53267
rect 1029 53251 1085 53267
rect 1137 53251 1193 53267
rect 1245 53251 1301 53267
rect 1353 53251 1409 53267
rect 1461 53251 1517 53267
rect 1569 53251 1625 53267
rect 1677 53251 1733 53267
rect 1785 53251 1841 53267
rect 1893 53251 1949 53267
rect 2001 53251 2057 53267
rect 2109 53251 2763 53267
rect 2815 53251 2871 53267
rect 2923 53251 2979 53267
rect 3031 53251 3087 53267
rect 3139 53251 3195 53267
rect 3247 53251 3303 53267
rect 3355 53251 3411 53267
rect 3463 53251 3519 53267
rect 3571 53251 3627 53267
rect 3679 53251 3735 53267
rect 3787 53251 3903 53267
rect 3955 53251 4027 53295
rect 4079 53251 4151 53295
rect 4203 53267 10775 53295
rect 4203 53251 5138 53267
rect 5190 53251 5246 53267
rect 5298 53251 5354 53267
rect 5406 53251 5462 53267
rect 5514 53251 5570 53267
rect 5622 53251 5678 53267
rect 5730 53251 5786 53267
rect 5838 53251 5894 53267
rect 5946 53251 6002 53267
rect 6054 53251 6110 53267
rect 6162 53251 6218 53267
rect 6270 53251 6326 53267
rect 6378 53251 6434 53267
rect 6486 53251 6542 53267
rect 6594 53251 6650 53267
rect 6702 53251 6758 53267
rect 6810 53251 6866 53267
rect 6918 53251 6974 53267
rect 7026 53251 7082 53267
rect 7134 53251 7844 53267
rect 7896 53251 7952 53267
rect 8004 53251 8060 53267
rect 8112 53251 8168 53267
rect 8220 53251 8276 53267
rect 8328 53251 8384 53267
rect 8436 53251 8492 53267
rect 8544 53251 8600 53267
rect 8652 53251 8708 53267
rect 8760 53251 8816 53267
rect 8868 53251 8924 53267
rect 8976 53251 9032 53267
rect 9084 53251 9140 53267
rect 9192 53251 9248 53267
rect 9300 53251 9356 53267
rect 9408 53251 9464 53267
rect 9516 53251 9572 53267
rect 9624 53251 9680 53267
rect 9732 53251 9788 53267
rect 9840 53251 10775 53267
rect 10827 53251 10899 53295
rect 10951 53251 11023 53295
rect 11075 53267 14185 53295
rect 11075 53251 11191 53267
rect 11243 53251 11299 53267
rect 11351 53251 11407 53267
rect 11459 53251 11515 53267
rect 11567 53251 11623 53267
rect 11675 53251 11731 53267
rect 11783 53251 11839 53267
rect 11891 53251 11947 53267
rect 11999 53251 12055 53267
rect 12107 53251 12163 53267
rect 12215 53251 12869 53267
rect 12921 53251 12977 53267
rect 13029 53251 13085 53267
rect 13137 53251 13193 53267
rect 13245 53251 13301 53267
rect 13353 53251 13409 53267
rect 13461 53251 13517 53267
rect 13569 53251 13625 53267
rect 13677 53251 13733 53267
rect 13785 53251 13841 53267
rect 13893 53251 13949 53267
rect 14001 53251 14057 53267
rect 14109 53251 14185 53267
rect 14237 53251 14309 53295
rect 14361 53251 14433 53295
rect 402 53205 510 53243
rect 14485 53243 14557 53295
rect 14468 53205 14576 53243
rect 14622 53205 14633 57105
rect 14892 57099 14904 57151
rect 14956 57099 14968 57151
rect 14892 57043 14968 57099
rect 14892 56991 14904 57043
rect 14956 56991 14968 57043
rect 14892 56935 14968 56991
rect 14892 56883 14904 56935
rect 14956 56883 14968 56935
rect 14892 56827 14968 56883
rect 14892 56775 14904 56827
rect 14956 56775 14968 56827
rect 14892 56719 14968 56775
rect 14892 56667 14904 56719
rect 14956 56667 14968 56719
rect 14892 56611 14968 56667
rect 14892 56559 14904 56611
rect 14956 56559 14968 56611
rect 14892 56503 14968 56559
rect 14892 56451 14904 56503
rect 14956 56451 14968 56503
rect 14892 56395 14968 56451
rect 14892 56343 14904 56395
rect 14956 56343 14968 56395
rect 14892 56287 14968 56343
rect 14892 56235 14904 56287
rect 14956 56235 14968 56287
rect 14892 56179 14968 56235
rect 14892 56127 14904 56179
rect 14956 56127 14968 56179
rect 14892 56071 14968 56127
rect 14892 56019 14904 56071
rect 14956 56019 14968 56071
rect 14892 56007 14968 56019
rect 345 53194 14633 53205
rect 14892 54174 14968 54186
rect 14892 54122 14904 54174
rect 14956 54122 14968 54174
rect 14892 54066 14968 54122
rect 14892 54014 14904 54066
rect 14956 54014 14968 54066
rect 14892 53958 14968 54014
rect 14892 53906 14904 53958
rect 14956 53906 14968 53958
rect 14892 53850 14968 53906
rect 14892 53798 14904 53850
rect 14956 53798 14968 53850
rect 14892 53742 14968 53798
rect 14892 53690 14904 53742
rect 14956 53690 14968 53742
rect 14892 53634 14968 53690
rect 14892 53582 14904 53634
rect 14956 53582 14968 53634
rect 14892 53526 14968 53582
rect 14892 53474 14904 53526
rect 14956 53474 14968 53526
rect 14892 53418 14968 53474
rect 14892 53366 14904 53418
rect 14956 53366 14968 53418
rect 14892 53310 14968 53366
rect 14892 53258 14904 53310
rect 14956 53258 14968 53310
rect 14892 53202 14968 53258
rect 10 53094 86 53150
rect 10 53042 22 53094
rect 74 53042 86 53094
rect 10 52986 86 53042
rect 10 52934 22 52986
rect 74 52934 86 52986
rect 10 52878 86 52934
rect 10 52826 22 52878
rect 74 52826 86 52878
rect 10 52814 86 52826
rect 14892 53150 14904 53202
rect 14956 53150 14968 53202
rect 14892 53094 14968 53150
rect 14892 53042 14904 53094
rect 14956 53042 14968 53094
rect 14892 52986 14968 53042
rect 14892 52934 14904 52986
rect 14956 52934 14968 52986
rect 14892 52878 14968 52934
rect 14892 52826 14904 52878
rect 14956 52826 14968 52878
rect 14892 52814 14968 52826
rect 71 52611 2225 52622
rect 71 52586 268 52611
rect 10 52574 268 52586
rect 10 52522 22 52574
rect 74 52522 268 52574
rect 10 52466 268 52522
rect 10 52414 22 52466
rect 74 52414 268 52466
rect 10 52358 268 52414
rect 10 52306 22 52358
rect 74 52306 268 52358
rect 10 52250 268 52306
rect 10 52198 22 52250
rect 74 52198 268 52250
rect 10 52142 268 52198
rect 10 52090 22 52142
rect 74 52090 268 52142
rect 10 52034 268 52090
rect 10 51982 22 52034
rect 74 51982 268 52034
rect 10 51926 268 51982
rect 10 51874 22 51926
rect 74 51874 268 51926
rect 10 51818 268 51874
rect 10 51766 22 51818
rect 74 51766 268 51818
rect 10 51710 268 51766
rect 10 51658 22 51710
rect 74 51658 268 51710
rect 10 51622 268 51658
rect 10 51602 86 51622
rect 10 51550 22 51602
rect 74 51550 86 51602
rect 10 51494 86 51550
rect 10 51442 22 51494
rect 74 51442 86 51494
rect 10 51422 86 51442
rect 257 51422 268 51622
rect 10 51386 268 51422
rect 10 51334 22 51386
rect 74 51334 268 51386
rect 10 51278 268 51334
rect 10 51226 22 51278
rect 74 51226 268 51278
rect 10 51214 268 51226
rect 71 50422 268 51214
rect 257 49854 268 50422
rect 71 49386 268 49854
rect 10 49374 268 49386
rect 10 49322 22 49374
rect 74 49322 268 49374
rect 10 49266 268 49322
rect 10 49214 22 49266
rect 74 49214 268 49266
rect 10 49158 268 49214
rect 10 49106 22 49158
rect 74 49106 268 49158
rect 10 49050 268 49106
rect 10 48998 22 49050
rect 74 48998 268 49050
rect 10 48942 268 48998
rect 10 48890 22 48942
rect 74 48890 268 48942
rect 10 48854 268 48890
rect 10 48834 86 48854
rect 10 48782 22 48834
rect 74 48782 86 48834
rect 10 48726 86 48782
rect 10 48674 22 48726
rect 74 48674 86 48726
rect 10 48654 86 48674
rect 257 48654 268 48854
rect 10 48618 268 48654
rect 10 48566 22 48618
rect 74 48566 268 48618
rect 10 48510 268 48566
rect 10 48458 22 48510
rect 74 48458 268 48510
rect 10 48402 268 48458
rect 10 48350 22 48402
rect 74 48350 268 48402
rect 10 48294 268 48350
rect 10 48242 22 48294
rect 74 48242 268 48294
rect 10 48186 268 48242
rect 10 48134 22 48186
rect 74 48134 268 48186
rect 10 48078 268 48134
rect 10 48026 22 48078
rect 74 48026 268 48078
rect 10 48014 268 48026
rect 71 47665 268 48014
rect 2214 47665 2225 52611
rect 71 47654 2225 47665
rect 2551 52611 12427 52622
rect 2551 47665 2562 52611
rect 2908 52265 3016 52611
rect 11962 52265 12070 52611
rect 2908 52254 12070 52265
rect 2908 48022 2919 52254
rect 3105 52029 11873 52040
rect 3105 51983 3142 52029
rect 11836 51983 11873 52029
rect 3105 51957 3161 51983
rect 3213 51957 3269 51983
rect 3321 51957 3377 51983
rect 3429 51957 3485 51983
rect 3537 51957 3593 51983
rect 3645 51957 3701 51983
rect 3753 51957 3809 51983
rect 3861 51957 3917 51983
rect 3969 51957 4025 51983
rect 4077 51957 4133 51983
rect 4185 51957 4241 51983
rect 4293 51957 4349 51983
rect 4401 51957 4457 51983
rect 4509 51957 4565 51983
rect 4617 51957 4673 51983
rect 4725 51957 5138 51983
rect 5190 51957 5246 51983
rect 5298 51957 5354 51983
rect 5406 51957 5462 51983
rect 5514 51957 5570 51983
rect 5622 51957 5678 51983
rect 5730 51957 5786 51983
rect 5838 51957 5894 51983
rect 5946 51957 6002 51983
rect 6054 51957 6110 51983
rect 6162 51957 6218 51983
rect 6270 51957 6326 51983
rect 6378 51957 6434 51983
rect 6486 51957 6542 51983
rect 6594 51957 6650 51983
rect 6702 51957 6758 51983
rect 6810 51957 6866 51983
rect 6918 51957 6974 51983
rect 7026 51957 7082 51983
rect 7134 51957 7844 51983
rect 7896 51957 7952 51983
rect 8004 51957 8060 51983
rect 8112 51957 8168 51983
rect 8220 51957 8276 51983
rect 8328 51957 8384 51983
rect 8436 51957 8492 51983
rect 8544 51957 8600 51983
rect 8652 51957 8708 51983
rect 8760 51957 8816 51983
rect 8868 51957 8924 51983
rect 8976 51957 9032 51983
rect 9084 51957 9140 51983
rect 9192 51957 9248 51983
rect 9300 51957 9356 51983
rect 9408 51957 9464 51983
rect 9516 51957 9572 51983
rect 9624 51957 9680 51983
rect 9732 51957 9788 51983
rect 9840 51957 10253 51983
rect 10305 51957 10361 51983
rect 10413 51957 10469 51983
rect 10521 51957 10577 51983
rect 10629 51957 10685 51983
rect 10737 51957 10793 51983
rect 10845 51957 10901 51983
rect 10953 51957 11009 51983
rect 11061 51957 11117 51983
rect 11169 51957 11225 51983
rect 11277 51957 11333 51983
rect 11385 51957 11441 51983
rect 11493 51957 11549 51983
rect 11601 51957 11657 51983
rect 11709 51957 11765 51983
rect 11817 51957 11873 51983
rect 3105 51901 11873 51957
rect 3105 51900 3161 51901
rect 3105 48376 3116 51900
rect 3213 51849 3269 51901
rect 3321 51849 3377 51901
rect 3429 51875 3485 51901
rect 3537 51875 3593 51901
rect 3645 51875 3701 51901
rect 3753 51875 3809 51901
rect 3861 51875 3917 51901
rect 3969 51875 4025 51901
rect 4077 51875 4133 51901
rect 4185 51875 4241 51901
rect 4293 51875 4349 51901
rect 4401 51875 4457 51901
rect 4509 51875 4565 51901
rect 4617 51875 4673 51901
rect 4725 51875 5138 51901
rect 5190 51875 5246 51901
rect 5298 51875 5354 51901
rect 5406 51875 5462 51901
rect 5514 51875 5570 51901
rect 5622 51875 5678 51901
rect 5730 51875 5786 51901
rect 5838 51875 5894 51901
rect 5946 51875 6002 51901
rect 6054 51875 6110 51901
rect 6162 51875 6218 51901
rect 6270 51875 6326 51901
rect 6378 51875 6434 51901
rect 6486 51875 6542 51901
rect 6594 51875 6650 51901
rect 6702 51875 6758 51901
rect 6810 51875 6866 51901
rect 6918 51875 6974 51901
rect 7026 51875 7082 51901
rect 7134 51875 7844 51901
rect 7896 51875 7952 51901
rect 8004 51875 8060 51901
rect 8112 51875 8168 51901
rect 8220 51875 8276 51901
rect 8328 51875 8384 51901
rect 8436 51875 8492 51901
rect 8544 51875 8600 51901
rect 8652 51875 8708 51901
rect 8760 51875 8816 51901
rect 8868 51875 8924 51901
rect 8976 51875 9032 51901
rect 9084 51875 9140 51901
rect 9192 51875 9248 51901
rect 9300 51875 9356 51901
rect 9408 51875 9464 51901
rect 9516 51875 9572 51901
rect 9624 51875 9680 51901
rect 9732 51875 9788 51901
rect 9840 51875 10253 51901
rect 10305 51875 10361 51901
rect 10413 51875 10469 51901
rect 10521 51875 10577 51901
rect 10629 51875 10685 51901
rect 10737 51875 10793 51901
rect 10845 51875 10901 51901
rect 10953 51875 11009 51901
rect 11061 51875 11117 51901
rect 11169 51875 11225 51901
rect 11277 51875 11333 51901
rect 11385 51875 11441 51901
rect 11493 51875 11549 51901
rect 11601 51849 11657 51901
rect 11709 51849 11765 51901
rect 11817 51900 11873 51901
rect 3162 51844 3424 51849
rect 3162 51234 3270 51844
rect 3316 51829 3424 51844
rect 11554 51844 11816 51849
rect 11554 51829 11662 51844
rect 3316 51818 11662 51829
rect 3316 51260 3327 51818
rect 3489 51626 11489 51639
rect 3489 51580 3502 51626
rect 11476 51580 11489 51626
rect 3489 51567 4871 51580
rect 4923 51567 4979 51580
rect 5031 51567 7247 51580
rect 7299 51567 7355 51580
rect 7407 51567 7463 51580
rect 7515 51567 7571 51580
rect 7623 51567 7679 51580
rect 7731 51567 9947 51580
rect 9999 51567 10055 51580
rect 10107 51567 11489 51580
rect 3489 51511 11489 51567
rect 3489 51498 4871 51511
rect 4923 51498 4979 51511
rect 5031 51498 7247 51511
rect 7299 51498 7355 51511
rect 7407 51498 7463 51511
rect 7515 51498 7571 51511
rect 7623 51498 7679 51511
rect 7731 51498 9947 51511
rect 9999 51498 10055 51511
rect 10107 51498 11489 51511
rect 3489 51452 3502 51498
rect 11476 51452 11489 51498
rect 3489 51439 11489 51452
rect 11651 51260 11662 51818
rect 3316 51249 11662 51260
rect 3316 51234 3424 51249
rect 3162 51206 3424 51234
rect 11554 51234 11662 51249
rect 11708 51234 11816 51844
rect 11554 51206 11816 51234
rect 3213 51154 3269 51206
rect 3321 51154 3377 51206
rect 3429 51154 3485 51203
rect 3537 51154 3593 51203
rect 3645 51154 3701 51203
rect 3753 51154 3809 51203
rect 3861 51154 3917 51203
rect 3969 51154 4025 51203
rect 4077 51154 4133 51203
rect 4185 51154 4241 51203
rect 4293 51154 4349 51203
rect 4401 51154 4457 51203
rect 4509 51154 4565 51203
rect 4617 51154 4673 51203
rect 4725 51154 5138 51203
rect 5190 51154 5246 51203
rect 5298 51154 5354 51203
rect 5406 51154 5462 51203
rect 5514 51154 5570 51203
rect 5622 51154 5678 51203
rect 5730 51154 5786 51203
rect 5838 51154 5894 51203
rect 5946 51154 6002 51203
rect 6054 51154 6110 51203
rect 6162 51154 6218 51203
rect 6270 51154 6326 51203
rect 6378 51154 6434 51203
rect 6486 51154 6542 51203
rect 6594 51154 6650 51203
rect 6702 51154 6758 51203
rect 6810 51154 6866 51203
rect 6918 51154 6974 51203
rect 7026 51154 7082 51203
rect 7134 51154 7844 51203
rect 7896 51154 7952 51203
rect 8004 51154 8060 51203
rect 8112 51154 8168 51203
rect 8220 51154 8276 51203
rect 8328 51154 8384 51203
rect 8436 51154 8492 51203
rect 8544 51154 8600 51203
rect 8652 51154 8708 51203
rect 8760 51154 8816 51203
rect 8868 51154 8924 51203
rect 8976 51154 9032 51203
rect 9084 51154 9140 51203
rect 9192 51154 9248 51203
rect 9300 51154 9356 51203
rect 9408 51154 9464 51203
rect 9516 51154 9572 51203
rect 9624 51154 9680 51203
rect 9732 51154 9788 51203
rect 9840 51154 10253 51203
rect 10305 51154 10361 51203
rect 10413 51154 10469 51203
rect 10521 51154 10577 51203
rect 10629 51154 10685 51203
rect 10737 51154 10793 51203
rect 10845 51154 10901 51203
rect 10953 51154 11009 51203
rect 11061 51154 11117 51203
rect 11169 51154 11225 51203
rect 11277 51154 11333 51203
rect 11385 51154 11441 51203
rect 11493 51154 11549 51203
rect 11601 51154 11657 51206
rect 11709 51154 11765 51206
rect 3162 51098 11816 51154
rect 3213 51046 3269 51098
rect 3321 51095 3377 51098
rect 3429 51095 3485 51098
rect 3537 51095 3593 51098
rect 3645 51095 3701 51098
rect 3753 51095 3809 51098
rect 3861 51095 3917 51098
rect 3969 51095 4025 51098
rect 4077 51095 4133 51098
rect 4185 51095 4241 51098
rect 4293 51095 4349 51098
rect 4401 51095 4457 51098
rect 4509 51095 4565 51098
rect 4617 51095 4673 51098
rect 4725 51095 5138 51098
rect 5190 51095 5246 51098
rect 5298 51095 5354 51098
rect 5406 51095 5462 51098
rect 5514 51095 5570 51098
rect 5622 51095 5678 51098
rect 5730 51095 5786 51098
rect 5838 51095 5894 51098
rect 5946 51095 6002 51098
rect 6054 51095 6110 51098
rect 6162 51095 6218 51098
rect 6270 51095 6326 51098
rect 6378 51095 6434 51098
rect 6486 51095 6542 51098
rect 6594 51095 6650 51098
rect 6702 51095 6758 51098
rect 6810 51095 6866 51098
rect 6918 51095 6974 51098
rect 7026 51095 7082 51098
rect 7134 51095 7844 51098
rect 7896 51095 7952 51098
rect 8004 51095 8060 51098
rect 8112 51095 8168 51098
rect 8220 51095 8276 51098
rect 8328 51095 8384 51098
rect 8436 51095 8492 51098
rect 8544 51095 8600 51098
rect 8652 51095 8708 51098
rect 8760 51095 8816 51098
rect 8868 51095 8924 51098
rect 8976 51095 9032 51098
rect 9084 51095 9140 51098
rect 9192 51095 9248 51098
rect 9300 51095 9356 51098
rect 9408 51095 9464 51098
rect 9516 51095 9572 51098
rect 9624 51095 9680 51098
rect 9732 51095 9788 51098
rect 9840 51095 10253 51098
rect 10305 51095 10361 51098
rect 10413 51095 10469 51098
rect 10521 51095 10577 51098
rect 10629 51095 10685 51098
rect 10737 51095 10793 51098
rect 10845 51095 10901 51098
rect 10953 51095 11009 51098
rect 11061 51095 11117 51098
rect 11169 51095 11225 51098
rect 11277 51095 11333 51098
rect 11385 51095 11441 51098
rect 11493 51095 11549 51098
rect 11601 51095 11657 51098
rect 3321 51049 3330 51095
rect 11648 51049 11657 51095
rect 3321 51046 3377 51049
rect 3429 51046 3485 51049
rect 3537 51046 3593 51049
rect 3645 51046 3701 51049
rect 3753 51046 3809 51049
rect 3861 51046 3917 51049
rect 3969 51046 4025 51049
rect 4077 51046 4133 51049
rect 4185 51046 4241 51049
rect 4293 51046 4349 51049
rect 4401 51046 4457 51049
rect 4509 51046 4565 51049
rect 4617 51046 4673 51049
rect 4725 51046 5138 51049
rect 5190 51046 5246 51049
rect 5298 51046 5354 51049
rect 5406 51046 5462 51049
rect 5514 51046 5570 51049
rect 5622 51046 5678 51049
rect 5730 51046 5786 51049
rect 5838 51046 5894 51049
rect 5946 51046 6002 51049
rect 6054 51046 6110 51049
rect 6162 51046 6218 51049
rect 6270 51046 6326 51049
rect 6378 51046 6434 51049
rect 6486 51046 6542 51049
rect 6594 51046 6650 51049
rect 6702 51046 6758 51049
rect 6810 51046 6866 51049
rect 6918 51046 6974 51049
rect 7026 51046 7082 51049
rect 7134 51046 7844 51049
rect 7896 51046 7952 51049
rect 8004 51046 8060 51049
rect 8112 51046 8168 51049
rect 8220 51046 8276 51049
rect 8328 51046 8384 51049
rect 8436 51046 8492 51049
rect 8544 51046 8600 51049
rect 8652 51046 8708 51049
rect 8760 51046 8816 51049
rect 8868 51046 8924 51049
rect 8976 51046 9032 51049
rect 9084 51046 9140 51049
rect 9192 51046 9248 51049
rect 9300 51046 9356 51049
rect 9408 51046 9464 51049
rect 9516 51046 9572 51049
rect 9624 51046 9680 51049
rect 9732 51046 9788 51049
rect 9840 51046 10253 51049
rect 10305 51046 10361 51049
rect 10413 51046 10469 51049
rect 10521 51046 10577 51049
rect 10629 51046 10685 51049
rect 10737 51046 10793 51049
rect 10845 51046 10901 51049
rect 10953 51046 11009 51049
rect 11061 51046 11117 51049
rect 11169 51046 11225 51049
rect 11277 51046 11333 51049
rect 11385 51046 11441 51049
rect 11493 51046 11549 51049
rect 11601 51046 11657 51049
rect 11709 51046 11765 51098
rect 3162 50990 11816 51046
rect 3213 50938 3269 50990
rect 3321 50938 3377 50990
rect 3429 50941 3485 50990
rect 3537 50941 3593 50990
rect 3645 50941 3701 50990
rect 3753 50941 3809 50990
rect 3861 50941 3917 50990
rect 3969 50941 4025 50990
rect 4077 50941 4133 50990
rect 4185 50941 4241 50990
rect 4293 50941 4349 50990
rect 4401 50941 4457 50990
rect 4509 50941 4565 50990
rect 4617 50941 4673 50990
rect 4725 50941 5138 50990
rect 5190 50941 5246 50990
rect 5298 50941 5354 50990
rect 5406 50941 5462 50990
rect 5514 50941 5570 50990
rect 5622 50941 5678 50990
rect 5730 50941 5786 50990
rect 5838 50941 5894 50990
rect 5946 50941 6002 50990
rect 6054 50941 6110 50990
rect 6162 50941 6218 50990
rect 6270 50941 6326 50990
rect 6378 50941 6434 50990
rect 6486 50941 6542 50990
rect 6594 50941 6650 50990
rect 6702 50941 6758 50990
rect 6810 50941 6866 50990
rect 6918 50941 6974 50990
rect 7026 50941 7082 50990
rect 7134 50941 7844 50990
rect 7896 50941 7952 50990
rect 8004 50941 8060 50990
rect 8112 50941 8168 50990
rect 8220 50941 8276 50990
rect 8328 50941 8384 50990
rect 8436 50941 8492 50990
rect 8544 50941 8600 50990
rect 8652 50941 8708 50990
rect 8760 50941 8816 50990
rect 8868 50941 8924 50990
rect 8976 50941 9032 50990
rect 9084 50941 9140 50990
rect 9192 50941 9248 50990
rect 9300 50941 9356 50990
rect 9408 50941 9464 50990
rect 9516 50941 9572 50990
rect 9624 50941 9680 50990
rect 9732 50941 9788 50990
rect 9840 50941 10253 50990
rect 10305 50941 10361 50990
rect 10413 50941 10469 50990
rect 10521 50941 10577 50990
rect 10629 50941 10685 50990
rect 10737 50941 10793 50990
rect 10845 50941 10901 50990
rect 10953 50941 11009 50990
rect 11061 50941 11117 50990
rect 11169 50941 11225 50990
rect 11277 50941 11333 50990
rect 11385 50941 11441 50990
rect 11493 50941 11549 50990
rect 11601 50938 11657 50990
rect 11709 50938 11765 50990
rect 3162 50910 3424 50938
rect 3162 50300 3270 50910
rect 3316 50895 3424 50910
rect 11554 50910 11816 50938
rect 11554 50895 11662 50910
rect 3316 50884 11662 50895
rect 3316 50326 3327 50884
rect 3489 50692 11489 50705
rect 3489 50646 3502 50692
rect 11476 50646 11489 50692
rect 3489 50633 4871 50646
rect 4923 50633 4979 50646
rect 5031 50633 7247 50646
rect 7299 50633 7355 50646
rect 7407 50633 7463 50646
rect 7515 50633 7571 50646
rect 7623 50633 7679 50646
rect 7731 50633 9947 50646
rect 9999 50633 10055 50646
rect 10107 50633 11489 50646
rect 3489 50577 11489 50633
rect 3489 50564 4871 50577
rect 4923 50564 4979 50577
rect 5031 50564 7247 50577
rect 7299 50564 7355 50577
rect 7407 50564 7463 50577
rect 7515 50564 7571 50577
rect 7623 50564 7679 50577
rect 7731 50564 9947 50577
rect 9999 50564 10055 50577
rect 10107 50564 11489 50577
rect 3489 50518 3502 50564
rect 11476 50518 11489 50564
rect 3489 50505 11489 50518
rect 11651 50326 11662 50884
rect 3316 50315 11662 50326
rect 3316 50300 3424 50315
rect 3162 50272 3424 50300
rect 11554 50300 11662 50315
rect 11708 50300 11816 50910
rect 11554 50272 11816 50300
rect 3213 50220 3269 50272
rect 3321 50220 3377 50272
rect 3429 50220 3485 50269
rect 3537 50220 3593 50269
rect 3645 50220 3701 50269
rect 3753 50220 3809 50269
rect 3861 50220 3917 50269
rect 3969 50220 4025 50269
rect 4077 50220 4133 50269
rect 4185 50220 4241 50269
rect 4293 50220 4349 50269
rect 4401 50220 4457 50269
rect 4509 50220 4565 50269
rect 4617 50220 4673 50269
rect 4725 50220 5138 50269
rect 5190 50220 5246 50269
rect 5298 50220 5354 50269
rect 5406 50220 5462 50269
rect 5514 50220 5570 50269
rect 5622 50220 5678 50269
rect 5730 50220 5786 50269
rect 5838 50220 5894 50269
rect 5946 50220 6002 50269
rect 6054 50220 6110 50269
rect 6162 50220 6218 50269
rect 6270 50220 6326 50269
rect 6378 50220 6434 50269
rect 6486 50220 6542 50269
rect 6594 50220 6650 50269
rect 6702 50220 6758 50269
rect 6810 50220 6866 50269
rect 6918 50220 6974 50269
rect 7026 50220 7082 50269
rect 7134 50220 7844 50269
rect 7896 50220 7952 50269
rect 8004 50220 8060 50269
rect 8112 50220 8168 50269
rect 8220 50220 8276 50269
rect 8328 50220 8384 50269
rect 8436 50220 8492 50269
rect 8544 50220 8600 50269
rect 8652 50220 8708 50269
rect 8760 50220 8816 50269
rect 8868 50220 8924 50269
rect 8976 50220 9032 50269
rect 9084 50220 9140 50269
rect 9192 50220 9248 50269
rect 9300 50220 9356 50269
rect 9408 50220 9464 50269
rect 9516 50220 9572 50269
rect 9624 50220 9680 50269
rect 9732 50220 9788 50269
rect 9840 50220 10253 50269
rect 10305 50220 10361 50269
rect 10413 50220 10469 50269
rect 10521 50220 10577 50269
rect 10629 50220 10685 50269
rect 10737 50220 10793 50269
rect 10845 50220 10901 50269
rect 10953 50220 11009 50269
rect 11061 50220 11117 50269
rect 11169 50220 11225 50269
rect 11277 50220 11333 50269
rect 11385 50220 11441 50269
rect 11493 50220 11549 50269
rect 11601 50220 11657 50272
rect 11709 50220 11765 50272
rect 3162 50164 11816 50220
rect 3213 50112 3269 50164
rect 3321 50161 3377 50164
rect 3429 50161 3485 50164
rect 3537 50161 3593 50164
rect 3645 50161 3701 50164
rect 3753 50161 3809 50164
rect 3861 50161 3917 50164
rect 3969 50161 4025 50164
rect 4077 50161 4133 50164
rect 4185 50161 4241 50164
rect 4293 50161 4349 50164
rect 4401 50161 4457 50164
rect 4509 50161 4565 50164
rect 4617 50161 4673 50164
rect 4725 50161 5138 50164
rect 5190 50161 5246 50164
rect 5298 50161 5354 50164
rect 5406 50161 5462 50164
rect 5514 50161 5570 50164
rect 5622 50161 5678 50164
rect 5730 50161 5786 50164
rect 5838 50161 5894 50164
rect 5946 50161 6002 50164
rect 6054 50161 6110 50164
rect 6162 50161 6218 50164
rect 6270 50161 6326 50164
rect 6378 50161 6434 50164
rect 6486 50161 6542 50164
rect 6594 50161 6650 50164
rect 6702 50161 6758 50164
rect 6810 50161 6866 50164
rect 6918 50161 6974 50164
rect 7026 50161 7082 50164
rect 7134 50161 7844 50164
rect 7896 50161 7952 50164
rect 8004 50161 8060 50164
rect 8112 50161 8168 50164
rect 8220 50161 8276 50164
rect 8328 50161 8384 50164
rect 8436 50161 8492 50164
rect 8544 50161 8600 50164
rect 8652 50161 8708 50164
rect 8760 50161 8816 50164
rect 8868 50161 8924 50164
rect 8976 50161 9032 50164
rect 9084 50161 9140 50164
rect 9192 50161 9248 50164
rect 9300 50161 9356 50164
rect 9408 50161 9464 50164
rect 9516 50161 9572 50164
rect 9624 50161 9680 50164
rect 9732 50161 9788 50164
rect 9840 50161 10253 50164
rect 10305 50161 10361 50164
rect 10413 50161 10469 50164
rect 10521 50161 10577 50164
rect 10629 50161 10685 50164
rect 10737 50161 10793 50164
rect 10845 50161 10901 50164
rect 10953 50161 11009 50164
rect 11061 50161 11117 50164
rect 11169 50161 11225 50164
rect 11277 50161 11333 50164
rect 11385 50161 11441 50164
rect 11493 50161 11549 50164
rect 11601 50161 11657 50164
rect 3321 50115 3330 50161
rect 11648 50115 11657 50161
rect 3321 50112 3377 50115
rect 3429 50112 3485 50115
rect 3537 50112 3593 50115
rect 3645 50112 3701 50115
rect 3753 50112 3809 50115
rect 3861 50112 3917 50115
rect 3969 50112 4025 50115
rect 4077 50112 4133 50115
rect 4185 50112 4241 50115
rect 4293 50112 4349 50115
rect 4401 50112 4457 50115
rect 4509 50112 4565 50115
rect 4617 50112 4673 50115
rect 4725 50112 5138 50115
rect 5190 50112 5246 50115
rect 5298 50112 5354 50115
rect 5406 50112 5462 50115
rect 5514 50112 5570 50115
rect 5622 50112 5678 50115
rect 5730 50112 5786 50115
rect 5838 50112 5894 50115
rect 5946 50112 6002 50115
rect 6054 50112 6110 50115
rect 6162 50112 6218 50115
rect 6270 50112 6326 50115
rect 6378 50112 6434 50115
rect 6486 50112 6542 50115
rect 6594 50112 6650 50115
rect 6702 50112 6758 50115
rect 6810 50112 6866 50115
rect 6918 50112 6974 50115
rect 7026 50112 7082 50115
rect 7134 50112 7844 50115
rect 7896 50112 7952 50115
rect 8004 50112 8060 50115
rect 8112 50112 8168 50115
rect 8220 50112 8276 50115
rect 8328 50112 8384 50115
rect 8436 50112 8492 50115
rect 8544 50112 8600 50115
rect 8652 50112 8708 50115
rect 8760 50112 8816 50115
rect 8868 50112 8924 50115
rect 8976 50112 9032 50115
rect 9084 50112 9140 50115
rect 9192 50112 9248 50115
rect 9300 50112 9356 50115
rect 9408 50112 9464 50115
rect 9516 50112 9572 50115
rect 9624 50112 9680 50115
rect 9732 50112 9788 50115
rect 9840 50112 10253 50115
rect 10305 50112 10361 50115
rect 10413 50112 10469 50115
rect 10521 50112 10577 50115
rect 10629 50112 10685 50115
rect 10737 50112 10793 50115
rect 10845 50112 10901 50115
rect 10953 50112 11009 50115
rect 11061 50112 11117 50115
rect 11169 50112 11225 50115
rect 11277 50112 11333 50115
rect 11385 50112 11441 50115
rect 11493 50112 11549 50115
rect 11601 50112 11657 50115
rect 11709 50112 11765 50164
rect 3162 50056 11816 50112
rect 3213 50004 3269 50056
rect 3321 50004 3377 50056
rect 3429 50007 3485 50056
rect 3537 50007 3593 50056
rect 3645 50007 3701 50056
rect 3753 50007 3809 50056
rect 3861 50007 3917 50056
rect 3969 50007 4025 50056
rect 4077 50007 4133 50056
rect 4185 50007 4241 50056
rect 4293 50007 4349 50056
rect 4401 50007 4457 50056
rect 4509 50007 4565 50056
rect 4617 50007 4673 50056
rect 4725 50007 5138 50056
rect 5190 50007 5246 50056
rect 5298 50007 5354 50056
rect 5406 50007 5462 50056
rect 5514 50007 5570 50056
rect 5622 50007 5678 50056
rect 5730 50007 5786 50056
rect 5838 50007 5894 50056
rect 5946 50007 6002 50056
rect 6054 50007 6110 50056
rect 6162 50007 6218 50056
rect 6270 50007 6326 50056
rect 6378 50007 6434 50056
rect 6486 50007 6542 50056
rect 6594 50007 6650 50056
rect 6702 50007 6758 50056
rect 6810 50007 6866 50056
rect 6918 50007 6974 50056
rect 7026 50007 7082 50056
rect 7134 50007 7844 50056
rect 7896 50007 7952 50056
rect 8004 50007 8060 50056
rect 8112 50007 8168 50056
rect 8220 50007 8276 50056
rect 8328 50007 8384 50056
rect 8436 50007 8492 50056
rect 8544 50007 8600 50056
rect 8652 50007 8708 50056
rect 8760 50007 8816 50056
rect 8868 50007 8924 50056
rect 8976 50007 9032 50056
rect 9084 50007 9140 50056
rect 9192 50007 9248 50056
rect 9300 50007 9356 50056
rect 9408 50007 9464 50056
rect 9516 50007 9572 50056
rect 9624 50007 9680 50056
rect 9732 50007 9788 50056
rect 9840 50007 10253 50056
rect 10305 50007 10361 50056
rect 10413 50007 10469 50056
rect 10521 50007 10577 50056
rect 10629 50007 10685 50056
rect 10737 50007 10793 50056
rect 10845 50007 10901 50056
rect 10953 50007 11009 50056
rect 11061 50007 11117 50056
rect 11169 50007 11225 50056
rect 11277 50007 11333 50056
rect 11385 50007 11441 50056
rect 11493 50007 11549 50056
rect 11601 50004 11657 50056
rect 11709 50004 11765 50056
rect 3162 49976 3424 50004
rect 3162 49366 3270 49976
rect 3316 49961 3424 49976
rect 11554 49976 11816 50004
rect 11554 49961 11662 49976
rect 3316 49950 11662 49961
rect 3316 49392 3327 49950
rect 3489 49758 11489 49771
rect 3489 49712 3502 49758
rect 11476 49712 11489 49758
rect 3489 49699 4871 49712
rect 4923 49699 4979 49712
rect 5031 49699 7247 49712
rect 7299 49699 7355 49712
rect 7407 49699 7463 49712
rect 7515 49699 7571 49712
rect 7623 49699 7679 49712
rect 7731 49699 9947 49712
rect 9999 49699 10055 49712
rect 10107 49699 11489 49712
rect 3489 49643 11489 49699
rect 3489 49630 4871 49643
rect 4923 49630 4979 49643
rect 5031 49630 7247 49643
rect 7299 49630 7355 49643
rect 7407 49630 7463 49643
rect 7515 49630 7571 49643
rect 7623 49630 7679 49643
rect 7731 49630 9947 49643
rect 9999 49630 10055 49643
rect 10107 49630 11489 49643
rect 3489 49584 3502 49630
rect 11476 49584 11489 49630
rect 3489 49571 11489 49584
rect 11651 49392 11662 49950
rect 3316 49381 11662 49392
rect 3316 49366 3424 49381
rect 3162 49338 3424 49366
rect 11554 49366 11662 49381
rect 11708 49366 11816 49976
rect 11554 49338 11816 49366
rect 3213 49286 3269 49338
rect 3321 49286 3377 49338
rect 3429 49286 3485 49335
rect 3537 49286 3593 49335
rect 3645 49286 3701 49335
rect 3753 49286 3809 49335
rect 3861 49286 3917 49335
rect 3969 49286 4025 49335
rect 4077 49286 4133 49335
rect 4185 49286 4241 49335
rect 4293 49286 4349 49335
rect 4401 49286 4457 49335
rect 4509 49286 4565 49335
rect 4617 49286 4673 49335
rect 4725 49286 5138 49335
rect 5190 49286 5246 49335
rect 5298 49286 5354 49335
rect 5406 49286 5462 49335
rect 5514 49286 5570 49335
rect 5622 49286 5678 49335
rect 5730 49286 5786 49335
rect 5838 49286 5894 49335
rect 5946 49286 6002 49335
rect 6054 49286 6110 49335
rect 6162 49286 6218 49335
rect 6270 49286 6326 49335
rect 6378 49286 6434 49335
rect 6486 49286 6542 49335
rect 6594 49286 6650 49335
rect 6702 49286 6758 49335
rect 6810 49286 6866 49335
rect 6918 49286 6974 49335
rect 7026 49286 7082 49335
rect 7134 49286 7844 49335
rect 7896 49286 7952 49335
rect 8004 49286 8060 49335
rect 8112 49286 8168 49335
rect 8220 49286 8276 49335
rect 8328 49286 8384 49335
rect 8436 49286 8492 49335
rect 8544 49286 8600 49335
rect 8652 49286 8708 49335
rect 8760 49286 8816 49335
rect 8868 49286 8924 49335
rect 8976 49286 9032 49335
rect 9084 49286 9140 49335
rect 9192 49286 9248 49335
rect 9300 49286 9356 49335
rect 9408 49286 9464 49335
rect 9516 49286 9572 49335
rect 9624 49286 9680 49335
rect 9732 49286 9788 49335
rect 9840 49286 10253 49335
rect 10305 49286 10361 49335
rect 10413 49286 10469 49335
rect 10521 49286 10577 49335
rect 10629 49286 10685 49335
rect 10737 49286 10793 49335
rect 10845 49286 10901 49335
rect 10953 49286 11009 49335
rect 11061 49286 11117 49335
rect 11169 49286 11225 49335
rect 11277 49286 11333 49335
rect 11385 49286 11441 49335
rect 11493 49286 11549 49335
rect 11601 49286 11657 49338
rect 11709 49286 11765 49338
rect 3162 49230 11816 49286
rect 3213 49178 3269 49230
rect 3321 49227 3377 49230
rect 3429 49227 3485 49230
rect 3537 49227 3593 49230
rect 3645 49227 3701 49230
rect 3753 49227 3809 49230
rect 3861 49227 3917 49230
rect 3969 49227 4025 49230
rect 4077 49227 4133 49230
rect 4185 49227 4241 49230
rect 4293 49227 4349 49230
rect 4401 49227 4457 49230
rect 4509 49227 4565 49230
rect 4617 49227 4673 49230
rect 4725 49227 5138 49230
rect 5190 49227 5246 49230
rect 5298 49227 5354 49230
rect 5406 49227 5462 49230
rect 5514 49227 5570 49230
rect 5622 49227 5678 49230
rect 5730 49227 5786 49230
rect 5838 49227 5894 49230
rect 5946 49227 6002 49230
rect 6054 49227 6110 49230
rect 6162 49227 6218 49230
rect 6270 49227 6326 49230
rect 6378 49227 6434 49230
rect 6486 49227 6542 49230
rect 6594 49227 6650 49230
rect 6702 49227 6758 49230
rect 6810 49227 6866 49230
rect 6918 49227 6974 49230
rect 7026 49227 7082 49230
rect 7134 49227 7844 49230
rect 7896 49227 7952 49230
rect 8004 49227 8060 49230
rect 8112 49227 8168 49230
rect 8220 49227 8276 49230
rect 8328 49227 8384 49230
rect 8436 49227 8492 49230
rect 8544 49227 8600 49230
rect 8652 49227 8708 49230
rect 8760 49227 8816 49230
rect 8868 49227 8924 49230
rect 8976 49227 9032 49230
rect 9084 49227 9140 49230
rect 9192 49227 9248 49230
rect 9300 49227 9356 49230
rect 9408 49227 9464 49230
rect 9516 49227 9572 49230
rect 9624 49227 9680 49230
rect 9732 49227 9788 49230
rect 9840 49227 10253 49230
rect 10305 49227 10361 49230
rect 10413 49227 10469 49230
rect 10521 49227 10577 49230
rect 10629 49227 10685 49230
rect 10737 49227 10793 49230
rect 10845 49227 10901 49230
rect 10953 49227 11009 49230
rect 11061 49227 11117 49230
rect 11169 49227 11225 49230
rect 11277 49227 11333 49230
rect 11385 49227 11441 49230
rect 11493 49227 11549 49230
rect 11601 49227 11657 49230
rect 3321 49181 3330 49227
rect 11648 49181 11657 49227
rect 3321 49178 3377 49181
rect 3429 49178 3485 49181
rect 3537 49178 3593 49181
rect 3645 49178 3701 49181
rect 3753 49178 3809 49181
rect 3861 49178 3917 49181
rect 3969 49178 4025 49181
rect 4077 49178 4133 49181
rect 4185 49178 4241 49181
rect 4293 49178 4349 49181
rect 4401 49178 4457 49181
rect 4509 49178 4565 49181
rect 4617 49178 4673 49181
rect 4725 49178 5138 49181
rect 5190 49178 5246 49181
rect 5298 49178 5354 49181
rect 5406 49178 5462 49181
rect 5514 49178 5570 49181
rect 5622 49178 5678 49181
rect 5730 49178 5786 49181
rect 5838 49178 5894 49181
rect 5946 49178 6002 49181
rect 6054 49178 6110 49181
rect 6162 49178 6218 49181
rect 6270 49178 6326 49181
rect 6378 49178 6434 49181
rect 6486 49178 6542 49181
rect 6594 49178 6650 49181
rect 6702 49178 6758 49181
rect 6810 49178 6866 49181
rect 6918 49178 6974 49181
rect 7026 49178 7082 49181
rect 7134 49178 7844 49181
rect 7896 49178 7952 49181
rect 8004 49178 8060 49181
rect 8112 49178 8168 49181
rect 8220 49178 8276 49181
rect 8328 49178 8384 49181
rect 8436 49178 8492 49181
rect 8544 49178 8600 49181
rect 8652 49178 8708 49181
rect 8760 49178 8816 49181
rect 8868 49178 8924 49181
rect 8976 49178 9032 49181
rect 9084 49178 9140 49181
rect 9192 49178 9248 49181
rect 9300 49178 9356 49181
rect 9408 49178 9464 49181
rect 9516 49178 9572 49181
rect 9624 49178 9680 49181
rect 9732 49178 9788 49181
rect 9840 49178 10253 49181
rect 10305 49178 10361 49181
rect 10413 49178 10469 49181
rect 10521 49178 10577 49181
rect 10629 49178 10685 49181
rect 10737 49178 10793 49181
rect 10845 49178 10901 49181
rect 10953 49178 11009 49181
rect 11061 49178 11117 49181
rect 11169 49178 11225 49181
rect 11277 49178 11333 49181
rect 11385 49178 11441 49181
rect 11493 49178 11549 49181
rect 11601 49178 11657 49181
rect 11709 49178 11765 49230
rect 3162 49122 11816 49178
rect 3213 49070 3269 49122
rect 3321 49070 3377 49122
rect 3429 49073 3485 49122
rect 3537 49073 3593 49122
rect 3645 49073 3701 49122
rect 3753 49073 3809 49122
rect 3861 49073 3917 49122
rect 3969 49073 4025 49122
rect 4077 49073 4133 49122
rect 4185 49073 4241 49122
rect 4293 49073 4349 49122
rect 4401 49073 4457 49122
rect 4509 49073 4565 49122
rect 4617 49073 4673 49122
rect 4725 49073 5138 49122
rect 5190 49073 5246 49122
rect 5298 49073 5354 49122
rect 5406 49073 5462 49122
rect 5514 49073 5570 49122
rect 5622 49073 5678 49122
rect 5730 49073 5786 49122
rect 5838 49073 5894 49122
rect 5946 49073 6002 49122
rect 6054 49073 6110 49122
rect 6162 49073 6218 49122
rect 6270 49073 6326 49122
rect 6378 49073 6434 49122
rect 6486 49073 6542 49122
rect 6594 49073 6650 49122
rect 6702 49073 6758 49122
rect 6810 49073 6866 49122
rect 6918 49073 6974 49122
rect 7026 49073 7082 49122
rect 7134 49073 7844 49122
rect 7896 49073 7952 49122
rect 8004 49073 8060 49122
rect 8112 49073 8168 49122
rect 8220 49073 8276 49122
rect 8328 49073 8384 49122
rect 8436 49073 8492 49122
rect 8544 49073 8600 49122
rect 8652 49073 8708 49122
rect 8760 49073 8816 49122
rect 8868 49073 8924 49122
rect 8976 49073 9032 49122
rect 9084 49073 9140 49122
rect 9192 49073 9248 49122
rect 9300 49073 9356 49122
rect 9408 49073 9464 49122
rect 9516 49073 9572 49122
rect 9624 49073 9680 49122
rect 9732 49073 9788 49122
rect 9840 49073 10253 49122
rect 10305 49073 10361 49122
rect 10413 49073 10469 49122
rect 10521 49073 10577 49122
rect 10629 49073 10685 49122
rect 10737 49073 10793 49122
rect 10845 49073 10901 49122
rect 10953 49073 11009 49122
rect 11061 49073 11117 49122
rect 11169 49073 11225 49122
rect 11277 49073 11333 49122
rect 11385 49073 11441 49122
rect 11493 49073 11549 49122
rect 11601 49070 11657 49122
rect 11709 49070 11765 49122
rect 3162 49042 3424 49070
rect 3162 48432 3270 49042
rect 3316 49027 3424 49042
rect 11554 49042 11816 49070
rect 11554 49027 11662 49042
rect 3316 49016 11662 49027
rect 3316 48458 3327 49016
rect 3489 48824 11489 48837
rect 3489 48778 3502 48824
rect 11476 48778 11489 48824
rect 3489 48765 4871 48778
rect 4923 48765 4979 48778
rect 5031 48765 7247 48778
rect 7299 48765 7355 48778
rect 7407 48765 7463 48778
rect 7515 48765 7571 48778
rect 7623 48765 7679 48778
rect 7731 48765 9947 48778
rect 9999 48765 10055 48778
rect 10107 48765 11489 48778
rect 3489 48709 11489 48765
rect 3489 48696 4871 48709
rect 4923 48696 4979 48709
rect 5031 48696 7247 48709
rect 7299 48696 7355 48709
rect 7407 48696 7463 48709
rect 7515 48696 7571 48709
rect 7623 48696 7679 48709
rect 7731 48696 9947 48709
rect 9999 48696 10055 48709
rect 10107 48696 11489 48709
rect 3489 48650 3502 48696
rect 11476 48650 11489 48696
rect 3489 48637 11489 48650
rect 11651 48458 11662 49016
rect 3316 48447 11662 48458
rect 3316 48432 3424 48447
rect 3162 48427 3424 48432
rect 11554 48432 11662 48447
rect 11708 48432 11816 49042
rect 11554 48427 11816 48432
rect 3105 48375 3161 48376
rect 3213 48375 3269 48427
rect 3321 48375 3377 48427
rect 3429 48375 3485 48401
rect 3537 48375 3593 48401
rect 3645 48375 3701 48401
rect 3753 48375 3809 48401
rect 3861 48375 3917 48401
rect 3969 48375 4025 48401
rect 4077 48375 4133 48401
rect 4185 48375 4241 48401
rect 4293 48375 4349 48401
rect 4401 48375 4457 48401
rect 4509 48375 4565 48401
rect 4617 48375 4673 48401
rect 4725 48375 5138 48401
rect 5190 48375 5246 48401
rect 5298 48375 5354 48401
rect 5406 48375 5462 48401
rect 5514 48375 5570 48401
rect 5622 48375 5678 48401
rect 5730 48375 5786 48401
rect 5838 48375 5894 48401
rect 5946 48375 6002 48401
rect 6054 48375 6110 48401
rect 6162 48375 6218 48401
rect 6270 48375 6326 48401
rect 6378 48375 6434 48401
rect 6486 48375 6542 48401
rect 6594 48375 6650 48401
rect 6702 48375 6758 48401
rect 6810 48375 6866 48401
rect 6918 48375 6974 48401
rect 7026 48375 7082 48401
rect 7134 48375 7844 48401
rect 7896 48375 7952 48401
rect 8004 48375 8060 48401
rect 8112 48375 8168 48401
rect 8220 48375 8276 48401
rect 8328 48375 8384 48401
rect 8436 48375 8492 48401
rect 8544 48375 8600 48401
rect 8652 48375 8708 48401
rect 8760 48375 8816 48401
rect 8868 48375 8924 48401
rect 8976 48375 9032 48401
rect 9084 48375 9140 48401
rect 9192 48375 9248 48401
rect 9300 48375 9356 48401
rect 9408 48375 9464 48401
rect 9516 48375 9572 48401
rect 9624 48375 9680 48401
rect 9732 48375 9788 48401
rect 9840 48375 10253 48401
rect 10305 48375 10361 48401
rect 10413 48375 10469 48401
rect 10521 48375 10577 48401
rect 10629 48375 10685 48401
rect 10737 48375 10793 48401
rect 10845 48375 10901 48401
rect 10953 48375 11009 48401
rect 11061 48375 11117 48401
rect 11169 48375 11225 48401
rect 11277 48375 11333 48401
rect 11385 48375 11441 48401
rect 11493 48375 11549 48401
rect 11601 48375 11657 48427
rect 11709 48375 11765 48427
rect 11862 48376 11873 51900
rect 11817 48375 11873 48376
rect 3105 48319 11873 48375
rect 3105 48293 3161 48319
rect 3213 48293 3269 48319
rect 3321 48293 3377 48319
rect 3429 48293 3485 48319
rect 3537 48293 3593 48319
rect 3645 48293 3701 48319
rect 3753 48293 3809 48319
rect 3861 48293 3917 48319
rect 3969 48293 4025 48319
rect 4077 48293 4133 48319
rect 4185 48293 4241 48319
rect 4293 48293 4349 48319
rect 4401 48293 4457 48319
rect 4509 48293 4565 48319
rect 4617 48293 4673 48319
rect 4725 48293 5138 48319
rect 5190 48293 5246 48319
rect 5298 48293 5354 48319
rect 5406 48293 5462 48319
rect 5514 48293 5570 48319
rect 5622 48293 5678 48319
rect 5730 48293 5786 48319
rect 5838 48293 5894 48319
rect 5946 48293 6002 48319
rect 6054 48293 6110 48319
rect 6162 48293 6218 48319
rect 6270 48293 6326 48319
rect 6378 48293 6434 48319
rect 6486 48293 6542 48319
rect 6594 48293 6650 48319
rect 6702 48293 6758 48319
rect 6810 48293 6866 48319
rect 6918 48293 6974 48319
rect 7026 48293 7082 48319
rect 7134 48293 7844 48319
rect 7896 48293 7952 48319
rect 8004 48293 8060 48319
rect 8112 48293 8168 48319
rect 8220 48293 8276 48319
rect 8328 48293 8384 48319
rect 8436 48293 8492 48319
rect 8544 48293 8600 48319
rect 8652 48293 8708 48319
rect 8760 48293 8816 48319
rect 8868 48293 8924 48319
rect 8976 48293 9032 48319
rect 9084 48293 9140 48319
rect 9192 48293 9248 48319
rect 9300 48293 9356 48319
rect 9408 48293 9464 48319
rect 9516 48293 9572 48319
rect 9624 48293 9680 48319
rect 9732 48293 9788 48319
rect 9840 48293 10253 48319
rect 10305 48293 10361 48319
rect 10413 48293 10469 48319
rect 10521 48293 10577 48319
rect 10629 48293 10685 48319
rect 10737 48293 10793 48319
rect 10845 48293 10901 48319
rect 10953 48293 11009 48319
rect 11061 48293 11117 48319
rect 11169 48293 11225 48319
rect 11277 48293 11333 48319
rect 11385 48293 11441 48319
rect 11493 48293 11549 48319
rect 11601 48293 11657 48319
rect 11709 48293 11765 48319
rect 11817 48293 11873 48319
rect 3105 48247 3142 48293
rect 11836 48247 11873 48293
rect 3105 48236 11873 48247
rect 12059 48022 12070 52254
rect 2908 48011 12070 48022
rect 2908 47665 3016 48011
rect 11962 47665 12070 48011
rect 12416 47665 12427 52611
rect 2551 47654 12427 47665
rect 12753 52611 14907 52622
rect 12753 47665 12764 52611
rect 14710 52586 14907 52611
rect 14710 52574 14968 52586
rect 14710 52522 14904 52574
rect 14956 52522 14968 52574
rect 14710 52466 14968 52522
rect 14710 52414 14904 52466
rect 14956 52414 14968 52466
rect 14710 52358 14968 52414
rect 14710 52306 14904 52358
rect 14956 52306 14968 52358
rect 14710 52250 14968 52306
rect 14710 52198 14904 52250
rect 14956 52198 14968 52250
rect 14710 52142 14968 52198
rect 14710 52090 14904 52142
rect 14956 52090 14968 52142
rect 14710 52034 14968 52090
rect 14710 51982 14904 52034
rect 14956 51982 14968 52034
rect 14710 51926 14968 51982
rect 14710 51874 14904 51926
rect 14956 51874 14968 51926
rect 14710 51818 14968 51874
rect 14710 51766 14904 51818
rect 14956 51766 14968 51818
rect 14710 51710 14968 51766
rect 14710 51658 14904 51710
rect 14956 51658 14968 51710
rect 14710 51622 14968 51658
rect 14710 51422 14721 51622
rect 14892 51602 14968 51622
rect 14892 51550 14904 51602
rect 14956 51550 14968 51602
rect 14892 51494 14968 51550
rect 14892 51442 14904 51494
rect 14956 51442 14968 51494
rect 14892 51422 14968 51442
rect 14710 51386 14968 51422
rect 14710 51334 14904 51386
rect 14956 51334 14968 51386
rect 14710 51278 14968 51334
rect 14710 51226 14904 51278
rect 14956 51226 14968 51278
rect 14710 51214 14968 51226
rect 14710 50422 14907 51214
rect 14710 49854 14721 50422
rect 14710 49386 14907 49854
rect 14710 49374 14968 49386
rect 14710 49322 14904 49374
rect 14956 49322 14968 49374
rect 14710 49266 14968 49322
rect 14710 49214 14904 49266
rect 14956 49214 14968 49266
rect 14710 49158 14968 49214
rect 14710 49106 14904 49158
rect 14956 49106 14968 49158
rect 14710 49050 14968 49106
rect 14710 48998 14904 49050
rect 14956 48998 14968 49050
rect 14710 48942 14968 48998
rect 14710 48890 14904 48942
rect 14956 48890 14968 48942
rect 14710 48854 14968 48890
rect 14710 48654 14721 48854
rect 14892 48834 14968 48854
rect 14892 48782 14904 48834
rect 14956 48782 14968 48834
rect 14892 48726 14968 48782
rect 14892 48674 14904 48726
rect 14956 48674 14968 48726
rect 14892 48654 14968 48674
rect 14710 48618 14968 48654
rect 14710 48566 14904 48618
rect 14956 48566 14968 48618
rect 14710 48510 14968 48566
rect 14710 48458 14904 48510
rect 14956 48458 14968 48510
rect 14710 48402 14968 48458
rect 14710 48350 14904 48402
rect 14956 48350 14968 48402
rect 14710 48294 14968 48350
rect 14710 48242 14904 48294
rect 14956 48242 14968 48294
rect 14710 48186 14968 48242
rect 14710 48134 14904 48186
rect 14956 48134 14968 48186
rect 14710 48078 14968 48134
rect 14710 48026 14904 48078
rect 14956 48026 14968 48078
rect 14710 48014 14968 48026
rect 14710 47665 14907 48014
rect 12753 47654 14907 47665
rect 10 46174 86 46186
rect 10 46122 22 46174
rect 74 46122 86 46174
rect 10 46066 86 46122
rect 10 46014 22 46066
rect 74 46014 86 46066
rect 10 45958 86 46014
rect 10 45906 22 45958
rect 74 45906 86 45958
rect 10 45850 86 45906
rect 10 45798 22 45850
rect 74 45798 86 45850
rect 10 45742 86 45798
rect 10 45690 22 45742
rect 74 45690 86 45742
rect 10 45634 86 45690
rect 10 45582 22 45634
rect 74 45582 86 45634
rect 10 45526 86 45582
rect 10 45474 22 45526
rect 74 45474 86 45526
rect 10 45418 86 45474
rect 10 45366 22 45418
rect 74 45366 86 45418
rect 10 45310 86 45366
rect 10 45258 22 45310
rect 74 45258 86 45310
rect 10 45202 86 45258
rect 10 45150 22 45202
rect 74 45150 86 45202
rect 10 45094 86 45150
rect 10 45042 22 45094
rect 74 45042 86 45094
rect 10 44986 86 45042
rect 10 44934 22 44986
rect 74 44934 86 44986
rect 10 44878 86 44934
rect 10 44826 22 44878
rect 74 44826 86 44878
rect 10 44814 86 44826
rect 14892 46174 14968 46186
rect 14892 46122 14904 46174
rect 14956 46122 14968 46174
rect 14892 46066 14968 46122
rect 14892 46014 14904 46066
rect 14956 46014 14968 46066
rect 14892 45958 14968 46014
rect 14892 45906 14904 45958
rect 14956 45906 14968 45958
rect 14892 45850 14968 45906
rect 14892 45798 14904 45850
rect 14956 45798 14968 45850
rect 14892 45742 14968 45798
rect 14892 45690 14904 45742
rect 14956 45690 14968 45742
rect 14892 45634 14968 45690
rect 14892 45582 14904 45634
rect 14956 45582 14968 45634
rect 14892 45526 14968 45582
rect 14892 45474 14904 45526
rect 14956 45474 14968 45526
rect 14892 45418 14968 45474
rect 14892 45366 14904 45418
rect 14956 45366 14968 45418
rect 14892 45310 14968 45366
rect 14892 45258 14904 45310
rect 14956 45258 14968 45310
rect 14892 45202 14968 45258
rect 14892 45150 14904 45202
rect 14956 45150 14968 45202
rect 14892 45094 14968 45150
rect 14892 45042 14904 45094
rect 14956 45042 14968 45094
rect 14892 44986 14968 45042
rect 14892 44934 14904 44986
rect 14956 44934 14968 44986
rect 14892 44878 14968 44934
rect 14892 44826 14904 44878
rect 14956 44826 14968 44878
rect 14892 44814 14968 44826
rect 71 42647 725 42658
rect 71 41658 268 42647
rect 257 41458 268 41658
rect 71 40458 268 41458
rect 257 40258 268 40458
rect 71 39258 268 40258
rect 257 39058 268 39258
rect 71 38186 268 39058
rect 10 38174 268 38186
rect 10 38122 22 38174
rect 74 38122 268 38174
rect 10 38066 268 38122
rect 10 38014 22 38066
rect 74 38058 268 38066
rect 74 38014 86 38058
rect 10 37958 86 38014
rect 10 37906 22 37958
rect 74 37906 86 37958
rect 10 37858 86 37906
rect 257 37858 268 38058
rect 10 37850 268 37858
rect 10 37798 22 37850
rect 74 37798 268 37850
rect 10 37742 268 37798
rect 10 37690 22 37742
rect 74 37690 268 37742
rect 10 37634 268 37690
rect 10 37582 22 37634
rect 74 37582 268 37634
rect 10 37526 268 37582
rect 10 37474 22 37526
rect 74 37474 268 37526
rect 10 37418 268 37474
rect 10 37366 22 37418
rect 74 37366 268 37418
rect 10 37310 268 37366
rect 10 37258 22 37310
rect 74 37258 268 37310
rect 10 37202 268 37258
rect 10 37150 22 37202
rect 74 37150 268 37202
rect 10 37094 268 37150
rect 10 37042 22 37094
rect 74 37042 268 37094
rect 10 36986 268 37042
rect 10 36934 22 36986
rect 74 36934 268 36986
rect 10 36878 268 36934
rect 10 36826 22 36878
rect 74 36858 268 36878
rect 74 36826 86 36858
rect 10 36814 86 36826
rect 257 36658 268 36858
rect 71 36596 268 36658
rect 10 36584 268 36596
rect 10 36532 22 36584
rect 74 36532 268 36584
rect 10 36476 268 36532
rect 10 36424 22 36476
rect 74 36424 268 36476
rect 10 36368 268 36424
rect 10 36316 22 36368
rect 74 36316 268 36368
rect 10 36260 268 36316
rect 10 36208 22 36260
rect 74 36208 268 36260
rect 10 36152 268 36208
rect 10 36100 22 36152
rect 74 36100 268 36152
rect 10 36044 268 36100
rect 10 35992 22 36044
rect 74 35992 268 36044
rect 10 35936 268 35992
rect 10 35884 22 35936
rect 74 35884 268 35936
rect 10 35828 268 35884
rect 10 35776 22 35828
rect 74 35776 268 35828
rect 10 35720 268 35776
rect 10 35668 22 35720
rect 74 35668 268 35720
rect 10 35658 268 35668
rect 10 35612 86 35658
rect 10 35560 22 35612
rect 74 35560 86 35612
rect 10 35504 86 35560
rect 10 35452 22 35504
rect 74 35458 86 35504
rect 257 35458 268 35658
rect 74 35452 268 35458
rect 10 35396 268 35452
rect 10 35344 22 35396
rect 74 35344 268 35396
rect 10 35288 268 35344
rect 10 35236 22 35288
rect 74 35236 268 35288
rect 10 35180 268 35236
rect 10 35128 22 35180
rect 74 35128 268 35180
rect 10 35072 268 35128
rect 10 35020 22 35072
rect 74 35020 268 35072
rect 10 34964 268 35020
rect 10 34912 22 34964
rect 74 34912 268 34964
rect 10 34856 268 34912
rect 10 34804 22 34856
rect 74 34804 268 34856
rect 10 34748 268 34804
rect 10 34696 22 34748
rect 74 34696 268 34748
rect 10 34640 268 34696
rect 10 34588 22 34640
rect 74 34588 268 34640
rect 10 34532 268 34588
rect 10 34480 22 34532
rect 74 34480 268 34532
rect 10 34458 268 34480
rect 10 34424 86 34458
rect 10 34372 22 34424
rect 74 34372 86 34424
rect 10 34316 86 34372
rect 10 34264 22 34316
rect 74 34264 86 34316
rect 10 34258 86 34264
rect 257 34258 268 34458
rect 10 34208 268 34258
rect 10 34156 22 34208
rect 74 34156 268 34208
rect 10 34100 268 34156
rect 10 34048 22 34100
rect 74 34048 268 34100
rect 10 33992 268 34048
rect 10 33940 22 33992
rect 74 33940 268 33992
rect 10 33884 268 33940
rect 10 33832 22 33884
rect 74 33832 268 33884
rect 10 33776 268 33832
rect 10 33724 22 33776
rect 74 33724 268 33776
rect 10 33668 268 33724
rect 10 33616 22 33668
rect 74 33616 268 33668
rect 10 33604 268 33616
rect 71 33258 268 33604
rect 257 33058 268 33258
rect 71 32058 268 33058
rect 257 31858 268 32058
rect 71 30858 268 31858
rect 257 30658 268 30858
rect 71 29658 268 30658
rect 257 29458 268 29658
rect 71 28586 268 29458
rect 10 28574 268 28586
rect 10 28522 22 28574
rect 74 28522 268 28574
rect 10 28466 268 28522
rect 10 28414 22 28466
rect 74 28458 268 28466
rect 74 28414 86 28458
rect 10 28358 86 28414
rect 10 28306 22 28358
rect 74 28306 86 28358
rect 10 28258 86 28306
rect 257 28258 268 28458
rect 10 28250 268 28258
rect 10 28198 22 28250
rect 74 28198 268 28250
rect 10 28142 268 28198
rect 10 28090 22 28142
rect 74 28090 268 28142
rect 10 28034 268 28090
rect 10 27982 22 28034
rect 74 27982 268 28034
rect 10 27926 268 27982
rect 10 27874 22 27926
rect 74 27874 268 27926
rect 10 27818 268 27874
rect 10 27766 22 27818
rect 74 27766 268 27818
rect 10 27710 268 27766
rect 10 27658 22 27710
rect 74 27658 268 27710
rect 10 27602 268 27658
rect 10 27550 22 27602
rect 74 27550 268 27602
rect 10 27494 268 27550
rect 10 27442 22 27494
rect 74 27442 268 27494
rect 10 27386 268 27442
rect 10 27334 22 27386
rect 74 27334 268 27386
rect 10 27278 268 27334
rect 10 27226 22 27278
rect 74 27258 268 27278
rect 74 27226 86 27258
rect 10 27214 86 27226
rect 257 27058 268 27258
rect 71 26058 268 27058
rect 257 25858 268 26058
rect 71 24858 268 25858
rect 257 24658 268 24858
rect 71 23658 268 24658
rect 257 23458 268 23658
rect 71 22458 268 23458
rect 257 21390 268 22458
rect 71 20390 268 21390
rect 257 20190 268 20390
rect 71 19190 268 20190
rect 257 18990 268 19190
rect 71 17990 268 18990
rect 257 17790 268 17990
rect 71 16790 268 17790
rect 257 16590 268 16790
rect 71 15590 268 16590
rect 257 15390 268 15590
rect 71 14390 268 15390
rect 257 14190 268 14390
rect 71 14186 268 14190
rect 10 14174 268 14186
rect 10 14122 22 14174
rect 74 14122 268 14174
rect 10 14066 268 14122
rect 10 14014 22 14066
rect 74 14014 268 14066
rect 10 13958 268 14014
rect 10 13906 22 13958
rect 74 13906 268 13958
rect 10 13850 268 13906
rect 10 13798 22 13850
rect 74 13798 268 13850
rect 10 13742 268 13798
rect 10 13690 22 13742
rect 74 13690 268 13742
rect 10 13634 268 13690
rect 10 13582 22 13634
rect 74 13582 268 13634
rect 10 13526 268 13582
rect 10 13474 22 13526
rect 74 13474 268 13526
rect 10 13418 268 13474
rect 10 13366 22 13418
rect 74 13366 268 13418
rect 10 13310 268 13366
rect 10 13258 22 13310
rect 74 13258 268 13310
rect 10 13202 268 13258
rect 10 13150 22 13202
rect 74 13190 268 13202
rect 74 13150 86 13190
rect 10 13094 86 13150
rect 10 13042 22 13094
rect 74 13042 86 13094
rect 10 12990 86 13042
rect 257 12990 268 13190
rect 10 12986 268 12990
rect 10 12934 22 12986
rect 74 12934 268 12986
rect 10 12878 268 12934
rect 10 12826 22 12878
rect 74 12826 268 12878
rect 10 12814 268 12826
rect 71 11990 268 12814
rect 257 11790 268 11990
rect 71 10996 268 11790
rect 10 10984 268 10996
rect 10 10932 22 10984
rect 74 10932 268 10984
rect 10 10876 268 10932
rect 10 10824 22 10876
rect 74 10824 268 10876
rect 10 10790 268 10824
rect 10 10768 86 10790
rect 10 10716 22 10768
rect 74 10716 86 10768
rect 10 10660 86 10716
rect 10 10608 22 10660
rect 74 10608 86 10660
rect 10 10590 86 10608
rect 257 10590 268 10790
rect 10 10552 268 10590
rect 10 10500 22 10552
rect 74 10500 268 10552
rect 10 10444 268 10500
rect 10 10392 22 10444
rect 74 10392 268 10444
rect 10 10336 268 10392
rect 10 10284 22 10336
rect 74 10284 268 10336
rect 10 10228 268 10284
rect 10 10176 22 10228
rect 74 10176 268 10228
rect 10 10120 268 10176
rect 10 10068 22 10120
rect 74 10068 268 10120
rect 10 10012 268 10068
rect 10 9960 22 10012
rect 74 9960 268 10012
rect 10 9904 268 9960
rect 10 9852 22 9904
rect 74 9852 268 9904
rect 10 9796 268 9852
rect 10 9744 22 9796
rect 74 9744 268 9796
rect 10 9688 268 9744
rect 10 9636 22 9688
rect 74 9636 268 9688
rect 10 9590 268 9636
rect 10 9580 86 9590
rect 10 9528 22 9580
rect 74 9528 86 9580
rect 10 9472 86 9528
rect 10 9420 22 9472
rect 74 9420 86 9472
rect 10 9390 86 9420
rect 257 9390 268 9590
rect 10 9364 268 9390
rect 10 9312 22 9364
rect 74 9312 268 9364
rect 10 9256 268 9312
rect 10 9204 22 9256
rect 74 9204 268 9256
rect 10 9148 268 9204
rect 10 9096 22 9148
rect 74 9096 268 9148
rect 10 9040 268 9096
rect 10 8988 22 9040
rect 74 8988 268 9040
rect 10 8932 268 8988
rect 10 8880 22 8932
rect 74 8880 268 8932
rect 10 8824 268 8880
rect 10 8772 22 8824
rect 74 8772 268 8824
rect 10 8716 268 8772
rect 10 8664 22 8716
rect 74 8664 268 8716
rect 10 8608 268 8664
rect 10 8556 22 8608
rect 74 8556 268 8608
rect 10 8500 268 8556
rect 10 8448 22 8500
rect 74 8448 268 8500
rect 10 8392 268 8448
rect 10 8340 22 8392
rect 74 8390 268 8392
rect 74 8340 86 8390
rect 10 8284 86 8340
rect 10 8232 22 8284
rect 74 8232 86 8284
rect 10 8190 86 8232
rect 257 8190 268 8390
rect 10 8176 268 8190
rect 10 8124 22 8176
rect 74 8124 268 8176
rect 10 8068 268 8124
rect 10 8016 22 8068
rect 74 8016 268 8068
rect 10 8004 268 8016
rect 71 7796 268 8004
rect 10 7784 268 7796
rect 10 7732 22 7784
rect 74 7732 268 7784
rect 10 7676 268 7732
rect 10 7624 22 7676
rect 74 7624 268 7676
rect 10 7568 268 7624
rect 10 7516 22 7568
rect 74 7516 268 7568
rect 10 7460 268 7516
rect 10 7408 22 7460
rect 74 7408 268 7460
rect 10 7352 268 7408
rect 10 7300 22 7352
rect 74 7300 268 7352
rect 10 7244 268 7300
rect 10 7192 22 7244
rect 74 7192 268 7244
rect 10 7190 268 7192
rect 10 7136 86 7190
rect 10 7084 22 7136
rect 74 7084 86 7136
rect 10 7028 86 7084
rect 10 6976 22 7028
rect 74 6990 86 7028
rect 257 6990 268 7190
rect 74 6976 268 6990
rect 10 6920 268 6976
rect 10 6868 22 6920
rect 74 6868 268 6920
rect 10 6812 268 6868
rect 10 6760 22 6812
rect 74 6760 268 6812
rect 10 6704 268 6760
rect 10 6652 22 6704
rect 74 6652 268 6704
rect 10 6596 268 6652
rect 10 6544 22 6596
rect 74 6544 268 6596
rect 10 6488 268 6544
rect 10 6436 22 6488
rect 74 6436 268 6488
rect 10 6380 268 6436
rect 10 6328 22 6380
rect 74 6328 268 6380
rect 10 6272 268 6328
rect 10 6220 22 6272
rect 74 6220 268 6272
rect 10 6164 268 6220
rect 10 6112 22 6164
rect 74 6112 268 6164
rect 10 6056 268 6112
rect 10 6004 22 6056
rect 74 6004 268 6056
rect 10 5990 268 6004
rect 10 5948 86 5990
rect 10 5896 22 5948
rect 74 5896 86 5948
rect 10 5840 86 5896
rect 10 5788 22 5840
rect 74 5790 86 5840
rect 257 5790 268 5990
rect 74 5788 268 5790
rect 10 5732 268 5788
rect 10 5680 22 5732
rect 74 5680 268 5732
rect 10 5624 268 5680
rect 10 5572 22 5624
rect 74 5572 268 5624
rect 10 5516 268 5572
rect 10 5464 22 5516
rect 74 5464 268 5516
rect 10 5408 268 5464
rect 10 5356 22 5408
rect 74 5356 268 5408
rect 10 5300 268 5356
rect 10 5248 22 5300
rect 74 5248 268 5300
rect 10 5192 268 5248
rect 10 5140 22 5192
rect 74 5140 268 5192
rect 10 5084 268 5140
rect 10 5032 22 5084
rect 74 5032 268 5084
rect 10 4976 268 5032
rect 10 4924 22 4976
rect 74 4924 268 4976
rect 10 4868 268 4924
rect 10 4816 22 4868
rect 74 4816 268 4868
rect 10 4804 268 4816
rect 71 4790 268 4804
rect 10 4590 86 4596
rect 257 4590 268 4790
rect 10 4584 268 4590
rect 10 4532 22 4584
rect 74 4532 268 4584
rect 10 4476 268 4532
rect 10 4424 22 4476
rect 74 4424 268 4476
rect 10 4368 268 4424
rect 10 4316 22 4368
rect 74 4316 268 4368
rect 10 4260 268 4316
rect 10 4208 22 4260
rect 74 4208 268 4260
rect 10 4152 268 4208
rect 10 4100 22 4152
rect 74 4100 268 4152
rect 10 4044 268 4100
rect 10 3992 22 4044
rect 74 3992 268 4044
rect 10 3936 268 3992
rect 10 3884 22 3936
rect 74 3884 268 3936
rect 10 3828 268 3884
rect 10 3776 22 3828
rect 74 3776 268 3828
rect 10 3720 268 3776
rect 10 3668 22 3720
rect 74 3668 268 3720
rect 10 3612 268 3668
rect 10 3560 22 3612
rect 74 3590 268 3612
rect 74 3560 86 3590
rect 10 3504 86 3560
rect 10 3452 22 3504
rect 74 3452 86 3504
rect 10 3396 86 3452
rect 10 3344 22 3396
rect 74 3390 86 3396
rect 257 3390 268 3590
rect 74 3344 268 3390
rect 10 3288 268 3344
rect 10 3236 22 3288
rect 74 3236 268 3288
rect 10 3180 268 3236
rect 10 3128 22 3180
rect 74 3128 268 3180
rect 10 3072 268 3128
rect 10 3020 22 3072
rect 74 3020 268 3072
rect 10 2964 268 3020
rect 10 2912 22 2964
rect 74 2912 268 2964
rect 10 2856 268 2912
rect 10 2804 22 2856
rect 74 2804 268 2856
rect 10 2748 268 2804
rect 10 2696 22 2748
rect 74 2696 268 2748
rect 10 2640 268 2696
rect 10 2588 22 2640
rect 74 2588 268 2640
rect 10 2532 268 2588
rect 10 2480 22 2532
rect 74 2480 268 2532
rect 10 2424 268 2480
rect 10 2372 22 2424
rect 74 2390 268 2424
rect 74 2372 86 2390
rect 10 2316 86 2372
rect 10 2264 22 2316
rect 74 2264 86 2316
rect 10 2208 86 2264
rect 10 2156 22 2208
rect 74 2190 86 2208
rect 257 2190 268 2390
rect 74 2156 268 2190
rect 10 2100 268 2156
rect 10 2048 22 2100
rect 74 2048 268 2100
rect 10 1992 268 2048
rect 10 1940 22 1992
rect 74 1940 268 1992
rect 10 1884 268 1940
rect 10 1832 22 1884
rect 74 1832 268 1884
rect 10 1776 268 1832
rect 10 1724 22 1776
rect 74 1724 268 1776
rect 10 1668 268 1724
rect 10 1616 22 1668
rect 74 1616 268 1668
rect 10 1604 268 1616
rect 71 1201 268 1604
rect 714 1201 725 42647
rect 13012 42647 14907 42658
rect 13012 27201 13023 42647
rect 13969 41658 14264 42647
rect 13969 41458 13980 41658
rect 14253 41458 14264 41658
rect 13969 40458 14264 41458
rect 13969 40258 13980 40458
rect 14253 40258 14264 40458
rect 13969 39258 14264 40258
rect 13969 39058 13980 39258
rect 14253 39058 14264 39258
rect 13969 38058 14264 39058
rect 13969 37858 13980 38058
rect 14253 37858 14264 38058
rect 13969 36858 14264 37858
rect 13969 36658 13980 36858
rect 14253 36658 14264 36858
rect 13969 35658 14264 36658
rect 13969 35458 13980 35658
rect 14253 35458 14264 35658
rect 13969 34458 14264 35458
rect 13969 34258 13980 34458
rect 14253 34258 14264 34458
rect 13969 33258 14264 34258
rect 13969 33058 13980 33258
rect 14253 33058 14264 33258
rect 13969 32058 14264 33058
rect 13969 31858 13980 32058
rect 14253 31858 14264 32058
rect 13969 30858 14264 31858
rect 13969 30658 13980 30858
rect 14253 30658 14264 30858
rect 13969 29658 14264 30658
rect 13969 29458 13980 29658
rect 14253 29458 14264 29658
rect 13969 28458 14264 29458
rect 13969 28190 13980 28458
rect 14253 28190 14264 28458
rect 13969 27201 14264 28190
rect 13012 27190 14264 27201
rect 71 1190 725 1201
rect 14253 1201 14264 27190
rect 14710 41658 14907 42647
rect 14710 41458 14721 41658
rect 14710 40458 14907 41458
rect 14710 40258 14721 40458
rect 14710 39258 14907 40258
rect 14710 39058 14721 39258
rect 14710 38186 14907 39058
rect 14710 38174 14968 38186
rect 14710 38122 14904 38174
rect 14956 38122 14968 38174
rect 14710 38066 14968 38122
rect 14710 38058 14904 38066
rect 14710 37858 14721 38058
rect 14892 38014 14904 38058
rect 14956 38014 14968 38066
rect 14892 37958 14968 38014
rect 14892 37906 14904 37958
rect 14956 37906 14968 37958
rect 14892 37858 14968 37906
rect 14710 37850 14968 37858
rect 14710 37798 14904 37850
rect 14956 37798 14968 37850
rect 14710 37742 14968 37798
rect 14710 37690 14904 37742
rect 14956 37690 14968 37742
rect 14710 37634 14968 37690
rect 14710 37582 14904 37634
rect 14956 37582 14968 37634
rect 14710 37526 14968 37582
rect 14710 37474 14904 37526
rect 14956 37474 14968 37526
rect 14710 37418 14968 37474
rect 14710 37366 14904 37418
rect 14956 37366 14968 37418
rect 14710 37310 14968 37366
rect 14710 37258 14904 37310
rect 14956 37258 14968 37310
rect 14710 37202 14968 37258
rect 14710 37150 14904 37202
rect 14956 37150 14968 37202
rect 14710 37094 14968 37150
rect 14710 37042 14904 37094
rect 14956 37042 14968 37094
rect 14710 36986 14968 37042
rect 14710 36934 14904 36986
rect 14956 36934 14968 36986
rect 14710 36878 14968 36934
rect 14710 36858 14904 36878
rect 14710 36658 14721 36858
rect 14892 36826 14904 36858
rect 14956 36826 14968 36878
rect 14892 36814 14968 36826
rect 14710 36596 14907 36658
rect 14710 36584 14968 36596
rect 14710 36532 14904 36584
rect 14956 36532 14968 36584
rect 14710 36476 14968 36532
rect 14710 36424 14904 36476
rect 14956 36424 14968 36476
rect 14710 36368 14968 36424
rect 14710 36316 14904 36368
rect 14956 36316 14968 36368
rect 14710 36260 14968 36316
rect 14710 36208 14904 36260
rect 14956 36208 14968 36260
rect 14710 36152 14968 36208
rect 14710 36100 14904 36152
rect 14956 36100 14968 36152
rect 14710 36044 14968 36100
rect 14710 35992 14904 36044
rect 14956 35992 14968 36044
rect 14710 35936 14968 35992
rect 14710 35884 14904 35936
rect 14956 35884 14968 35936
rect 14710 35828 14968 35884
rect 14710 35776 14904 35828
rect 14956 35776 14968 35828
rect 14710 35720 14968 35776
rect 14710 35668 14904 35720
rect 14956 35668 14968 35720
rect 14710 35658 14968 35668
rect 14710 35458 14721 35658
rect 14892 35612 14968 35658
rect 14892 35560 14904 35612
rect 14956 35560 14968 35612
rect 14892 35504 14968 35560
rect 14892 35458 14904 35504
rect 14710 35452 14904 35458
rect 14956 35452 14968 35504
rect 14710 35396 14968 35452
rect 14710 35344 14904 35396
rect 14956 35344 14968 35396
rect 14710 35288 14968 35344
rect 14710 35236 14904 35288
rect 14956 35236 14968 35288
rect 14710 35180 14968 35236
rect 14710 35128 14904 35180
rect 14956 35128 14968 35180
rect 14710 35072 14968 35128
rect 14710 35020 14904 35072
rect 14956 35020 14968 35072
rect 14710 34964 14968 35020
rect 14710 34912 14904 34964
rect 14956 34912 14968 34964
rect 14710 34856 14968 34912
rect 14710 34804 14904 34856
rect 14956 34804 14968 34856
rect 14710 34748 14968 34804
rect 14710 34696 14904 34748
rect 14956 34696 14968 34748
rect 14710 34640 14968 34696
rect 14710 34588 14904 34640
rect 14956 34588 14968 34640
rect 14710 34532 14968 34588
rect 14710 34480 14904 34532
rect 14956 34480 14968 34532
rect 14710 34458 14968 34480
rect 14710 34258 14721 34458
rect 14892 34424 14968 34458
rect 14892 34372 14904 34424
rect 14956 34372 14968 34424
rect 14892 34316 14968 34372
rect 14892 34264 14904 34316
rect 14956 34264 14968 34316
rect 14892 34258 14968 34264
rect 14710 34208 14968 34258
rect 14710 34156 14904 34208
rect 14956 34156 14968 34208
rect 14710 34100 14968 34156
rect 14710 34048 14904 34100
rect 14956 34048 14968 34100
rect 14710 33992 14968 34048
rect 14710 33940 14904 33992
rect 14956 33940 14968 33992
rect 14710 33884 14968 33940
rect 14710 33832 14904 33884
rect 14956 33832 14968 33884
rect 14710 33776 14968 33832
rect 14710 33724 14904 33776
rect 14956 33724 14968 33776
rect 14710 33668 14968 33724
rect 14710 33616 14904 33668
rect 14956 33616 14968 33668
rect 14710 33604 14968 33616
rect 14710 33258 14907 33604
rect 14710 33058 14721 33258
rect 14710 32058 14907 33058
rect 14710 31858 14721 32058
rect 14710 30858 14907 31858
rect 14710 30658 14721 30858
rect 14710 29658 14907 30658
rect 14710 29458 14721 29658
rect 14710 28586 14907 29458
rect 14710 28574 14968 28586
rect 14710 28522 14904 28574
rect 14956 28522 14968 28574
rect 14710 28466 14968 28522
rect 14710 28458 14904 28466
rect 14710 28258 14721 28458
rect 14892 28414 14904 28458
rect 14956 28414 14968 28466
rect 14892 28358 14968 28414
rect 14892 28306 14904 28358
rect 14956 28306 14968 28358
rect 14892 28258 14968 28306
rect 14710 28250 14968 28258
rect 14710 28198 14904 28250
rect 14956 28198 14968 28250
rect 14710 28142 14968 28198
rect 14710 28090 14904 28142
rect 14956 28090 14968 28142
rect 14710 28034 14968 28090
rect 14710 27982 14904 28034
rect 14956 27982 14968 28034
rect 14710 27926 14968 27982
rect 14710 27874 14904 27926
rect 14956 27874 14968 27926
rect 14710 27818 14968 27874
rect 14710 27766 14904 27818
rect 14956 27766 14968 27818
rect 14710 27710 14968 27766
rect 14710 27658 14904 27710
rect 14956 27658 14968 27710
rect 14710 27602 14968 27658
rect 14710 27550 14904 27602
rect 14956 27550 14968 27602
rect 14710 27494 14968 27550
rect 14710 27442 14904 27494
rect 14956 27442 14968 27494
rect 14710 27386 14968 27442
rect 14710 27334 14904 27386
rect 14956 27334 14968 27386
rect 14710 27278 14968 27334
rect 14710 27258 14904 27278
rect 14710 27058 14721 27258
rect 14892 27226 14904 27258
rect 14956 27226 14968 27278
rect 14892 27214 14968 27226
rect 14710 26058 14907 27058
rect 14710 25858 14721 26058
rect 14710 24858 14907 25858
rect 14710 24658 14721 24858
rect 14710 23658 14907 24658
rect 14710 23458 14721 23658
rect 14710 22458 14907 23458
rect 14710 21390 14721 22458
rect 14710 20390 14907 21390
rect 14710 20190 14721 20390
rect 14710 19190 14907 20190
rect 14710 18990 14721 19190
rect 14710 17990 14907 18990
rect 14710 17790 14721 17990
rect 14710 16790 14907 17790
rect 14710 16590 14721 16790
rect 14710 15590 14907 16590
rect 14710 15390 14721 15590
rect 14710 14390 14907 15390
rect 14710 14190 14721 14390
rect 14710 14186 14907 14190
rect 14710 14174 14968 14186
rect 14710 14122 14904 14174
rect 14956 14122 14968 14174
rect 14710 14066 14968 14122
rect 14710 14014 14904 14066
rect 14956 14014 14968 14066
rect 14710 13958 14968 14014
rect 14710 13906 14904 13958
rect 14956 13906 14968 13958
rect 14710 13850 14968 13906
rect 14710 13798 14904 13850
rect 14956 13798 14968 13850
rect 14710 13742 14968 13798
rect 14710 13690 14904 13742
rect 14956 13690 14968 13742
rect 14710 13634 14968 13690
rect 14710 13582 14904 13634
rect 14956 13582 14968 13634
rect 14710 13526 14968 13582
rect 14710 13474 14904 13526
rect 14956 13474 14968 13526
rect 14710 13418 14968 13474
rect 14710 13366 14904 13418
rect 14956 13366 14968 13418
rect 14710 13310 14968 13366
rect 14710 13258 14904 13310
rect 14956 13258 14968 13310
rect 14710 13202 14968 13258
rect 14710 13190 14904 13202
rect 14710 12990 14721 13190
rect 14892 13150 14904 13190
rect 14956 13150 14968 13202
rect 14892 13094 14968 13150
rect 14892 13042 14904 13094
rect 14956 13042 14968 13094
rect 14892 12990 14968 13042
rect 14710 12986 14968 12990
rect 14710 12934 14904 12986
rect 14956 12934 14968 12986
rect 14710 12878 14968 12934
rect 14710 12826 14904 12878
rect 14956 12826 14968 12878
rect 14710 12814 14968 12826
rect 14710 11990 14907 12814
rect 14710 11790 14721 11990
rect 14710 10996 14907 11790
rect 14710 10984 14968 10996
rect 14710 10932 14904 10984
rect 14956 10932 14968 10984
rect 14710 10876 14968 10932
rect 14710 10824 14904 10876
rect 14956 10824 14968 10876
rect 14710 10790 14968 10824
rect 14710 10590 14721 10790
rect 14892 10768 14968 10790
rect 14892 10716 14904 10768
rect 14956 10716 14968 10768
rect 14892 10660 14968 10716
rect 14892 10608 14904 10660
rect 14956 10608 14968 10660
rect 14892 10590 14968 10608
rect 14710 10552 14968 10590
rect 14710 10500 14904 10552
rect 14956 10500 14968 10552
rect 14710 10444 14968 10500
rect 14710 10392 14904 10444
rect 14956 10392 14968 10444
rect 14710 10336 14968 10392
rect 14710 10284 14904 10336
rect 14956 10284 14968 10336
rect 14710 10228 14968 10284
rect 14710 10176 14904 10228
rect 14956 10176 14968 10228
rect 14710 10120 14968 10176
rect 14710 10068 14904 10120
rect 14956 10068 14968 10120
rect 14710 10012 14968 10068
rect 14710 9960 14904 10012
rect 14956 9960 14968 10012
rect 14710 9904 14968 9960
rect 14710 9852 14904 9904
rect 14956 9852 14968 9904
rect 14710 9796 14968 9852
rect 14710 9744 14904 9796
rect 14956 9744 14968 9796
rect 14710 9688 14968 9744
rect 14710 9636 14904 9688
rect 14956 9636 14968 9688
rect 14710 9590 14968 9636
rect 14710 9390 14721 9590
rect 14892 9580 14968 9590
rect 14892 9528 14904 9580
rect 14956 9528 14968 9580
rect 14892 9472 14968 9528
rect 14892 9420 14904 9472
rect 14956 9420 14968 9472
rect 14892 9390 14968 9420
rect 14710 9364 14968 9390
rect 14710 9312 14904 9364
rect 14956 9312 14968 9364
rect 14710 9256 14968 9312
rect 14710 9204 14904 9256
rect 14956 9204 14968 9256
rect 14710 9148 14968 9204
rect 14710 9096 14904 9148
rect 14956 9096 14968 9148
rect 14710 9040 14968 9096
rect 14710 8988 14904 9040
rect 14956 8988 14968 9040
rect 14710 8932 14968 8988
rect 14710 8880 14904 8932
rect 14956 8880 14968 8932
rect 14710 8824 14968 8880
rect 14710 8772 14904 8824
rect 14956 8772 14968 8824
rect 14710 8716 14968 8772
rect 14710 8664 14904 8716
rect 14956 8664 14968 8716
rect 14710 8608 14968 8664
rect 14710 8556 14904 8608
rect 14956 8556 14968 8608
rect 14710 8500 14968 8556
rect 14710 8448 14904 8500
rect 14956 8448 14968 8500
rect 14710 8392 14968 8448
rect 14710 8390 14904 8392
rect 14710 8190 14721 8390
rect 14892 8340 14904 8390
rect 14956 8340 14968 8392
rect 14892 8284 14968 8340
rect 14892 8232 14904 8284
rect 14956 8232 14968 8284
rect 14892 8190 14968 8232
rect 14710 8176 14968 8190
rect 14710 8124 14904 8176
rect 14956 8124 14968 8176
rect 14710 8068 14968 8124
rect 14710 8016 14904 8068
rect 14956 8016 14968 8068
rect 14710 8004 14968 8016
rect 14710 7796 14907 8004
rect 14710 7784 14968 7796
rect 14710 7732 14904 7784
rect 14956 7732 14968 7784
rect 14710 7676 14968 7732
rect 14710 7624 14904 7676
rect 14956 7624 14968 7676
rect 14710 7568 14968 7624
rect 14710 7516 14904 7568
rect 14956 7516 14968 7568
rect 14710 7460 14968 7516
rect 14710 7408 14904 7460
rect 14956 7408 14968 7460
rect 14710 7352 14968 7408
rect 14710 7300 14904 7352
rect 14956 7300 14968 7352
rect 14710 7244 14968 7300
rect 14710 7192 14904 7244
rect 14956 7192 14968 7244
rect 14710 7190 14968 7192
rect 14710 6990 14721 7190
rect 14892 7136 14968 7190
rect 14892 7084 14904 7136
rect 14956 7084 14968 7136
rect 14892 7028 14968 7084
rect 14892 6990 14904 7028
rect 14710 6976 14904 6990
rect 14956 6976 14968 7028
rect 14710 6920 14968 6976
rect 14710 6868 14904 6920
rect 14956 6868 14968 6920
rect 14710 6812 14968 6868
rect 14710 6760 14904 6812
rect 14956 6760 14968 6812
rect 14710 6704 14968 6760
rect 14710 6652 14904 6704
rect 14956 6652 14968 6704
rect 14710 6596 14968 6652
rect 14710 6544 14904 6596
rect 14956 6544 14968 6596
rect 14710 6488 14968 6544
rect 14710 6436 14904 6488
rect 14956 6436 14968 6488
rect 14710 6380 14968 6436
rect 14710 6328 14904 6380
rect 14956 6328 14968 6380
rect 14710 6272 14968 6328
rect 14710 6220 14904 6272
rect 14956 6220 14968 6272
rect 14710 6164 14968 6220
rect 14710 6112 14904 6164
rect 14956 6112 14968 6164
rect 14710 6056 14968 6112
rect 14710 6004 14904 6056
rect 14956 6004 14968 6056
rect 14710 5990 14968 6004
rect 14710 5790 14721 5990
rect 14892 5948 14968 5990
rect 14892 5896 14904 5948
rect 14956 5896 14968 5948
rect 14892 5840 14968 5896
rect 14892 5790 14904 5840
rect 14710 5788 14904 5790
rect 14956 5788 14968 5840
rect 14710 5732 14968 5788
rect 14710 5680 14904 5732
rect 14956 5680 14968 5732
rect 14710 5624 14968 5680
rect 14710 5572 14904 5624
rect 14956 5572 14968 5624
rect 14710 5516 14968 5572
rect 14710 5464 14904 5516
rect 14956 5464 14968 5516
rect 14710 5408 14968 5464
rect 14710 5356 14904 5408
rect 14956 5356 14968 5408
rect 14710 5300 14968 5356
rect 14710 5248 14904 5300
rect 14956 5248 14968 5300
rect 14710 5192 14968 5248
rect 14710 5140 14904 5192
rect 14956 5140 14968 5192
rect 14710 5084 14968 5140
rect 14710 5032 14904 5084
rect 14956 5032 14968 5084
rect 14710 4976 14968 5032
rect 14710 4924 14904 4976
rect 14956 4924 14968 4976
rect 14710 4868 14968 4924
rect 14710 4816 14904 4868
rect 14956 4816 14968 4868
rect 14710 4804 14968 4816
rect 14710 4790 14907 4804
rect 14710 4590 14721 4790
rect 14892 4590 14968 4596
rect 14710 4584 14968 4590
rect 14710 4532 14904 4584
rect 14956 4532 14968 4584
rect 14710 4476 14968 4532
rect 14710 4424 14904 4476
rect 14956 4424 14968 4476
rect 14710 4368 14968 4424
rect 14710 4316 14904 4368
rect 14956 4316 14968 4368
rect 14710 4260 14968 4316
rect 14710 4208 14904 4260
rect 14956 4208 14968 4260
rect 14710 4152 14968 4208
rect 14710 4100 14904 4152
rect 14956 4100 14968 4152
rect 14710 4044 14968 4100
rect 14710 3992 14904 4044
rect 14956 3992 14968 4044
rect 14710 3936 14968 3992
rect 14710 3884 14904 3936
rect 14956 3884 14968 3936
rect 14710 3828 14968 3884
rect 14710 3776 14904 3828
rect 14956 3776 14968 3828
rect 14710 3720 14968 3776
rect 14710 3668 14904 3720
rect 14956 3668 14968 3720
rect 14710 3612 14968 3668
rect 14710 3590 14904 3612
rect 14710 3390 14721 3590
rect 14892 3560 14904 3590
rect 14956 3560 14968 3612
rect 14892 3504 14968 3560
rect 14892 3452 14904 3504
rect 14956 3452 14968 3504
rect 14892 3396 14968 3452
rect 14892 3390 14904 3396
rect 14710 3344 14904 3390
rect 14956 3344 14968 3396
rect 14710 3288 14968 3344
rect 14710 3236 14904 3288
rect 14956 3236 14968 3288
rect 14710 3180 14968 3236
rect 14710 3128 14904 3180
rect 14956 3128 14968 3180
rect 14710 3072 14968 3128
rect 14710 3020 14904 3072
rect 14956 3020 14968 3072
rect 14710 2964 14968 3020
rect 14710 2912 14904 2964
rect 14956 2912 14968 2964
rect 14710 2856 14968 2912
rect 14710 2804 14904 2856
rect 14956 2804 14968 2856
rect 14710 2748 14968 2804
rect 14710 2696 14904 2748
rect 14956 2696 14968 2748
rect 14710 2640 14968 2696
rect 14710 2588 14904 2640
rect 14956 2588 14968 2640
rect 14710 2532 14968 2588
rect 14710 2480 14904 2532
rect 14956 2480 14968 2532
rect 14710 2424 14968 2480
rect 14710 2390 14904 2424
rect 14710 2190 14721 2390
rect 14892 2372 14904 2390
rect 14956 2372 14968 2424
rect 14892 2316 14968 2372
rect 14892 2264 14904 2316
rect 14956 2264 14968 2316
rect 14892 2208 14968 2264
rect 14892 2190 14904 2208
rect 14710 2156 14904 2190
rect 14956 2156 14968 2208
rect 14710 2100 14968 2156
rect 14710 2048 14904 2100
rect 14956 2048 14968 2100
rect 14710 1992 14968 2048
rect 14710 1940 14904 1992
rect 14956 1940 14968 1992
rect 14710 1884 14968 1940
rect 14710 1832 14904 1884
rect 14956 1832 14968 1884
rect 14710 1776 14968 1832
rect 14710 1724 14904 1776
rect 14956 1724 14968 1776
rect 14710 1668 14968 1724
rect 14710 1616 14904 1668
rect 14956 1616 14968 1668
rect 14710 1604 14968 1616
rect 14710 1201 14907 1604
rect 14253 1190 14907 1201
<< via1 >>
rect 22 57207 74 57259
rect 22 57099 74 57151
rect 14904 57207 14956 57259
rect 22 56991 74 57043
rect 22 56883 74 56935
rect 22 56775 74 56827
rect 22 56667 74 56719
rect 22 56559 74 56611
rect 22 56451 74 56503
rect 22 56343 74 56395
rect 22 56235 74 56287
rect 22 56127 74 56179
rect 22 56019 74 56071
rect 22 54122 74 54174
rect 22 54014 74 54066
rect 22 53906 74 53958
rect 22 53798 74 53850
rect 22 53690 74 53742
rect 22 53582 74 53634
rect 22 53474 74 53526
rect 22 53366 74 53418
rect 22 53258 74 53310
rect 22 53150 74 53202
rect 375 57052 402 57104
rect 402 57052 427 57104
rect 483 57059 510 57104
rect 510 57059 535 57104
rect 591 57059 643 57104
rect 699 57059 751 57104
rect 807 57059 859 57104
rect 915 57059 967 57104
rect 1023 57059 1075 57104
rect 1131 57059 1183 57104
rect 1239 57059 1291 57104
rect 1347 57059 1399 57104
rect 1455 57059 1507 57104
rect 1563 57059 1615 57104
rect 1671 57059 1723 57104
rect 1779 57059 1831 57104
rect 1887 57059 1939 57104
rect 1995 57059 2047 57104
rect 2768 57059 2820 57104
rect 2876 57059 2928 57104
rect 2984 57059 3036 57104
rect 3092 57059 3144 57104
rect 3200 57059 3252 57104
rect 3308 57059 3360 57104
rect 3416 57059 3468 57104
rect 3524 57059 3576 57104
rect 3632 57059 3684 57104
rect 3740 57059 3792 57104
rect 3848 57059 3900 57104
rect 3956 57059 4008 57104
rect 4064 57059 4116 57104
rect 4172 57059 4224 57104
rect 4280 57059 4332 57104
rect 4388 57059 4440 57104
rect 4496 57059 4548 57104
rect 4604 57059 4656 57104
rect 4712 57059 4764 57104
rect 5138 57059 5190 57104
rect 5246 57059 5298 57104
rect 5354 57059 5406 57104
rect 5462 57059 5514 57104
rect 5570 57059 5622 57104
rect 5678 57059 5730 57104
rect 5786 57059 5838 57104
rect 5894 57059 5946 57104
rect 6002 57059 6054 57104
rect 6110 57059 6162 57104
rect 6218 57059 6270 57104
rect 6326 57059 6378 57104
rect 6434 57059 6486 57104
rect 6542 57059 6594 57104
rect 6650 57059 6702 57104
rect 6758 57059 6810 57104
rect 6866 57059 6918 57104
rect 6974 57059 7026 57104
rect 7082 57059 7134 57104
rect 7844 57059 7896 57104
rect 7952 57059 8004 57104
rect 8060 57059 8112 57104
rect 8168 57059 8220 57104
rect 8276 57059 8328 57104
rect 8384 57059 8436 57104
rect 8492 57059 8544 57104
rect 8600 57059 8652 57104
rect 8708 57059 8760 57104
rect 8816 57059 8868 57104
rect 8924 57059 8976 57104
rect 9032 57059 9084 57104
rect 9140 57059 9192 57104
rect 9248 57059 9300 57104
rect 9356 57059 9408 57104
rect 9464 57059 9516 57104
rect 9572 57059 9624 57104
rect 9680 57059 9732 57104
rect 9788 57059 9840 57104
rect 10214 57059 10266 57104
rect 10322 57059 10374 57104
rect 10430 57059 10482 57104
rect 10538 57059 10590 57104
rect 10646 57059 10698 57104
rect 10754 57059 10806 57104
rect 10862 57059 10914 57104
rect 10970 57059 11022 57104
rect 11078 57059 11130 57104
rect 11186 57059 11238 57104
rect 11294 57059 11346 57104
rect 11402 57059 11454 57104
rect 11510 57059 11562 57104
rect 11618 57059 11670 57104
rect 11726 57059 11778 57104
rect 11834 57059 11886 57104
rect 11942 57059 11994 57104
rect 12050 57059 12102 57104
rect 12158 57059 12210 57104
rect 12931 57059 12983 57104
rect 13039 57059 13091 57104
rect 13147 57059 13199 57104
rect 13255 57059 13307 57104
rect 13363 57059 13415 57104
rect 13471 57059 13523 57104
rect 13579 57059 13631 57104
rect 13687 57059 13739 57104
rect 13795 57059 13847 57104
rect 13903 57059 13955 57104
rect 14011 57059 14063 57104
rect 14119 57059 14171 57104
rect 14227 57059 14279 57104
rect 14335 57059 14387 57104
rect 14443 57059 14468 57104
rect 14468 57059 14495 57104
rect 483 57052 535 57059
rect 591 57052 643 57059
rect 699 57052 751 57059
rect 807 57052 859 57059
rect 915 57052 967 57059
rect 1023 57052 1075 57059
rect 1131 57052 1183 57059
rect 1239 57052 1291 57059
rect 1347 57052 1399 57059
rect 1455 57052 1507 57059
rect 1563 57052 1615 57059
rect 1671 57052 1723 57059
rect 1779 57052 1831 57059
rect 1887 57052 1939 57059
rect 1995 57052 2047 57059
rect 2768 57052 2820 57059
rect 2876 57052 2928 57059
rect 2984 57052 3036 57059
rect 3092 57052 3144 57059
rect 3200 57052 3252 57059
rect 3308 57052 3360 57059
rect 3416 57052 3468 57059
rect 3524 57052 3576 57059
rect 3632 57052 3684 57059
rect 3740 57052 3792 57059
rect 3848 57052 3900 57059
rect 3956 57052 4008 57059
rect 4064 57052 4116 57059
rect 4172 57052 4224 57059
rect 4280 57052 4332 57059
rect 4388 57052 4440 57059
rect 4496 57052 4548 57059
rect 4604 57052 4656 57059
rect 4712 57052 4764 57059
rect 5138 57052 5190 57059
rect 5246 57052 5298 57059
rect 5354 57052 5406 57059
rect 5462 57052 5514 57059
rect 5570 57052 5622 57059
rect 5678 57052 5730 57059
rect 5786 57052 5838 57059
rect 5894 57052 5946 57059
rect 6002 57052 6054 57059
rect 6110 57052 6162 57059
rect 6218 57052 6270 57059
rect 6326 57052 6378 57059
rect 6434 57052 6486 57059
rect 6542 57052 6594 57059
rect 6650 57052 6702 57059
rect 6758 57052 6810 57059
rect 6866 57052 6918 57059
rect 6974 57052 7026 57059
rect 7082 57052 7134 57059
rect 7844 57052 7896 57059
rect 7952 57052 8004 57059
rect 8060 57052 8112 57059
rect 8168 57052 8220 57059
rect 8276 57052 8328 57059
rect 8384 57052 8436 57059
rect 8492 57052 8544 57059
rect 8600 57052 8652 57059
rect 8708 57052 8760 57059
rect 8816 57052 8868 57059
rect 8924 57052 8976 57059
rect 9032 57052 9084 57059
rect 9140 57052 9192 57059
rect 9248 57052 9300 57059
rect 9356 57052 9408 57059
rect 9464 57052 9516 57059
rect 9572 57052 9624 57059
rect 9680 57052 9732 57059
rect 9788 57052 9840 57059
rect 10214 57052 10266 57059
rect 10322 57052 10374 57059
rect 10430 57052 10482 57059
rect 10538 57052 10590 57059
rect 10646 57052 10698 57059
rect 10754 57052 10806 57059
rect 10862 57052 10914 57059
rect 10970 57052 11022 57059
rect 11078 57052 11130 57059
rect 11186 57052 11238 57059
rect 11294 57052 11346 57059
rect 11402 57052 11454 57059
rect 11510 57052 11562 57059
rect 11618 57052 11670 57059
rect 11726 57052 11778 57059
rect 11834 57052 11886 57059
rect 11942 57052 11994 57059
rect 12050 57052 12102 57059
rect 12158 57052 12210 57059
rect 12931 57052 12983 57059
rect 13039 57052 13091 57059
rect 13147 57052 13199 57059
rect 13255 57052 13307 57059
rect 13363 57052 13415 57059
rect 13471 57052 13523 57059
rect 13579 57052 13631 57059
rect 13687 57052 13739 57059
rect 13795 57052 13847 57059
rect 13903 57052 13955 57059
rect 14011 57052 14063 57059
rect 14119 57052 14171 57059
rect 14227 57052 14279 57059
rect 14335 57052 14387 57059
rect 14443 57052 14495 57059
rect 14551 57052 14576 57104
rect 14576 57052 14603 57104
rect 2501 56734 2553 56741
rect 2609 56734 2661 56741
rect 2501 56689 2553 56734
rect 2609 56689 2661 56734
rect 369 56591 402 56643
rect 402 56591 421 56643
rect 493 56591 545 56643
rect 617 56591 669 56643
rect 741 56618 793 56643
rect 741 56591 760 56618
rect 760 56591 793 56618
rect 369 56467 402 56519
rect 402 56467 421 56519
rect 493 56467 545 56519
rect 617 56467 669 56519
rect 741 56467 760 56519
rect 760 56467 793 56519
rect 369 56343 402 56395
rect 402 56343 421 56395
rect 493 56343 545 56395
rect 617 56343 669 56395
rect 741 56343 760 56395
rect 760 56343 793 56395
rect 369 56219 402 56271
rect 402 56219 421 56271
rect 493 56219 545 56271
rect 617 56219 669 56271
rect 741 56219 760 56271
rect 760 56219 793 56271
rect 369 56095 402 56147
rect 402 56095 421 56147
rect 493 56095 545 56147
rect 617 56095 669 56147
rect 741 56095 760 56147
rect 760 56095 793 56147
rect 369 55971 402 56023
rect 402 55971 421 56023
rect 493 55971 545 56023
rect 617 55971 669 56023
rect 741 55971 760 56023
rect 760 55971 793 56023
rect 369 55847 402 55899
rect 402 55847 421 55899
rect 493 55847 545 55899
rect 617 55847 669 55899
rect 741 55847 760 55899
rect 760 55847 793 55899
rect 369 55723 402 55775
rect 402 55723 421 55775
rect 493 55723 545 55775
rect 617 55723 669 55775
rect 741 55723 760 55775
rect 760 55723 793 55775
rect 369 55599 402 55651
rect 402 55599 421 55651
rect 493 55599 545 55651
rect 617 55599 669 55651
rect 741 55599 760 55651
rect 760 55599 793 55651
rect 369 55475 402 55527
rect 402 55475 421 55527
rect 493 55475 545 55527
rect 617 55475 669 55527
rect 741 55475 760 55527
rect 760 55475 793 55527
rect 369 55351 402 55403
rect 402 55351 421 55403
rect 493 55351 545 55403
rect 617 55351 669 55403
rect 741 55351 760 55403
rect 760 55351 793 55403
rect 369 55227 402 55279
rect 402 55227 421 55279
rect 493 55227 545 55279
rect 617 55227 669 55279
rect 741 55227 760 55279
rect 760 55227 793 55279
rect 369 55103 402 55155
rect 402 55103 421 55155
rect 493 55103 545 55155
rect 617 55103 669 55155
rect 741 55103 760 55155
rect 760 55103 793 55155
rect 369 54979 402 55031
rect 402 54979 421 55031
rect 493 54979 545 55031
rect 617 54979 669 55031
rect 741 54979 760 55031
rect 760 54979 793 55031
rect 369 54855 402 54907
rect 402 54855 421 54907
rect 493 54855 545 54907
rect 617 54855 669 54907
rect 741 54855 760 54907
rect 760 54855 793 54907
rect 369 54731 402 54783
rect 402 54731 421 54783
rect 493 54731 545 54783
rect 617 54731 669 54783
rect 741 54731 760 54783
rect 760 54731 793 54783
rect 369 54607 402 54659
rect 402 54607 421 54659
rect 493 54607 545 54659
rect 617 54607 669 54659
rect 741 54607 760 54659
rect 760 54607 793 54659
rect 369 54483 402 54535
rect 402 54483 421 54535
rect 493 54483 545 54535
rect 617 54483 669 54535
rect 741 54483 760 54535
rect 760 54483 793 54535
rect 369 54359 402 54411
rect 402 54359 421 54411
rect 493 54359 545 54411
rect 617 54359 669 54411
rect 741 54359 760 54411
rect 760 54359 793 54411
rect 369 54235 402 54287
rect 402 54235 421 54287
rect 493 54235 545 54287
rect 617 54235 669 54287
rect 741 54235 760 54287
rect 760 54235 793 54287
rect 369 54111 402 54163
rect 402 54111 421 54163
rect 493 54111 545 54163
rect 617 54111 669 54163
rect 741 54111 760 54163
rect 760 54111 793 54163
rect 369 53987 402 54039
rect 402 53987 421 54039
rect 493 53987 545 54039
rect 617 53987 669 54039
rect 741 53987 760 54039
rect 760 53987 793 54039
rect 369 53863 402 53915
rect 402 53863 421 53915
rect 493 53863 545 53915
rect 617 53863 669 53915
rect 741 53863 760 53915
rect 760 53863 793 53915
rect 369 53739 402 53791
rect 402 53739 421 53791
rect 493 53739 545 53791
rect 617 53739 669 53791
rect 741 53739 760 53791
rect 760 53739 793 53791
rect 369 53615 402 53667
rect 402 53615 421 53667
rect 493 53615 545 53667
rect 617 53615 669 53667
rect 741 53615 793 53667
rect 4871 56688 4923 56693
rect 4979 56688 5031 56693
rect 2501 53576 2553 53621
rect 2609 53576 2661 53621
rect 2501 53569 2553 53576
rect 2609 53569 2661 53576
rect 3903 56618 3955 56643
rect 3903 56591 3910 56618
rect 3910 56591 3955 56618
rect 4027 56591 4079 56643
rect 4151 56618 4203 56643
rect 4151 56591 4196 56618
rect 4196 56591 4203 56618
rect 3903 56467 3910 56519
rect 3910 56467 3955 56519
rect 4027 56467 4079 56519
rect 4151 56467 4196 56519
rect 4196 56467 4203 56519
rect 3903 56343 3910 56395
rect 3910 56343 3955 56395
rect 4027 56343 4079 56395
rect 4151 56343 4196 56395
rect 4196 56343 4203 56395
rect 3903 56219 3910 56271
rect 3910 56219 3955 56271
rect 4027 56219 4079 56271
rect 4151 56219 4196 56271
rect 4196 56219 4203 56271
rect 3903 56095 3910 56147
rect 3910 56095 3955 56147
rect 4027 56095 4079 56147
rect 4151 56095 4196 56147
rect 4196 56095 4203 56147
rect 3903 55971 3910 56023
rect 3910 55971 3955 56023
rect 4027 55971 4079 56023
rect 4151 55971 4196 56023
rect 4196 55971 4203 56023
rect 3903 55847 3910 55899
rect 3910 55847 3955 55899
rect 4027 55847 4079 55899
rect 4151 55847 4196 55899
rect 4196 55847 4203 55899
rect 3903 55723 3910 55775
rect 3910 55723 3955 55775
rect 4027 55723 4079 55775
rect 4151 55723 4196 55775
rect 4196 55723 4203 55775
rect 3903 55599 3910 55651
rect 3910 55599 3955 55651
rect 4027 55599 4079 55651
rect 4151 55599 4196 55651
rect 4196 55599 4203 55651
rect 3903 55475 3910 55527
rect 3910 55475 3955 55527
rect 4027 55475 4079 55527
rect 4151 55475 4196 55527
rect 4196 55475 4203 55527
rect 3903 55351 3910 55403
rect 3910 55351 3955 55403
rect 4027 55351 4079 55403
rect 4151 55351 4196 55403
rect 4196 55351 4203 55403
rect 3903 55227 3910 55279
rect 3910 55227 3955 55279
rect 4027 55227 4079 55279
rect 4151 55227 4196 55279
rect 4196 55227 4203 55279
rect 3903 55103 3910 55155
rect 3910 55103 3955 55155
rect 4027 55103 4079 55155
rect 4151 55103 4196 55155
rect 4196 55103 4203 55155
rect 3903 54979 3910 55031
rect 3910 54979 3955 55031
rect 4027 54979 4079 55031
rect 4151 54979 4196 55031
rect 4196 54979 4203 55031
rect 3903 54855 3910 54907
rect 3910 54855 3955 54907
rect 4027 54855 4079 54907
rect 4151 54855 4196 54907
rect 4196 54855 4203 54907
rect 3903 54731 3910 54783
rect 3910 54731 3955 54783
rect 4027 54731 4079 54783
rect 4151 54731 4196 54783
rect 4196 54731 4203 54783
rect 3903 54607 3910 54659
rect 3910 54607 3955 54659
rect 4027 54607 4079 54659
rect 4151 54607 4196 54659
rect 4196 54607 4203 54659
rect 3903 54483 3910 54535
rect 3910 54483 3955 54535
rect 4027 54483 4079 54535
rect 4151 54483 4196 54535
rect 4196 54483 4203 54535
rect 3903 54359 3910 54411
rect 3910 54359 3955 54411
rect 4027 54359 4079 54411
rect 4151 54359 4196 54411
rect 4196 54359 4203 54411
rect 3903 54235 3910 54287
rect 3910 54235 3955 54287
rect 4027 54235 4079 54287
rect 4151 54235 4196 54287
rect 4196 54235 4203 54287
rect 3903 54111 3910 54163
rect 3910 54111 3955 54163
rect 4027 54111 4079 54163
rect 4151 54111 4196 54163
rect 4196 54111 4203 54163
rect 3903 53987 3910 54039
rect 3910 53987 3955 54039
rect 4027 53987 4079 54039
rect 4151 53987 4196 54039
rect 4196 53987 4203 54039
rect 3903 53863 3910 53915
rect 3910 53863 3955 53915
rect 4027 53863 4079 53915
rect 4151 53863 4196 53915
rect 4196 53863 4203 53915
rect 3903 53739 3910 53791
rect 3910 53739 3955 53791
rect 4027 53739 4079 53791
rect 4151 53739 4196 53791
rect 4196 53739 4203 53791
rect 3903 53615 3955 53667
rect 4027 53615 4079 53667
rect 4151 53615 4203 53667
rect 369 53491 402 53543
rect 402 53491 421 53543
rect 493 53491 545 53543
rect 617 53491 669 53543
rect 741 53491 793 53543
rect 4871 56641 4923 56688
rect 4979 56641 5031 56688
rect 4871 56533 4923 56585
rect 4979 56533 5031 56585
rect 4871 56425 4923 56477
rect 4979 56425 5031 56477
rect 4871 56317 4923 56369
rect 4979 56317 5031 56369
rect 4871 56209 4923 56261
rect 4979 56209 5031 56261
rect 4871 56101 4923 56153
rect 4979 56101 5031 56153
rect 4871 55993 4923 56045
rect 4979 55993 5031 56045
rect 4871 55885 4923 55937
rect 4979 55885 5031 55937
rect 4871 55777 4923 55829
rect 4979 55777 5031 55829
rect 4871 55669 4923 55721
rect 4979 55669 5031 55721
rect 4871 55561 4923 55613
rect 4979 55561 5031 55613
rect 4871 55453 4923 55505
rect 4979 55453 5031 55505
rect 4871 55345 4923 55397
rect 4979 55345 5031 55397
rect 4871 55237 4923 55289
rect 4979 55237 5031 55289
rect 4871 55129 4923 55181
rect 4979 55129 5031 55181
rect 4871 55021 4923 55073
rect 4979 55021 5031 55073
rect 4871 54913 4923 54965
rect 4979 54913 5031 54965
rect 4871 54805 4923 54857
rect 4979 54805 5031 54857
rect 4871 54697 4923 54749
rect 4979 54697 5031 54749
rect 4871 54589 4923 54641
rect 4979 54589 5031 54641
rect 4871 54481 4923 54533
rect 4979 54481 5031 54533
rect 4871 54373 4923 54425
rect 4979 54373 5031 54425
rect 4871 54265 4923 54317
rect 4979 54265 5031 54317
rect 4871 54157 4923 54209
rect 4979 54157 5031 54209
rect 4871 54049 4923 54101
rect 4979 54049 5031 54101
rect 4871 53941 4923 53993
rect 4979 53941 5031 53993
rect 4871 53833 4923 53885
rect 4979 53833 5031 53885
rect 4871 53725 4923 53777
rect 4979 53725 5031 53777
rect 4871 53622 4923 53669
rect 4979 53622 5031 53669
rect 9947 56688 9999 56693
rect 10055 56688 10107 56693
rect 4871 53617 4923 53622
rect 4979 53617 5031 53622
rect 3903 53491 3955 53543
rect 4027 53491 4079 53543
rect 4151 53491 4203 53543
rect 9947 56641 9999 56688
rect 10055 56641 10107 56688
rect 12317 56734 12369 56741
rect 12425 56734 12477 56741
rect 12317 56689 12369 56734
rect 12425 56689 12477 56734
rect 9947 56533 9999 56585
rect 10055 56533 10107 56585
rect 9947 56425 9999 56477
rect 10055 56425 10107 56477
rect 9947 56317 9999 56369
rect 10055 56317 10107 56369
rect 9947 56209 9999 56261
rect 10055 56209 10107 56261
rect 9947 56101 9999 56153
rect 10055 56101 10107 56153
rect 9947 55993 9999 56045
rect 10055 55993 10107 56045
rect 9947 55885 9999 55937
rect 10055 55885 10107 55937
rect 9947 55777 9999 55829
rect 10055 55777 10107 55829
rect 9947 55669 9999 55721
rect 10055 55669 10107 55721
rect 9947 55561 9999 55613
rect 10055 55561 10107 55613
rect 9947 55453 9999 55505
rect 10055 55453 10107 55505
rect 9947 55345 9999 55397
rect 10055 55345 10107 55397
rect 9947 55237 9999 55289
rect 10055 55237 10107 55289
rect 9947 55129 9999 55181
rect 10055 55129 10107 55181
rect 9947 55021 9999 55073
rect 10055 55021 10107 55073
rect 9947 54913 9999 54965
rect 10055 54913 10107 54965
rect 9947 54805 9999 54857
rect 10055 54805 10107 54857
rect 9947 54697 9999 54749
rect 10055 54697 10107 54749
rect 9947 54589 9999 54641
rect 10055 54589 10107 54641
rect 9947 54481 9999 54533
rect 10055 54481 10107 54533
rect 9947 54373 9999 54425
rect 10055 54373 10107 54425
rect 9947 54265 9999 54317
rect 10055 54265 10107 54317
rect 9947 54157 9999 54209
rect 10055 54157 10107 54209
rect 9947 54049 9999 54101
rect 10055 54049 10107 54101
rect 9947 53941 9999 53993
rect 10055 53941 10107 53993
rect 9947 53833 9999 53885
rect 10055 53833 10107 53885
rect 9947 53725 9999 53777
rect 10055 53725 10107 53777
rect 9947 53622 9999 53669
rect 10055 53622 10107 53669
rect 9947 53617 9999 53622
rect 10055 53617 10107 53622
rect 10775 56618 10827 56643
rect 10775 56591 10782 56618
rect 10782 56591 10827 56618
rect 10899 56591 10951 56643
rect 11023 56618 11075 56643
rect 11023 56591 11068 56618
rect 11068 56591 11075 56618
rect 10775 56467 10782 56519
rect 10782 56467 10827 56519
rect 10899 56467 10951 56519
rect 11023 56467 11068 56519
rect 11068 56467 11075 56519
rect 10775 56343 10782 56395
rect 10782 56343 10827 56395
rect 10899 56343 10951 56395
rect 11023 56343 11068 56395
rect 11068 56343 11075 56395
rect 10775 56219 10782 56271
rect 10782 56219 10827 56271
rect 10899 56219 10951 56271
rect 11023 56219 11068 56271
rect 11068 56219 11075 56271
rect 10775 56095 10782 56147
rect 10782 56095 10827 56147
rect 10899 56095 10951 56147
rect 11023 56095 11068 56147
rect 11068 56095 11075 56147
rect 10775 55971 10782 56023
rect 10782 55971 10827 56023
rect 10899 55971 10951 56023
rect 11023 55971 11068 56023
rect 11068 55971 11075 56023
rect 10775 55847 10782 55899
rect 10782 55847 10827 55899
rect 10899 55847 10951 55899
rect 11023 55847 11068 55899
rect 11068 55847 11075 55899
rect 10775 55723 10782 55775
rect 10782 55723 10827 55775
rect 10899 55723 10951 55775
rect 11023 55723 11068 55775
rect 11068 55723 11075 55775
rect 10775 55599 10782 55651
rect 10782 55599 10827 55651
rect 10899 55599 10951 55651
rect 11023 55599 11068 55651
rect 11068 55599 11075 55651
rect 10775 55475 10782 55527
rect 10782 55475 10827 55527
rect 10899 55475 10951 55527
rect 11023 55475 11068 55527
rect 11068 55475 11075 55527
rect 10775 55351 10782 55403
rect 10782 55351 10827 55403
rect 10899 55351 10951 55403
rect 11023 55351 11068 55403
rect 11068 55351 11075 55403
rect 10775 55227 10782 55279
rect 10782 55227 10827 55279
rect 10899 55227 10951 55279
rect 11023 55227 11068 55279
rect 11068 55227 11075 55279
rect 10775 55103 10782 55155
rect 10782 55103 10827 55155
rect 10899 55103 10951 55155
rect 11023 55103 11068 55155
rect 11068 55103 11075 55155
rect 10775 54979 10782 55031
rect 10782 54979 10827 55031
rect 10899 54979 10951 55031
rect 11023 54979 11068 55031
rect 11068 54979 11075 55031
rect 10775 54855 10782 54907
rect 10782 54855 10827 54907
rect 10899 54855 10951 54907
rect 11023 54855 11068 54907
rect 11068 54855 11075 54907
rect 10775 54731 10782 54783
rect 10782 54731 10827 54783
rect 10899 54731 10951 54783
rect 11023 54731 11068 54783
rect 11068 54731 11075 54783
rect 10775 54607 10782 54659
rect 10782 54607 10827 54659
rect 10899 54607 10951 54659
rect 11023 54607 11068 54659
rect 11068 54607 11075 54659
rect 10775 54483 10782 54535
rect 10782 54483 10827 54535
rect 10899 54483 10951 54535
rect 11023 54483 11068 54535
rect 11068 54483 11075 54535
rect 10775 54359 10782 54411
rect 10782 54359 10827 54411
rect 10899 54359 10951 54411
rect 11023 54359 11068 54411
rect 11068 54359 11075 54411
rect 10775 54235 10782 54287
rect 10782 54235 10827 54287
rect 10899 54235 10951 54287
rect 11023 54235 11068 54287
rect 11068 54235 11075 54287
rect 10775 54111 10782 54163
rect 10782 54111 10827 54163
rect 10899 54111 10951 54163
rect 11023 54111 11068 54163
rect 11068 54111 11075 54163
rect 10775 53987 10782 54039
rect 10782 53987 10827 54039
rect 10899 53987 10951 54039
rect 11023 53987 11068 54039
rect 11068 53987 11075 54039
rect 10775 53863 10782 53915
rect 10782 53863 10827 53915
rect 10899 53863 10951 53915
rect 11023 53863 11068 53915
rect 11068 53863 11075 53915
rect 10775 53739 10782 53791
rect 10782 53739 10827 53791
rect 10899 53739 10951 53791
rect 11023 53739 11068 53791
rect 11068 53739 11075 53791
rect 10775 53615 10827 53667
rect 10899 53615 10951 53667
rect 11023 53615 11075 53667
rect 12317 53576 12369 53621
rect 12425 53576 12477 53621
rect 12317 53569 12369 53576
rect 12425 53569 12477 53576
rect 14185 56618 14237 56643
rect 14185 56591 14218 56618
rect 14218 56591 14237 56618
rect 14309 56591 14361 56643
rect 14433 56591 14485 56643
rect 14557 56591 14576 56643
rect 14576 56591 14609 56643
rect 14185 56467 14218 56519
rect 14218 56467 14237 56519
rect 14309 56467 14361 56519
rect 14433 56467 14485 56519
rect 14557 56467 14576 56519
rect 14576 56467 14609 56519
rect 14185 56343 14218 56395
rect 14218 56343 14237 56395
rect 14309 56343 14361 56395
rect 14433 56343 14485 56395
rect 14557 56343 14576 56395
rect 14576 56343 14609 56395
rect 14185 56219 14218 56271
rect 14218 56219 14237 56271
rect 14309 56219 14361 56271
rect 14433 56219 14485 56271
rect 14557 56219 14576 56271
rect 14576 56219 14609 56271
rect 14185 56095 14218 56147
rect 14218 56095 14237 56147
rect 14309 56095 14361 56147
rect 14433 56095 14485 56147
rect 14557 56095 14576 56147
rect 14576 56095 14609 56147
rect 14185 55971 14218 56023
rect 14218 55971 14237 56023
rect 14309 55971 14361 56023
rect 14433 55971 14485 56023
rect 14557 55971 14576 56023
rect 14576 55971 14609 56023
rect 14185 55847 14218 55899
rect 14218 55847 14237 55899
rect 14309 55847 14361 55899
rect 14433 55847 14485 55899
rect 14557 55847 14576 55899
rect 14576 55847 14609 55899
rect 14185 55723 14218 55775
rect 14218 55723 14237 55775
rect 14309 55723 14361 55775
rect 14433 55723 14485 55775
rect 14557 55723 14576 55775
rect 14576 55723 14609 55775
rect 14185 55599 14218 55651
rect 14218 55599 14237 55651
rect 14309 55599 14361 55651
rect 14433 55599 14485 55651
rect 14557 55599 14576 55651
rect 14576 55599 14609 55651
rect 14185 55475 14218 55527
rect 14218 55475 14237 55527
rect 14309 55475 14361 55527
rect 14433 55475 14485 55527
rect 14557 55475 14576 55527
rect 14576 55475 14609 55527
rect 14185 55351 14218 55403
rect 14218 55351 14237 55403
rect 14309 55351 14361 55403
rect 14433 55351 14485 55403
rect 14557 55351 14576 55403
rect 14576 55351 14609 55403
rect 14185 55227 14218 55279
rect 14218 55227 14237 55279
rect 14309 55227 14361 55279
rect 14433 55227 14485 55279
rect 14557 55227 14576 55279
rect 14576 55227 14609 55279
rect 14185 55103 14218 55155
rect 14218 55103 14237 55155
rect 14309 55103 14361 55155
rect 14433 55103 14485 55155
rect 14557 55103 14576 55155
rect 14576 55103 14609 55155
rect 14185 54979 14218 55031
rect 14218 54979 14237 55031
rect 14309 54979 14361 55031
rect 14433 54979 14485 55031
rect 14557 54979 14576 55031
rect 14576 54979 14609 55031
rect 14185 54855 14218 54907
rect 14218 54855 14237 54907
rect 14309 54855 14361 54907
rect 14433 54855 14485 54907
rect 14557 54855 14576 54907
rect 14576 54855 14609 54907
rect 14185 54731 14218 54783
rect 14218 54731 14237 54783
rect 14309 54731 14361 54783
rect 14433 54731 14485 54783
rect 14557 54731 14576 54783
rect 14576 54731 14609 54783
rect 14185 54607 14218 54659
rect 14218 54607 14237 54659
rect 14309 54607 14361 54659
rect 14433 54607 14485 54659
rect 14557 54607 14576 54659
rect 14576 54607 14609 54659
rect 14185 54483 14218 54535
rect 14218 54483 14237 54535
rect 14309 54483 14361 54535
rect 14433 54483 14485 54535
rect 14557 54483 14576 54535
rect 14576 54483 14609 54535
rect 14185 54359 14218 54411
rect 14218 54359 14237 54411
rect 14309 54359 14361 54411
rect 14433 54359 14485 54411
rect 14557 54359 14576 54411
rect 14576 54359 14609 54411
rect 14185 54235 14218 54287
rect 14218 54235 14237 54287
rect 14309 54235 14361 54287
rect 14433 54235 14485 54287
rect 14557 54235 14576 54287
rect 14576 54235 14609 54287
rect 14185 54111 14218 54163
rect 14218 54111 14237 54163
rect 14309 54111 14361 54163
rect 14433 54111 14485 54163
rect 14557 54111 14576 54163
rect 14576 54111 14609 54163
rect 14185 53987 14218 54039
rect 14218 53987 14237 54039
rect 14309 53987 14361 54039
rect 14433 53987 14485 54039
rect 14557 53987 14576 54039
rect 14576 53987 14609 54039
rect 14185 53863 14218 53915
rect 14218 53863 14237 53915
rect 14309 53863 14361 53915
rect 14433 53863 14485 53915
rect 14557 53863 14576 53915
rect 14576 53863 14609 53915
rect 14185 53739 14218 53791
rect 14218 53739 14237 53791
rect 14309 53739 14361 53791
rect 14433 53739 14485 53791
rect 14557 53739 14576 53791
rect 14576 53739 14609 53791
rect 14185 53615 14237 53667
rect 14309 53615 14361 53667
rect 14433 53615 14485 53667
rect 14557 53615 14576 53667
rect 14576 53615 14609 53667
rect 10775 53491 10827 53543
rect 10899 53491 10951 53543
rect 11023 53491 11075 53543
rect 14185 53491 14237 53543
rect 14309 53491 14361 53543
rect 14433 53491 14485 53543
rect 14557 53491 14576 53543
rect 14576 53491 14609 53543
rect 869 53431 921 53483
rect 977 53431 1029 53483
rect 1085 53431 1137 53483
rect 1193 53431 1245 53483
rect 1301 53431 1353 53483
rect 1409 53431 1461 53483
rect 1517 53431 1569 53483
rect 1625 53431 1677 53483
rect 1733 53431 1785 53483
rect 1841 53431 1893 53483
rect 1949 53431 2001 53483
rect 2057 53431 2109 53483
rect 2763 53431 2815 53483
rect 2871 53431 2923 53483
rect 2979 53431 3031 53483
rect 3087 53431 3139 53483
rect 3195 53431 3247 53483
rect 3303 53431 3355 53483
rect 3411 53431 3463 53483
rect 3519 53431 3571 53483
rect 3627 53431 3679 53483
rect 3735 53431 3787 53483
rect 5138 53431 5190 53483
rect 5246 53431 5298 53483
rect 5354 53431 5406 53483
rect 5462 53431 5514 53483
rect 5570 53431 5622 53483
rect 5678 53431 5730 53483
rect 5786 53431 5838 53483
rect 5894 53431 5946 53483
rect 6002 53431 6054 53483
rect 6110 53431 6162 53483
rect 6218 53431 6270 53483
rect 6326 53431 6378 53483
rect 6434 53431 6486 53483
rect 6542 53431 6594 53483
rect 6650 53431 6702 53483
rect 6758 53431 6810 53483
rect 6866 53431 6918 53483
rect 6974 53431 7026 53483
rect 7082 53431 7134 53483
rect 7844 53431 7896 53483
rect 7952 53431 8004 53483
rect 8060 53431 8112 53483
rect 8168 53431 8220 53483
rect 8276 53431 8328 53483
rect 8384 53431 8436 53483
rect 8492 53431 8544 53483
rect 8600 53431 8652 53483
rect 8708 53431 8760 53483
rect 8816 53431 8868 53483
rect 8924 53431 8976 53483
rect 9032 53431 9084 53483
rect 9140 53431 9192 53483
rect 9248 53431 9300 53483
rect 9356 53431 9408 53483
rect 9464 53431 9516 53483
rect 9572 53431 9624 53483
rect 9680 53431 9732 53483
rect 9788 53431 9840 53483
rect 11191 53431 11243 53483
rect 11299 53431 11351 53483
rect 11407 53431 11459 53483
rect 11515 53431 11567 53483
rect 11623 53431 11675 53483
rect 11731 53431 11783 53483
rect 11839 53431 11891 53483
rect 11947 53431 11999 53483
rect 12055 53431 12107 53483
rect 12163 53431 12215 53483
rect 12869 53431 12921 53483
rect 12977 53431 13029 53483
rect 13085 53431 13137 53483
rect 13193 53431 13245 53483
rect 13301 53431 13353 53483
rect 13409 53431 13461 53483
rect 13517 53431 13569 53483
rect 13625 53431 13677 53483
rect 13733 53431 13785 53483
rect 13841 53431 13893 53483
rect 13949 53431 14001 53483
rect 14057 53431 14109 53483
rect 369 53367 402 53419
rect 402 53367 421 53419
rect 493 53367 545 53419
rect 617 53367 669 53419
rect 741 53367 793 53419
rect 869 53323 921 53375
rect 977 53323 1029 53375
rect 1085 53323 1137 53375
rect 1193 53323 1245 53375
rect 1301 53323 1353 53375
rect 1409 53323 1461 53375
rect 1517 53323 1569 53375
rect 1625 53323 1677 53375
rect 1733 53323 1785 53375
rect 1841 53323 1893 53375
rect 1949 53323 2001 53375
rect 2057 53323 2109 53375
rect 2763 53323 2815 53375
rect 2871 53323 2923 53375
rect 2979 53323 3031 53375
rect 3087 53323 3139 53375
rect 3195 53323 3247 53375
rect 3303 53323 3355 53375
rect 3411 53323 3463 53375
rect 3519 53323 3571 53375
rect 3627 53323 3679 53375
rect 3735 53323 3787 53375
rect 3903 53367 3955 53419
rect 4027 53367 4079 53419
rect 4151 53367 4203 53419
rect 5138 53323 5190 53375
rect 5246 53323 5298 53375
rect 5354 53323 5406 53375
rect 5462 53323 5514 53375
rect 5570 53323 5622 53375
rect 5678 53323 5730 53375
rect 5786 53323 5838 53375
rect 5894 53323 5946 53375
rect 6002 53323 6054 53375
rect 6110 53323 6162 53375
rect 6218 53323 6270 53375
rect 6326 53323 6378 53375
rect 6434 53323 6486 53375
rect 6542 53323 6594 53375
rect 6650 53323 6702 53375
rect 6758 53323 6810 53375
rect 6866 53323 6918 53375
rect 6974 53323 7026 53375
rect 7082 53323 7134 53375
rect 7844 53323 7896 53375
rect 7952 53323 8004 53375
rect 8060 53323 8112 53375
rect 8168 53323 8220 53375
rect 8276 53323 8328 53375
rect 8384 53323 8436 53375
rect 8492 53323 8544 53375
rect 8600 53323 8652 53375
rect 8708 53323 8760 53375
rect 8816 53323 8868 53375
rect 8924 53323 8976 53375
rect 9032 53323 9084 53375
rect 9140 53323 9192 53375
rect 9248 53323 9300 53375
rect 9356 53323 9408 53375
rect 9464 53323 9516 53375
rect 9572 53323 9624 53375
rect 9680 53323 9732 53375
rect 9788 53323 9840 53375
rect 10775 53367 10827 53419
rect 10899 53367 10951 53419
rect 11023 53367 11075 53419
rect 11191 53323 11243 53375
rect 11299 53323 11351 53375
rect 11407 53323 11459 53375
rect 11515 53323 11567 53375
rect 11623 53323 11675 53375
rect 11731 53323 11783 53375
rect 11839 53323 11891 53375
rect 11947 53323 11999 53375
rect 12055 53323 12107 53375
rect 12163 53323 12215 53375
rect 12869 53323 12921 53375
rect 12977 53323 13029 53375
rect 13085 53323 13137 53375
rect 13193 53323 13245 53375
rect 13301 53323 13353 53375
rect 13409 53323 13461 53375
rect 13517 53323 13569 53375
rect 13625 53323 13677 53375
rect 13733 53323 13785 53375
rect 13841 53323 13893 53375
rect 13949 53323 14001 53375
rect 14057 53323 14109 53375
rect 14185 53367 14237 53419
rect 14309 53367 14361 53419
rect 14433 53367 14485 53419
rect 14557 53367 14576 53419
rect 14576 53367 14609 53419
rect 369 53243 402 53295
rect 402 53243 421 53295
rect 493 53251 545 53295
rect 617 53251 669 53295
rect 741 53251 793 53295
rect 869 53251 921 53267
rect 977 53251 1029 53267
rect 1085 53251 1137 53267
rect 1193 53251 1245 53267
rect 1301 53251 1353 53267
rect 1409 53251 1461 53267
rect 1517 53251 1569 53267
rect 1625 53251 1677 53267
rect 1733 53251 1785 53267
rect 1841 53251 1893 53267
rect 1949 53251 2001 53267
rect 2057 53251 2109 53267
rect 2763 53251 2815 53267
rect 2871 53251 2923 53267
rect 2979 53251 3031 53267
rect 3087 53251 3139 53267
rect 3195 53251 3247 53267
rect 3303 53251 3355 53267
rect 3411 53251 3463 53267
rect 3519 53251 3571 53267
rect 3627 53251 3679 53267
rect 3735 53251 3787 53267
rect 3903 53251 3955 53295
rect 4027 53251 4079 53295
rect 4151 53251 4203 53295
rect 5138 53251 5190 53267
rect 5246 53251 5298 53267
rect 5354 53251 5406 53267
rect 5462 53251 5514 53267
rect 5570 53251 5622 53267
rect 5678 53251 5730 53267
rect 5786 53251 5838 53267
rect 5894 53251 5946 53267
rect 6002 53251 6054 53267
rect 6110 53251 6162 53267
rect 6218 53251 6270 53267
rect 6326 53251 6378 53267
rect 6434 53251 6486 53267
rect 6542 53251 6594 53267
rect 6650 53251 6702 53267
rect 6758 53251 6810 53267
rect 6866 53251 6918 53267
rect 6974 53251 7026 53267
rect 7082 53251 7134 53267
rect 7844 53251 7896 53267
rect 7952 53251 8004 53267
rect 8060 53251 8112 53267
rect 8168 53251 8220 53267
rect 8276 53251 8328 53267
rect 8384 53251 8436 53267
rect 8492 53251 8544 53267
rect 8600 53251 8652 53267
rect 8708 53251 8760 53267
rect 8816 53251 8868 53267
rect 8924 53251 8976 53267
rect 9032 53251 9084 53267
rect 9140 53251 9192 53267
rect 9248 53251 9300 53267
rect 9356 53251 9408 53267
rect 9464 53251 9516 53267
rect 9572 53251 9624 53267
rect 9680 53251 9732 53267
rect 9788 53251 9840 53267
rect 10775 53251 10827 53295
rect 10899 53251 10951 53295
rect 11023 53251 11075 53295
rect 11191 53251 11243 53267
rect 11299 53251 11351 53267
rect 11407 53251 11459 53267
rect 11515 53251 11567 53267
rect 11623 53251 11675 53267
rect 11731 53251 11783 53267
rect 11839 53251 11891 53267
rect 11947 53251 11999 53267
rect 12055 53251 12107 53267
rect 12163 53251 12215 53267
rect 12869 53251 12921 53267
rect 12977 53251 13029 53267
rect 13085 53251 13137 53267
rect 13193 53251 13245 53267
rect 13301 53251 13353 53267
rect 13409 53251 13461 53267
rect 13517 53251 13569 53267
rect 13625 53251 13677 53267
rect 13733 53251 13785 53267
rect 13841 53251 13893 53267
rect 13949 53251 14001 53267
rect 14057 53251 14109 53267
rect 14185 53251 14237 53295
rect 14309 53251 14361 53295
rect 14433 53251 14485 53295
rect 493 53243 510 53251
rect 510 53243 545 53251
rect 617 53243 669 53251
rect 741 53243 793 53251
rect 869 53215 921 53251
rect 977 53215 1029 53251
rect 1085 53215 1137 53251
rect 1193 53215 1245 53251
rect 1301 53215 1353 53251
rect 1409 53215 1461 53251
rect 1517 53215 1569 53251
rect 1625 53215 1677 53251
rect 1733 53215 1785 53251
rect 1841 53215 1893 53251
rect 1949 53215 2001 53251
rect 2057 53215 2109 53251
rect 2763 53215 2815 53251
rect 2871 53215 2923 53251
rect 2979 53215 3031 53251
rect 3087 53215 3139 53251
rect 3195 53215 3247 53251
rect 3303 53215 3355 53251
rect 3411 53215 3463 53251
rect 3519 53215 3571 53251
rect 3627 53215 3679 53251
rect 3735 53215 3787 53251
rect 3903 53243 3955 53251
rect 4027 53243 4079 53251
rect 4151 53243 4203 53251
rect 5138 53215 5190 53251
rect 5246 53215 5298 53251
rect 5354 53215 5406 53251
rect 5462 53215 5514 53251
rect 5570 53215 5622 53251
rect 5678 53215 5730 53251
rect 5786 53215 5838 53251
rect 5894 53215 5946 53251
rect 6002 53215 6054 53251
rect 6110 53215 6162 53251
rect 6218 53215 6270 53251
rect 6326 53215 6378 53251
rect 6434 53215 6486 53251
rect 6542 53215 6594 53251
rect 6650 53215 6702 53251
rect 6758 53215 6810 53251
rect 6866 53215 6918 53251
rect 6974 53215 7026 53251
rect 7082 53215 7134 53251
rect 7844 53215 7896 53251
rect 7952 53215 8004 53251
rect 8060 53215 8112 53251
rect 8168 53215 8220 53251
rect 8276 53215 8328 53251
rect 8384 53215 8436 53251
rect 8492 53215 8544 53251
rect 8600 53215 8652 53251
rect 8708 53215 8760 53251
rect 8816 53215 8868 53251
rect 8924 53215 8976 53251
rect 9032 53215 9084 53251
rect 9140 53215 9192 53251
rect 9248 53215 9300 53251
rect 9356 53215 9408 53251
rect 9464 53215 9516 53251
rect 9572 53215 9624 53251
rect 9680 53215 9732 53251
rect 9788 53215 9840 53251
rect 10775 53243 10827 53251
rect 10899 53243 10951 53251
rect 11023 53243 11075 53251
rect 11191 53215 11243 53251
rect 11299 53215 11351 53251
rect 11407 53215 11459 53251
rect 11515 53215 11567 53251
rect 11623 53215 11675 53251
rect 11731 53215 11783 53251
rect 11839 53215 11891 53251
rect 11947 53215 11999 53251
rect 12055 53215 12107 53251
rect 12163 53215 12215 53251
rect 12869 53215 12921 53251
rect 12977 53215 13029 53251
rect 13085 53215 13137 53251
rect 13193 53215 13245 53251
rect 13301 53215 13353 53251
rect 13409 53215 13461 53251
rect 13517 53215 13569 53251
rect 13625 53215 13677 53251
rect 13733 53215 13785 53251
rect 13841 53215 13893 53251
rect 13949 53215 14001 53251
rect 14057 53215 14109 53251
rect 14185 53243 14237 53251
rect 14309 53243 14361 53251
rect 14433 53243 14468 53251
rect 14468 53243 14485 53251
rect 14557 53243 14576 53295
rect 14576 53243 14609 53295
rect 14904 57099 14956 57151
rect 14904 56991 14956 57043
rect 14904 56883 14956 56935
rect 14904 56775 14956 56827
rect 14904 56667 14956 56719
rect 14904 56559 14956 56611
rect 14904 56451 14956 56503
rect 14904 56343 14956 56395
rect 14904 56235 14956 56287
rect 14904 56127 14956 56179
rect 14904 56019 14956 56071
rect 14904 54122 14956 54174
rect 14904 54014 14956 54066
rect 14904 53906 14956 53958
rect 14904 53798 14956 53850
rect 14904 53690 14956 53742
rect 14904 53582 14956 53634
rect 14904 53474 14956 53526
rect 14904 53366 14956 53418
rect 14904 53258 14956 53310
rect 22 53042 74 53094
rect 22 52934 74 52986
rect 22 52826 74 52878
rect 14904 53150 14956 53202
rect 14904 53042 14956 53094
rect 14904 52934 14956 52986
rect 14904 52826 14956 52878
rect 22 52522 74 52574
rect 22 52414 74 52466
rect 22 52306 74 52358
rect 22 52198 74 52250
rect 22 52090 74 52142
rect 22 51982 74 52034
rect 22 51874 74 51926
rect 22 51766 74 51818
rect 22 51658 74 51710
rect 22 51550 74 51602
rect 22 51442 74 51494
rect 22 51334 74 51386
rect 22 51226 74 51278
rect 22 49322 74 49374
rect 22 49214 74 49266
rect 22 49106 74 49158
rect 22 48998 74 49050
rect 22 48890 74 48942
rect 22 48782 74 48834
rect 22 48674 74 48726
rect 22 48566 74 48618
rect 22 48458 74 48510
rect 22 48350 74 48402
rect 22 48242 74 48294
rect 22 48134 74 48186
rect 22 48026 74 48078
rect 2590 52542 2642 52594
rect 2590 52434 2642 52486
rect 2590 52326 2642 52378
rect 2590 52218 2642 52270
rect 4871 52520 4923 52572
rect 4979 52520 5031 52572
rect 7247 52520 7299 52572
rect 7355 52520 7407 52572
rect 7463 52520 7515 52572
rect 7571 52520 7623 52572
rect 7679 52520 7731 52572
rect 9947 52520 9999 52572
rect 10055 52520 10107 52572
rect 4871 52412 4923 52464
rect 4979 52412 5031 52464
rect 7247 52412 7299 52464
rect 7355 52412 7407 52464
rect 7463 52412 7515 52464
rect 7571 52412 7623 52464
rect 7679 52412 7731 52464
rect 9947 52412 9999 52464
rect 10055 52412 10107 52464
rect 4871 52304 4923 52356
rect 4979 52304 5031 52356
rect 7247 52304 7299 52356
rect 7355 52304 7407 52356
rect 7463 52304 7515 52356
rect 7571 52304 7623 52356
rect 7679 52304 7731 52356
rect 9947 52304 9999 52356
rect 10055 52304 10107 52356
rect 12336 52542 12388 52594
rect 12336 52434 12388 52486
rect 12336 52326 12388 52378
rect 2590 52110 2642 52162
rect 2590 52002 2642 52054
rect 2590 51894 2642 51946
rect 2590 51786 2642 51838
rect 2590 51678 2642 51730
rect 2590 51570 2642 51622
rect 2590 51462 2642 51514
rect 2590 51354 2642 51406
rect 2590 51246 2642 51298
rect 2590 51138 2642 51190
rect 2590 51030 2642 51082
rect 2590 50922 2642 50974
rect 2590 50814 2642 50866
rect 2590 50706 2642 50758
rect 2590 50598 2642 50650
rect 2590 50490 2642 50542
rect 2590 50382 2642 50434
rect 2590 50274 2642 50326
rect 2590 50166 2642 50218
rect 2590 50058 2642 50110
rect 2590 49950 2642 50002
rect 2590 49842 2642 49894
rect 2590 49734 2642 49786
rect 2590 49626 2642 49678
rect 2590 49518 2642 49570
rect 2590 49410 2642 49462
rect 2590 49302 2642 49354
rect 2590 49194 2642 49246
rect 2590 49086 2642 49138
rect 2590 48978 2642 49030
rect 2590 48870 2642 48922
rect 2590 48762 2642 48814
rect 2590 48654 2642 48706
rect 2590 48546 2642 48598
rect 2590 48438 2642 48490
rect 2590 48330 2642 48382
rect 2590 48222 2642 48274
rect 2590 48114 2642 48166
rect 2590 48006 2642 48058
rect 3161 51983 3213 52009
rect 3269 51983 3321 52009
rect 3377 51983 3429 52009
rect 3485 51983 3537 52009
rect 3593 51983 3645 52009
rect 3701 51983 3753 52009
rect 3809 51983 3861 52009
rect 3917 51983 3969 52009
rect 4025 51983 4077 52009
rect 4133 51983 4185 52009
rect 4241 51983 4293 52009
rect 4349 51983 4401 52009
rect 4457 51983 4509 52009
rect 4565 51983 4617 52009
rect 4673 51983 4725 52009
rect 5138 51983 5190 52009
rect 5246 51983 5298 52009
rect 5354 51983 5406 52009
rect 5462 51983 5514 52009
rect 5570 51983 5622 52009
rect 5678 51983 5730 52009
rect 5786 51983 5838 52009
rect 5894 51983 5946 52009
rect 6002 51983 6054 52009
rect 6110 51983 6162 52009
rect 6218 51983 6270 52009
rect 6326 51983 6378 52009
rect 6434 51983 6486 52009
rect 6542 51983 6594 52009
rect 6650 51983 6702 52009
rect 6758 51983 6810 52009
rect 6866 51983 6918 52009
rect 6974 51983 7026 52009
rect 7082 51983 7134 52009
rect 7844 51983 7896 52009
rect 7952 51983 8004 52009
rect 8060 51983 8112 52009
rect 8168 51983 8220 52009
rect 8276 51983 8328 52009
rect 8384 51983 8436 52009
rect 8492 51983 8544 52009
rect 8600 51983 8652 52009
rect 8708 51983 8760 52009
rect 8816 51983 8868 52009
rect 8924 51983 8976 52009
rect 9032 51983 9084 52009
rect 9140 51983 9192 52009
rect 9248 51983 9300 52009
rect 9356 51983 9408 52009
rect 9464 51983 9516 52009
rect 9572 51983 9624 52009
rect 9680 51983 9732 52009
rect 9788 51983 9840 52009
rect 10253 51983 10305 52009
rect 10361 51983 10413 52009
rect 10469 51983 10521 52009
rect 10577 51983 10629 52009
rect 10685 51983 10737 52009
rect 10793 51983 10845 52009
rect 10901 51983 10953 52009
rect 11009 51983 11061 52009
rect 11117 51983 11169 52009
rect 11225 51983 11277 52009
rect 11333 51983 11385 52009
rect 11441 51983 11493 52009
rect 11549 51983 11601 52009
rect 11657 51983 11709 52009
rect 11765 51983 11817 52009
rect 3161 51957 3213 51983
rect 3269 51957 3321 51983
rect 3377 51957 3429 51983
rect 3485 51957 3537 51983
rect 3593 51957 3645 51983
rect 3701 51957 3753 51983
rect 3809 51957 3861 51983
rect 3917 51957 3969 51983
rect 4025 51957 4077 51983
rect 4133 51957 4185 51983
rect 4241 51957 4293 51983
rect 4349 51957 4401 51983
rect 4457 51957 4509 51983
rect 4565 51957 4617 51983
rect 4673 51957 4725 51983
rect 5138 51957 5190 51983
rect 5246 51957 5298 51983
rect 5354 51957 5406 51983
rect 5462 51957 5514 51983
rect 5570 51957 5622 51983
rect 5678 51957 5730 51983
rect 5786 51957 5838 51983
rect 5894 51957 5946 51983
rect 6002 51957 6054 51983
rect 6110 51957 6162 51983
rect 6218 51957 6270 51983
rect 6326 51957 6378 51983
rect 6434 51957 6486 51983
rect 6542 51957 6594 51983
rect 6650 51957 6702 51983
rect 6758 51957 6810 51983
rect 6866 51957 6918 51983
rect 6974 51957 7026 51983
rect 7082 51957 7134 51983
rect 7844 51957 7896 51983
rect 7952 51957 8004 51983
rect 8060 51957 8112 51983
rect 8168 51957 8220 51983
rect 8276 51957 8328 51983
rect 8384 51957 8436 51983
rect 8492 51957 8544 51983
rect 8600 51957 8652 51983
rect 8708 51957 8760 51983
rect 8816 51957 8868 51983
rect 8924 51957 8976 51983
rect 9032 51957 9084 51983
rect 9140 51957 9192 51983
rect 9248 51957 9300 51983
rect 9356 51957 9408 51983
rect 9464 51957 9516 51983
rect 9572 51957 9624 51983
rect 9680 51957 9732 51983
rect 9788 51957 9840 51983
rect 10253 51957 10305 51983
rect 10361 51957 10413 51983
rect 10469 51957 10521 51983
rect 10577 51957 10629 51983
rect 10685 51957 10737 51983
rect 10793 51957 10845 51983
rect 10901 51957 10953 51983
rect 11009 51957 11061 51983
rect 11117 51957 11169 51983
rect 11225 51957 11277 51983
rect 11333 51957 11385 51983
rect 11441 51957 11493 51983
rect 11549 51957 11601 51983
rect 11657 51957 11709 51983
rect 11765 51957 11817 51983
rect 3161 51900 3213 51901
rect 3161 51849 3162 51900
rect 3162 51849 3213 51900
rect 3269 51849 3321 51901
rect 3377 51875 3429 51901
rect 3485 51875 3537 51901
rect 3593 51875 3645 51901
rect 3701 51875 3753 51901
rect 3809 51875 3861 51901
rect 3917 51875 3969 51901
rect 4025 51875 4077 51901
rect 4133 51875 4185 51901
rect 4241 51875 4293 51901
rect 4349 51875 4401 51901
rect 4457 51875 4509 51901
rect 4565 51875 4617 51901
rect 4673 51875 4725 51901
rect 5138 51875 5190 51901
rect 5246 51875 5298 51901
rect 5354 51875 5406 51901
rect 5462 51875 5514 51901
rect 5570 51875 5622 51901
rect 5678 51875 5730 51901
rect 5786 51875 5838 51901
rect 5894 51875 5946 51901
rect 6002 51875 6054 51901
rect 6110 51875 6162 51901
rect 6218 51875 6270 51901
rect 6326 51875 6378 51901
rect 6434 51875 6486 51901
rect 6542 51875 6594 51901
rect 6650 51875 6702 51901
rect 6758 51875 6810 51901
rect 6866 51875 6918 51901
rect 6974 51875 7026 51901
rect 7082 51875 7134 51901
rect 7844 51875 7896 51901
rect 7952 51875 8004 51901
rect 8060 51875 8112 51901
rect 8168 51875 8220 51901
rect 8276 51875 8328 51901
rect 8384 51875 8436 51901
rect 8492 51875 8544 51901
rect 8600 51875 8652 51901
rect 8708 51875 8760 51901
rect 8816 51875 8868 51901
rect 8924 51875 8976 51901
rect 9032 51875 9084 51901
rect 9140 51875 9192 51901
rect 9248 51875 9300 51901
rect 9356 51875 9408 51901
rect 9464 51875 9516 51901
rect 9572 51875 9624 51901
rect 9680 51875 9732 51901
rect 9788 51875 9840 51901
rect 10253 51875 10305 51901
rect 10361 51875 10413 51901
rect 10469 51875 10521 51901
rect 10577 51875 10629 51901
rect 10685 51875 10737 51901
rect 10793 51875 10845 51901
rect 10901 51875 10953 51901
rect 11009 51875 11061 51901
rect 11117 51875 11169 51901
rect 11225 51875 11277 51901
rect 11333 51875 11385 51901
rect 11441 51875 11493 51901
rect 11549 51875 11601 51901
rect 3377 51849 3424 51875
rect 3424 51849 3429 51875
rect 3485 51849 3537 51875
rect 3593 51849 3645 51875
rect 3701 51849 3753 51875
rect 3809 51849 3861 51875
rect 3917 51849 3969 51875
rect 4025 51849 4077 51875
rect 4133 51849 4185 51875
rect 4241 51849 4293 51875
rect 4349 51849 4401 51875
rect 4457 51849 4509 51875
rect 4565 51849 4617 51875
rect 4673 51849 4725 51875
rect 5138 51849 5190 51875
rect 5246 51849 5298 51875
rect 5354 51849 5406 51875
rect 5462 51849 5514 51875
rect 5570 51849 5622 51875
rect 5678 51849 5730 51875
rect 5786 51849 5838 51875
rect 5894 51849 5946 51875
rect 6002 51849 6054 51875
rect 6110 51849 6162 51875
rect 6218 51849 6270 51875
rect 6326 51849 6378 51875
rect 6434 51849 6486 51875
rect 6542 51849 6594 51875
rect 6650 51849 6702 51875
rect 6758 51849 6810 51875
rect 6866 51849 6918 51875
rect 6974 51849 7026 51875
rect 7082 51849 7134 51875
rect 7844 51849 7896 51875
rect 7952 51849 8004 51875
rect 8060 51849 8112 51875
rect 8168 51849 8220 51875
rect 8276 51849 8328 51875
rect 8384 51849 8436 51875
rect 8492 51849 8544 51875
rect 8600 51849 8652 51875
rect 8708 51849 8760 51875
rect 8816 51849 8868 51875
rect 8924 51849 8976 51875
rect 9032 51849 9084 51875
rect 9140 51849 9192 51875
rect 9248 51849 9300 51875
rect 9356 51849 9408 51875
rect 9464 51849 9516 51875
rect 9572 51849 9624 51875
rect 9680 51849 9732 51875
rect 9788 51849 9840 51875
rect 10253 51849 10305 51875
rect 10361 51849 10413 51875
rect 10469 51849 10521 51875
rect 10577 51849 10629 51875
rect 10685 51849 10737 51875
rect 10793 51849 10845 51875
rect 10901 51849 10953 51875
rect 11009 51849 11061 51875
rect 11117 51849 11169 51875
rect 11225 51849 11277 51875
rect 11333 51849 11385 51875
rect 11441 51849 11493 51875
rect 11549 51849 11554 51875
rect 11554 51849 11601 51875
rect 11657 51849 11709 51901
rect 11765 51900 11817 51901
rect 11765 51849 11816 51900
rect 11816 51849 11817 51900
rect 4871 51580 4923 51619
rect 4979 51580 5031 51619
rect 7247 51580 7299 51619
rect 7355 51580 7407 51619
rect 7463 51580 7515 51619
rect 7571 51580 7623 51619
rect 7679 51580 7731 51619
rect 9947 51580 9999 51619
rect 10055 51580 10107 51619
rect 4871 51567 4923 51580
rect 4979 51567 5031 51580
rect 7247 51567 7299 51580
rect 7355 51567 7407 51580
rect 7463 51567 7515 51580
rect 7571 51567 7623 51580
rect 7679 51567 7731 51580
rect 9947 51567 9999 51580
rect 10055 51567 10107 51580
rect 4871 51498 4923 51511
rect 4979 51498 5031 51511
rect 7247 51498 7299 51511
rect 7355 51498 7407 51511
rect 7463 51498 7515 51511
rect 7571 51498 7623 51511
rect 7679 51498 7731 51511
rect 9947 51498 9999 51511
rect 10055 51498 10107 51511
rect 4871 51459 4923 51498
rect 4979 51459 5031 51498
rect 7247 51459 7299 51498
rect 7355 51459 7407 51498
rect 7463 51459 7515 51498
rect 7571 51459 7623 51498
rect 7679 51459 7731 51498
rect 9947 51459 9999 51498
rect 10055 51459 10107 51498
rect 3161 51154 3162 51206
rect 3162 51154 3213 51206
rect 3269 51154 3321 51206
rect 3377 51203 3424 51206
rect 3424 51203 3429 51206
rect 3485 51203 3537 51206
rect 3593 51203 3645 51206
rect 3701 51203 3753 51206
rect 3809 51203 3861 51206
rect 3917 51203 3969 51206
rect 4025 51203 4077 51206
rect 4133 51203 4185 51206
rect 4241 51203 4293 51206
rect 4349 51203 4401 51206
rect 4457 51203 4509 51206
rect 4565 51203 4617 51206
rect 4673 51203 4725 51206
rect 5138 51203 5190 51206
rect 5246 51203 5298 51206
rect 5354 51203 5406 51206
rect 5462 51203 5514 51206
rect 5570 51203 5622 51206
rect 5678 51203 5730 51206
rect 5786 51203 5838 51206
rect 5894 51203 5946 51206
rect 6002 51203 6054 51206
rect 6110 51203 6162 51206
rect 6218 51203 6270 51206
rect 6326 51203 6378 51206
rect 6434 51203 6486 51206
rect 6542 51203 6594 51206
rect 6650 51203 6702 51206
rect 6758 51203 6810 51206
rect 6866 51203 6918 51206
rect 6974 51203 7026 51206
rect 7082 51203 7134 51206
rect 7844 51203 7896 51206
rect 7952 51203 8004 51206
rect 8060 51203 8112 51206
rect 8168 51203 8220 51206
rect 8276 51203 8328 51206
rect 8384 51203 8436 51206
rect 8492 51203 8544 51206
rect 8600 51203 8652 51206
rect 8708 51203 8760 51206
rect 8816 51203 8868 51206
rect 8924 51203 8976 51206
rect 9032 51203 9084 51206
rect 9140 51203 9192 51206
rect 9248 51203 9300 51206
rect 9356 51203 9408 51206
rect 9464 51203 9516 51206
rect 9572 51203 9624 51206
rect 9680 51203 9732 51206
rect 9788 51203 9840 51206
rect 10253 51203 10305 51206
rect 10361 51203 10413 51206
rect 10469 51203 10521 51206
rect 10577 51203 10629 51206
rect 10685 51203 10737 51206
rect 10793 51203 10845 51206
rect 10901 51203 10953 51206
rect 11009 51203 11061 51206
rect 11117 51203 11169 51206
rect 11225 51203 11277 51206
rect 11333 51203 11385 51206
rect 11441 51203 11493 51206
rect 11549 51203 11554 51206
rect 11554 51203 11601 51206
rect 3377 51154 3429 51203
rect 3485 51154 3537 51203
rect 3593 51154 3645 51203
rect 3701 51154 3753 51203
rect 3809 51154 3861 51203
rect 3917 51154 3969 51203
rect 4025 51154 4077 51203
rect 4133 51154 4185 51203
rect 4241 51154 4293 51203
rect 4349 51154 4401 51203
rect 4457 51154 4509 51203
rect 4565 51154 4617 51203
rect 4673 51154 4725 51203
rect 5138 51154 5190 51203
rect 5246 51154 5298 51203
rect 5354 51154 5406 51203
rect 5462 51154 5514 51203
rect 5570 51154 5622 51203
rect 5678 51154 5730 51203
rect 5786 51154 5838 51203
rect 5894 51154 5946 51203
rect 6002 51154 6054 51203
rect 6110 51154 6162 51203
rect 6218 51154 6270 51203
rect 6326 51154 6378 51203
rect 6434 51154 6486 51203
rect 6542 51154 6594 51203
rect 6650 51154 6702 51203
rect 6758 51154 6810 51203
rect 6866 51154 6918 51203
rect 6974 51154 7026 51203
rect 7082 51154 7134 51203
rect 7844 51154 7896 51203
rect 7952 51154 8004 51203
rect 8060 51154 8112 51203
rect 8168 51154 8220 51203
rect 8276 51154 8328 51203
rect 8384 51154 8436 51203
rect 8492 51154 8544 51203
rect 8600 51154 8652 51203
rect 8708 51154 8760 51203
rect 8816 51154 8868 51203
rect 8924 51154 8976 51203
rect 9032 51154 9084 51203
rect 9140 51154 9192 51203
rect 9248 51154 9300 51203
rect 9356 51154 9408 51203
rect 9464 51154 9516 51203
rect 9572 51154 9624 51203
rect 9680 51154 9732 51203
rect 9788 51154 9840 51203
rect 10253 51154 10305 51203
rect 10361 51154 10413 51203
rect 10469 51154 10521 51203
rect 10577 51154 10629 51203
rect 10685 51154 10737 51203
rect 10793 51154 10845 51203
rect 10901 51154 10953 51203
rect 11009 51154 11061 51203
rect 11117 51154 11169 51203
rect 11225 51154 11277 51203
rect 11333 51154 11385 51203
rect 11441 51154 11493 51203
rect 11549 51154 11601 51203
rect 11657 51154 11709 51206
rect 11765 51154 11816 51206
rect 11816 51154 11817 51206
rect 3161 51046 3162 51098
rect 3162 51046 3213 51098
rect 3269 51046 3321 51098
rect 3377 51095 3429 51098
rect 3485 51095 3537 51098
rect 3593 51095 3645 51098
rect 3701 51095 3753 51098
rect 3809 51095 3861 51098
rect 3917 51095 3969 51098
rect 4025 51095 4077 51098
rect 4133 51095 4185 51098
rect 4241 51095 4293 51098
rect 4349 51095 4401 51098
rect 4457 51095 4509 51098
rect 4565 51095 4617 51098
rect 4673 51095 4725 51098
rect 5138 51095 5190 51098
rect 5246 51095 5298 51098
rect 5354 51095 5406 51098
rect 5462 51095 5514 51098
rect 5570 51095 5622 51098
rect 5678 51095 5730 51098
rect 5786 51095 5838 51098
rect 5894 51095 5946 51098
rect 6002 51095 6054 51098
rect 6110 51095 6162 51098
rect 6218 51095 6270 51098
rect 6326 51095 6378 51098
rect 6434 51095 6486 51098
rect 6542 51095 6594 51098
rect 6650 51095 6702 51098
rect 6758 51095 6810 51098
rect 6866 51095 6918 51098
rect 6974 51095 7026 51098
rect 7082 51095 7134 51098
rect 7844 51095 7896 51098
rect 7952 51095 8004 51098
rect 8060 51095 8112 51098
rect 8168 51095 8220 51098
rect 8276 51095 8328 51098
rect 8384 51095 8436 51098
rect 8492 51095 8544 51098
rect 8600 51095 8652 51098
rect 8708 51095 8760 51098
rect 8816 51095 8868 51098
rect 8924 51095 8976 51098
rect 9032 51095 9084 51098
rect 9140 51095 9192 51098
rect 9248 51095 9300 51098
rect 9356 51095 9408 51098
rect 9464 51095 9516 51098
rect 9572 51095 9624 51098
rect 9680 51095 9732 51098
rect 9788 51095 9840 51098
rect 10253 51095 10305 51098
rect 10361 51095 10413 51098
rect 10469 51095 10521 51098
rect 10577 51095 10629 51098
rect 10685 51095 10737 51098
rect 10793 51095 10845 51098
rect 10901 51095 10953 51098
rect 11009 51095 11061 51098
rect 11117 51095 11169 51098
rect 11225 51095 11277 51098
rect 11333 51095 11385 51098
rect 11441 51095 11493 51098
rect 11549 51095 11601 51098
rect 3377 51049 3429 51095
rect 3485 51049 3537 51095
rect 3593 51049 3645 51095
rect 3701 51049 3753 51095
rect 3809 51049 3861 51095
rect 3917 51049 3969 51095
rect 4025 51049 4077 51095
rect 4133 51049 4185 51095
rect 4241 51049 4293 51095
rect 4349 51049 4401 51095
rect 4457 51049 4509 51095
rect 4565 51049 4617 51095
rect 4673 51049 4725 51095
rect 5138 51049 5190 51095
rect 5246 51049 5298 51095
rect 5354 51049 5406 51095
rect 5462 51049 5514 51095
rect 5570 51049 5622 51095
rect 5678 51049 5730 51095
rect 5786 51049 5838 51095
rect 5894 51049 5946 51095
rect 6002 51049 6054 51095
rect 6110 51049 6162 51095
rect 6218 51049 6270 51095
rect 6326 51049 6378 51095
rect 6434 51049 6486 51095
rect 6542 51049 6594 51095
rect 6650 51049 6702 51095
rect 6758 51049 6810 51095
rect 6866 51049 6918 51095
rect 6974 51049 7026 51095
rect 7082 51049 7134 51095
rect 7844 51049 7896 51095
rect 7952 51049 8004 51095
rect 8060 51049 8112 51095
rect 8168 51049 8220 51095
rect 8276 51049 8328 51095
rect 8384 51049 8436 51095
rect 8492 51049 8544 51095
rect 8600 51049 8652 51095
rect 8708 51049 8760 51095
rect 8816 51049 8868 51095
rect 8924 51049 8976 51095
rect 9032 51049 9084 51095
rect 9140 51049 9192 51095
rect 9248 51049 9300 51095
rect 9356 51049 9408 51095
rect 9464 51049 9516 51095
rect 9572 51049 9624 51095
rect 9680 51049 9732 51095
rect 9788 51049 9840 51095
rect 10253 51049 10305 51095
rect 10361 51049 10413 51095
rect 10469 51049 10521 51095
rect 10577 51049 10629 51095
rect 10685 51049 10737 51095
rect 10793 51049 10845 51095
rect 10901 51049 10953 51095
rect 11009 51049 11061 51095
rect 11117 51049 11169 51095
rect 11225 51049 11277 51095
rect 11333 51049 11385 51095
rect 11441 51049 11493 51095
rect 11549 51049 11601 51095
rect 3377 51046 3429 51049
rect 3485 51046 3537 51049
rect 3593 51046 3645 51049
rect 3701 51046 3753 51049
rect 3809 51046 3861 51049
rect 3917 51046 3969 51049
rect 4025 51046 4077 51049
rect 4133 51046 4185 51049
rect 4241 51046 4293 51049
rect 4349 51046 4401 51049
rect 4457 51046 4509 51049
rect 4565 51046 4617 51049
rect 4673 51046 4725 51049
rect 5138 51046 5190 51049
rect 5246 51046 5298 51049
rect 5354 51046 5406 51049
rect 5462 51046 5514 51049
rect 5570 51046 5622 51049
rect 5678 51046 5730 51049
rect 5786 51046 5838 51049
rect 5894 51046 5946 51049
rect 6002 51046 6054 51049
rect 6110 51046 6162 51049
rect 6218 51046 6270 51049
rect 6326 51046 6378 51049
rect 6434 51046 6486 51049
rect 6542 51046 6594 51049
rect 6650 51046 6702 51049
rect 6758 51046 6810 51049
rect 6866 51046 6918 51049
rect 6974 51046 7026 51049
rect 7082 51046 7134 51049
rect 7844 51046 7896 51049
rect 7952 51046 8004 51049
rect 8060 51046 8112 51049
rect 8168 51046 8220 51049
rect 8276 51046 8328 51049
rect 8384 51046 8436 51049
rect 8492 51046 8544 51049
rect 8600 51046 8652 51049
rect 8708 51046 8760 51049
rect 8816 51046 8868 51049
rect 8924 51046 8976 51049
rect 9032 51046 9084 51049
rect 9140 51046 9192 51049
rect 9248 51046 9300 51049
rect 9356 51046 9408 51049
rect 9464 51046 9516 51049
rect 9572 51046 9624 51049
rect 9680 51046 9732 51049
rect 9788 51046 9840 51049
rect 10253 51046 10305 51049
rect 10361 51046 10413 51049
rect 10469 51046 10521 51049
rect 10577 51046 10629 51049
rect 10685 51046 10737 51049
rect 10793 51046 10845 51049
rect 10901 51046 10953 51049
rect 11009 51046 11061 51049
rect 11117 51046 11169 51049
rect 11225 51046 11277 51049
rect 11333 51046 11385 51049
rect 11441 51046 11493 51049
rect 11549 51046 11601 51049
rect 11657 51046 11709 51098
rect 11765 51046 11816 51098
rect 11816 51046 11817 51098
rect 3161 50938 3162 50990
rect 3162 50938 3213 50990
rect 3269 50938 3321 50990
rect 3377 50941 3429 50990
rect 3485 50941 3537 50990
rect 3593 50941 3645 50990
rect 3701 50941 3753 50990
rect 3809 50941 3861 50990
rect 3917 50941 3969 50990
rect 4025 50941 4077 50990
rect 4133 50941 4185 50990
rect 4241 50941 4293 50990
rect 4349 50941 4401 50990
rect 4457 50941 4509 50990
rect 4565 50941 4617 50990
rect 4673 50941 4725 50990
rect 5138 50941 5190 50990
rect 5246 50941 5298 50990
rect 5354 50941 5406 50990
rect 5462 50941 5514 50990
rect 5570 50941 5622 50990
rect 5678 50941 5730 50990
rect 5786 50941 5838 50990
rect 5894 50941 5946 50990
rect 6002 50941 6054 50990
rect 6110 50941 6162 50990
rect 6218 50941 6270 50990
rect 6326 50941 6378 50990
rect 6434 50941 6486 50990
rect 6542 50941 6594 50990
rect 6650 50941 6702 50990
rect 6758 50941 6810 50990
rect 6866 50941 6918 50990
rect 6974 50941 7026 50990
rect 7082 50941 7134 50990
rect 7844 50941 7896 50990
rect 7952 50941 8004 50990
rect 8060 50941 8112 50990
rect 8168 50941 8220 50990
rect 8276 50941 8328 50990
rect 8384 50941 8436 50990
rect 8492 50941 8544 50990
rect 8600 50941 8652 50990
rect 8708 50941 8760 50990
rect 8816 50941 8868 50990
rect 8924 50941 8976 50990
rect 9032 50941 9084 50990
rect 9140 50941 9192 50990
rect 9248 50941 9300 50990
rect 9356 50941 9408 50990
rect 9464 50941 9516 50990
rect 9572 50941 9624 50990
rect 9680 50941 9732 50990
rect 9788 50941 9840 50990
rect 10253 50941 10305 50990
rect 10361 50941 10413 50990
rect 10469 50941 10521 50990
rect 10577 50941 10629 50990
rect 10685 50941 10737 50990
rect 10793 50941 10845 50990
rect 10901 50941 10953 50990
rect 11009 50941 11061 50990
rect 11117 50941 11169 50990
rect 11225 50941 11277 50990
rect 11333 50941 11385 50990
rect 11441 50941 11493 50990
rect 11549 50941 11601 50990
rect 3377 50938 3424 50941
rect 3424 50938 3429 50941
rect 3485 50938 3537 50941
rect 3593 50938 3645 50941
rect 3701 50938 3753 50941
rect 3809 50938 3861 50941
rect 3917 50938 3969 50941
rect 4025 50938 4077 50941
rect 4133 50938 4185 50941
rect 4241 50938 4293 50941
rect 4349 50938 4401 50941
rect 4457 50938 4509 50941
rect 4565 50938 4617 50941
rect 4673 50938 4725 50941
rect 5138 50938 5190 50941
rect 5246 50938 5298 50941
rect 5354 50938 5406 50941
rect 5462 50938 5514 50941
rect 5570 50938 5622 50941
rect 5678 50938 5730 50941
rect 5786 50938 5838 50941
rect 5894 50938 5946 50941
rect 6002 50938 6054 50941
rect 6110 50938 6162 50941
rect 6218 50938 6270 50941
rect 6326 50938 6378 50941
rect 6434 50938 6486 50941
rect 6542 50938 6594 50941
rect 6650 50938 6702 50941
rect 6758 50938 6810 50941
rect 6866 50938 6918 50941
rect 6974 50938 7026 50941
rect 7082 50938 7134 50941
rect 7844 50938 7896 50941
rect 7952 50938 8004 50941
rect 8060 50938 8112 50941
rect 8168 50938 8220 50941
rect 8276 50938 8328 50941
rect 8384 50938 8436 50941
rect 8492 50938 8544 50941
rect 8600 50938 8652 50941
rect 8708 50938 8760 50941
rect 8816 50938 8868 50941
rect 8924 50938 8976 50941
rect 9032 50938 9084 50941
rect 9140 50938 9192 50941
rect 9248 50938 9300 50941
rect 9356 50938 9408 50941
rect 9464 50938 9516 50941
rect 9572 50938 9624 50941
rect 9680 50938 9732 50941
rect 9788 50938 9840 50941
rect 10253 50938 10305 50941
rect 10361 50938 10413 50941
rect 10469 50938 10521 50941
rect 10577 50938 10629 50941
rect 10685 50938 10737 50941
rect 10793 50938 10845 50941
rect 10901 50938 10953 50941
rect 11009 50938 11061 50941
rect 11117 50938 11169 50941
rect 11225 50938 11277 50941
rect 11333 50938 11385 50941
rect 11441 50938 11493 50941
rect 11549 50938 11554 50941
rect 11554 50938 11601 50941
rect 11657 50938 11709 50990
rect 11765 50938 11816 50990
rect 11816 50938 11817 50990
rect 4871 50646 4923 50685
rect 4979 50646 5031 50685
rect 7247 50646 7299 50685
rect 7355 50646 7407 50685
rect 7463 50646 7515 50685
rect 7571 50646 7623 50685
rect 7679 50646 7731 50685
rect 9947 50646 9999 50685
rect 10055 50646 10107 50685
rect 4871 50633 4923 50646
rect 4979 50633 5031 50646
rect 7247 50633 7299 50646
rect 7355 50633 7407 50646
rect 7463 50633 7515 50646
rect 7571 50633 7623 50646
rect 7679 50633 7731 50646
rect 9947 50633 9999 50646
rect 10055 50633 10107 50646
rect 4871 50564 4923 50577
rect 4979 50564 5031 50577
rect 7247 50564 7299 50577
rect 7355 50564 7407 50577
rect 7463 50564 7515 50577
rect 7571 50564 7623 50577
rect 7679 50564 7731 50577
rect 9947 50564 9999 50577
rect 10055 50564 10107 50577
rect 4871 50525 4923 50564
rect 4979 50525 5031 50564
rect 7247 50525 7299 50564
rect 7355 50525 7407 50564
rect 7463 50525 7515 50564
rect 7571 50525 7623 50564
rect 7679 50525 7731 50564
rect 9947 50525 9999 50564
rect 10055 50525 10107 50564
rect 3161 50220 3162 50272
rect 3162 50220 3213 50272
rect 3269 50220 3321 50272
rect 3377 50269 3424 50272
rect 3424 50269 3429 50272
rect 3485 50269 3537 50272
rect 3593 50269 3645 50272
rect 3701 50269 3753 50272
rect 3809 50269 3861 50272
rect 3917 50269 3969 50272
rect 4025 50269 4077 50272
rect 4133 50269 4185 50272
rect 4241 50269 4293 50272
rect 4349 50269 4401 50272
rect 4457 50269 4509 50272
rect 4565 50269 4617 50272
rect 4673 50269 4725 50272
rect 5138 50269 5190 50272
rect 5246 50269 5298 50272
rect 5354 50269 5406 50272
rect 5462 50269 5514 50272
rect 5570 50269 5622 50272
rect 5678 50269 5730 50272
rect 5786 50269 5838 50272
rect 5894 50269 5946 50272
rect 6002 50269 6054 50272
rect 6110 50269 6162 50272
rect 6218 50269 6270 50272
rect 6326 50269 6378 50272
rect 6434 50269 6486 50272
rect 6542 50269 6594 50272
rect 6650 50269 6702 50272
rect 6758 50269 6810 50272
rect 6866 50269 6918 50272
rect 6974 50269 7026 50272
rect 7082 50269 7134 50272
rect 7844 50269 7896 50272
rect 7952 50269 8004 50272
rect 8060 50269 8112 50272
rect 8168 50269 8220 50272
rect 8276 50269 8328 50272
rect 8384 50269 8436 50272
rect 8492 50269 8544 50272
rect 8600 50269 8652 50272
rect 8708 50269 8760 50272
rect 8816 50269 8868 50272
rect 8924 50269 8976 50272
rect 9032 50269 9084 50272
rect 9140 50269 9192 50272
rect 9248 50269 9300 50272
rect 9356 50269 9408 50272
rect 9464 50269 9516 50272
rect 9572 50269 9624 50272
rect 9680 50269 9732 50272
rect 9788 50269 9840 50272
rect 10253 50269 10305 50272
rect 10361 50269 10413 50272
rect 10469 50269 10521 50272
rect 10577 50269 10629 50272
rect 10685 50269 10737 50272
rect 10793 50269 10845 50272
rect 10901 50269 10953 50272
rect 11009 50269 11061 50272
rect 11117 50269 11169 50272
rect 11225 50269 11277 50272
rect 11333 50269 11385 50272
rect 11441 50269 11493 50272
rect 11549 50269 11554 50272
rect 11554 50269 11601 50272
rect 3377 50220 3429 50269
rect 3485 50220 3537 50269
rect 3593 50220 3645 50269
rect 3701 50220 3753 50269
rect 3809 50220 3861 50269
rect 3917 50220 3969 50269
rect 4025 50220 4077 50269
rect 4133 50220 4185 50269
rect 4241 50220 4293 50269
rect 4349 50220 4401 50269
rect 4457 50220 4509 50269
rect 4565 50220 4617 50269
rect 4673 50220 4725 50269
rect 5138 50220 5190 50269
rect 5246 50220 5298 50269
rect 5354 50220 5406 50269
rect 5462 50220 5514 50269
rect 5570 50220 5622 50269
rect 5678 50220 5730 50269
rect 5786 50220 5838 50269
rect 5894 50220 5946 50269
rect 6002 50220 6054 50269
rect 6110 50220 6162 50269
rect 6218 50220 6270 50269
rect 6326 50220 6378 50269
rect 6434 50220 6486 50269
rect 6542 50220 6594 50269
rect 6650 50220 6702 50269
rect 6758 50220 6810 50269
rect 6866 50220 6918 50269
rect 6974 50220 7026 50269
rect 7082 50220 7134 50269
rect 7844 50220 7896 50269
rect 7952 50220 8004 50269
rect 8060 50220 8112 50269
rect 8168 50220 8220 50269
rect 8276 50220 8328 50269
rect 8384 50220 8436 50269
rect 8492 50220 8544 50269
rect 8600 50220 8652 50269
rect 8708 50220 8760 50269
rect 8816 50220 8868 50269
rect 8924 50220 8976 50269
rect 9032 50220 9084 50269
rect 9140 50220 9192 50269
rect 9248 50220 9300 50269
rect 9356 50220 9408 50269
rect 9464 50220 9516 50269
rect 9572 50220 9624 50269
rect 9680 50220 9732 50269
rect 9788 50220 9840 50269
rect 10253 50220 10305 50269
rect 10361 50220 10413 50269
rect 10469 50220 10521 50269
rect 10577 50220 10629 50269
rect 10685 50220 10737 50269
rect 10793 50220 10845 50269
rect 10901 50220 10953 50269
rect 11009 50220 11061 50269
rect 11117 50220 11169 50269
rect 11225 50220 11277 50269
rect 11333 50220 11385 50269
rect 11441 50220 11493 50269
rect 11549 50220 11601 50269
rect 11657 50220 11709 50272
rect 11765 50220 11816 50272
rect 11816 50220 11817 50272
rect 3161 50112 3162 50164
rect 3162 50112 3213 50164
rect 3269 50112 3321 50164
rect 3377 50161 3429 50164
rect 3485 50161 3537 50164
rect 3593 50161 3645 50164
rect 3701 50161 3753 50164
rect 3809 50161 3861 50164
rect 3917 50161 3969 50164
rect 4025 50161 4077 50164
rect 4133 50161 4185 50164
rect 4241 50161 4293 50164
rect 4349 50161 4401 50164
rect 4457 50161 4509 50164
rect 4565 50161 4617 50164
rect 4673 50161 4725 50164
rect 5138 50161 5190 50164
rect 5246 50161 5298 50164
rect 5354 50161 5406 50164
rect 5462 50161 5514 50164
rect 5570 50161 5622 50164
rect 5678 50161 5730 50164
rect 5786 50161 5838 50164
rect 5894 50161 5946 50164
rect 6002 50161 6054 50164
rect 6110 50161 6162 50164
rect 6218 50161 6270 50164
rect 6326 50161 6378 50164
rect 6434 50161 6486 50164
rect 6542 50161 6594 50164
rect 6650 50161 6702 50164
rect 6758 50161 6810 50164
rect 6866 50161 6918 50164
rect 6974 50161 7026 50164
rect 7082 50161 7134 50164
rect 7844 50161 7896 50164
rect 7952 50161 8004 50164
rect 8060 50161 8112 50164
rect 8168 50161 8220 50164
rect 8276 50161 8328 50164
rect 8384 50161 8436 50164
rect 8492 50161 8544 50164
rect 8600 50161 8652 50164
rect 8708 50161 8760 50164
rect 8816 50161 8868 50164
rect 8924 50161 8976 50164
rect 9032 50161 9084 50164
rect 9140 50161 9192 50164
rect 9248 50161 9300 50164
rect 9356 50161 9408 50164
rect 9464 50161 9516 50164
rect 9572 50161 9624 50164
rect 9680 50161 9732 50164
rect 9788 50161 9840 50164
rect 10253 50161 10305 50164
rect 10361 50161 10413 50164
rect 10469 50161 10521 50164
rect 10577 50161 10629 50164
rect 10685 50161 10737 50164
rect 10793 50161 10845 50164
rect 10901 50161 10953 50164
rect 11009 50161 11061 50164
rect 11117 50161 11169 50164
rect 11225 50161 11277 50164
rect 11333 50161 11385 50164
rect 11441 50161 11493 50164
rect 11549 50161 11601 50164
rect 3377 50115 3429 50161
rect 3485 50115 3537 50161
rect 3593 50115 3645 50161
rect 3701 50115 3753 50161
rect 3809 50115 3861 50161
rect 3917 50115 3969 50161
rect 4025 50115 4077 50161
rect 4133 50115 4185 50161
rect 4241 50115 4293 50161
rect 4349 50115 4401 50161
rect 4457 50115 4509 50161
rect 4565 50115 4617 50161
rect 4673 50115 4725 50161
rect 5138 50115 5190 50161
rect 5246 50115 5298 50161
rect 5354 50115 5406 50161
rect 5462 50115 5514 50161
rect 5570 50115 5622 50161
rect 5678 50115 5730 50161
rect 5786 50115 5838 50161
rect 5894 50115 5946 50161
rect 6002 50115 6054 50161
rect 6110 50115 6162 50161
rect 6218 50115 6270 50161
rect 6326 50115 6378 50161
rect 6434 50115 6486 50161
rect 6542 50115 6594 50161
rect 6650 50115 6702 50161
rect 6758 50115 6810 50161
rect 6866 50115 6918 50161
rect 6974 50115 7026 50161
rect 7082 50115 7134 50161
rect 7844 50115 7896 50161
rect 7952 50115 8004 50161
rect 8060 50115 8112 50161
rect 8168 50115 8220 50161
rect 8276 50115 8328 50161
rect 8384 50115 8436 50161
rect 8492 50115 8544 50161
rect 8600 50115 8652 50161
rect 8708 50115 8760 50161
rect 8816 50115 8868 50161
rect 8924 50115 8976 50161
rect 9032 50115 9084 50161
rect 9140 50115 9192 50161
rect 9248 50115 9300 50161
rect 9356 50115 9408 50161
rect 9464 50115 9516 50161
rect 9572 50115 9624 50161
rect 9680 50115 9732 50161
rect 9788 50115 9840 50161
rect 10253 50115 10305 50161
rect 10361 50115 10413 50161
rect 10469 50115 10521 50161
rect 10577 50115 10629 50161
rect 10685 50115 10737 50161
rect 10793 50115 10845 50161
rect 10901 50115 10953 50161
rect 11009 50115 11061 50161
rect 11117 50115 11169 50161
rect 11225 50115 11277 50161
rect 11333 50115 11385 50161
rect 11441 50115 11493 50161
rect 11549 50115 11601 50161
rect 3377 50112 3429 50115
rect 3485 50112 3537 50115
rect 3593 50112 3645 50115
rect 3701 50112 3753 50115
rect 3809 50112 3861 50115
rect 3917 50112 3969 50115
rect 4025 50112 4077 50115
rect 4133 50112 4185 50115
rect 4241 50112 4293 50115
rect 4349 50112 4401 50115
rect 4457 50112 4509 50115
rect 4565 50112 4617 50115
rect 4673 50112 4725 50115
rect 5138 50112 5190 50115
rect 5246 50112 5298 50115
rect 5354 50112 5406 50115
rect 5462 50112 5514 50115
rect 5570 50112 5622 50115
rect 5678 50112 5730 50115
rect 5786 50112 5838 50115
rect 5894 50112 5946 50115
rect 6002 50112 6054 50115
rect 6110 50112 6162 50115
rect 6218 50112 6270 50115
rect 6326 50112 6378 50115
rect 6434 50112 6486 50115
rect 6542 50112 6594 50115
rect 6650 50112 6702 50115
rect 6758 50112 6810 50115
rect 6866 50112 6918 50115
rect 6974 50112 7026 50115
rect 7082 50112 7134 50115
rect 7844 50112 7896 50115
rect 7952 50112 8004 50115
rect 8060 50112 8112 50115
rect 8168 50112 8220 50115
rect 8276 50112 8328 50115
rect 8384 50112 8436 50115
rect 8492 50112 8544 50115
rect 8600 50112 8652 50115
rect 8708 50112 8760 50115
rect 8816 50112 8868 50115
rect 8924 50112 8976 50115
rect 9032 50112 9084 50115
rect 9140 50112 9192 50115
rect 9248 50112 9300 50115
rect 9356 50112 9408 50115
rect 9464 50112 9516 50115
rect 9572 50112 9624 50115
rect 9680 50112 9732 50115
rect 9788 50112 9840 50115
rect 10253 50112 10305 50115
rect 10361 50112 10413 50115
rect 10469 50112 10521 50115
rect 10577 50112 10629 50115
rect 10685 50112 10737 50115
rect 10793 50112 10845 50115
rect 10901 50112 10953 50115
rect 11009 50112 11061 50115
rect 11117 50112 11169 50115
rect 11225 50112 11277 50115
rect 11333 50112 11385 50115
rect 11441 50112 11493 50115
rect 11549 50112 11601 50115
rect 11657 50112 11709 50164
rect 11765 50112 11816 50164
rect 11816 50112 11817 50164
rect 3161 50004 3162 50056
rect 3162 50004 3213 50056
rect 3269 50004 3321 50056
rect 3377 50007 3429 50056
rect 3485 50007 3537 50056
rect 3593 50007 3645 50056
rect 3701 50007 3753 50056
rect 3809 50007 3861 50056
rect 3917 50007 3969 50056
rect 4025 50007 4077 50056
rect 4133 50007 4185 50056
rect 4241 50007 4293 50056
rect 4349 50007 4401 50056
rect 4457 50007 4509 50056
rect 4565 50007 4617 50056
rect 4673 50007 4725 50056
rect 5138 50007 5190 50056
rect 5246 50007 5298 50056
rect 5354 50007 5406 50056
rect 5462 50007 5514 50056
rect 5570 50007 5622 50056
rect 5678 50007 5730 50056
rect 5786 50007 5838 50056
rect 5894 50007 5946 50056
rect 6002 50007 6054 50056
rect 6110 50007 6162 50056
rect 6218 50007 6270 50056
rect 6326 50007 6378 50056
rect 6434 50007 6486 50056
rect 6542 50007 6594 50056
rect 6650 50007 6702 50056
rect 6758 50007 6810 50056
rect 6866 50007 6918 50056
rect 6974 50007 7026 50056
rect 7082 50007 7134 50056
rect 7844 50007 7896 50056
rect 7952 50007 8004 50056
rect 8060 50007 8112 50056
rect 8168 50007 8220 50056
rect 8276 50007 8328 50056
rect 8384 50007 8436 50056
rect 8492 50007 8544 50056
rect 8600 50007 8652 50056
rect 8708 50007 8760 50056
rect 8816 50007 8868 50056
rect 8924 50007 8976 50056
rect 9032 50007 9084 50056
rect 9140 50007 9192 50056
rect 9248 50007 9300 50056
rect 9356 50007 9408 50056
rect 9464 50007 9516 50056
rect 9572 50007 9624 50056
rect 9680 50007 9732 50056
rect 9788 50007 9840 50056
rect 10253 50007 10305 50056
rect 10361 50007 10413 50056
rect 10469 50007 10521 50056
rect 10577 50007 10629 50056
rect 10685 50007 10737 50056
rect 10793 50007 10845 50056
rect 10901 50007 10953 50056
rect 11009 50007 11061 50056
rect 11117 50007 11169 50056
rect 11225 50007 11277 50056
rect 11333 50007 11385 50056
rect 11441 50007 11493 50056
rect 11549 50007 11601 50056
rect 3377 50004 3424 50007
rect 3424 50004 3429 50007
rect 3485 50004 3537 50007
rect 3593 50004 3645 50007
rect 3701 50004 3753 50007
rect 3809 50004 3861 50007
rect 3917 50004 3969 50007
rect 4025 50004 4077 50007
rect 4133 50004 4185 50007
rect 4241 50004 4293 50007
rect 4349 50004 4401 50007
rect 4457 50004 4509 50007
rect 4565 50004 4617 50007
rect 4673 50004 4725 50007
rect 5138 50004 5190 50007
rect 5246 50004 5298 50007
rect 5354 50004 5406 50007
rect 5462 50004 5514 50007
rect 5570 50004 5622 50007
rect 5678 50004 5730 50007
rect 5786 50004 5838 50007
rect 5894 50004 5946 50007
rect 6002 50004 6054 50007
rect 6110 50004 6162 50007
rect 6218 50004 6270 50007
rect 6326 50004 6378 50007
rect 6434 50004 6486 50007
rect 6542 50004 6594 50007
rect 6650 50004 6702 50007
rect 6758 50004 6810 50007
rect 6866 50004 6918 50007
rect 6974 50004 7026 50007
rect 7082 50004 7134 50007
rect 7844 50004 7896 50007
rect 7952 50004 8004 50007
rect 8060 50004 8112 50007
rect 8168 50004 8220 50007
rect 8276 50004 8328 50007
rect 8384 50004 8436 50007
rect 8492 50004 8544 50007
rect 8600 50004 8652 50007
rect 8708 50004 8760 50007
rect 8816 50004 8868 50007
rect 8924 50004 8976 50007
rect 9032 50004 9084 50007
rect 9140 50004 9192 50007
rect 9248 50004 9300 50007
rect 9356 50004 9408 50007
rect 9464 50004 9516 50007
rect 9572 50004 9624 50007
rect 9680 50004 9732 50007
rect 9788 50004 9840 50007
rect 10253 50004 10305 50007
rect 10361 50004 10413 50007
rect 10469 50004 10521 50007
rect 10577 50004 10629 50007
rect 10685 50004 10737 50007
rect 10793 50004 10845 50007
rect 10901 50004 10953 50007
rect 11009 50004 11061 50007
rect 11117 50004 11169 50007
rect 11225 50004 11277 50007
rect 11333 50004 11385 50007
rect 11441 50004 11493 50007
rect 11549 50004 11554 50007
rect 11554 50004 11601 50007
rect 11657 50004 11709 50056
rect 11765 50004 11816 50056
rect 11816 50004 11817 50056
rect 4871 49712 4923 49751
rect 4979 49712 5031 49751
rect 7247 49712 7299 49751
rect 7355 49712 7407 49751
rect 7463 49712 7515 49751
rect 7571 49712 7623 49751
rect 7679 49712 7731 49751
rect 9947 49712 9999 49751
rect 10055 49712 10107 49751
rect 4871 49699 4923 49712
rect 4979 49699 5031 49712
rect 7247 49699 7299 49712
rect 7355 49699 7407 49712
rect 7463 49699 7515 49712
rect 7571 49699 7623 49712
rect 7679 49699 7731 49712
rect 9947 49699 9999 49712
rect 10055 49699 10107 49712
rect 4871 49630 4923 49643
rect 4979 49630 5031 49643
rect 7247 49630 7299 49643
rect 7355 49630 7407 49643
rect 7463 49630 7515 49643
rect 7571 49630 7623 49643
rect 7679 49630 7731 49643
rect 9947 49630 9999 49643
rect 10055 49630 10107 49643
rect 4871 49591 4923 49630
rect 4979 49591 5031 49630
rect 7247 49591 7299 49630
rect 7355 49591 7407 49630
rect 7463 49591 7515 49630
rect 7571 49591 7623 49630
rect 7679 49591 7731 49630
rect 9947 49591 9999 49630
rect 10055 49591 10107 49630
rect 3161 49286 3162 49338
rect 3162 49286 3213 49338
rect 3269 49286 3321 49338
rect 3377 49335 3424 49338
rect 3424 49335 3429 49338
rect 3485 49335 3537 49338
rect 3593 49335 3645 49338
rect 3701 49335 3753 49338
rect 3809 49335 3861 49338
rect 3917 49335 3969 49338
rect 4025 49335 4077 49338
rect 4133 49335 4185 49338
rect 4241 49335 4293 49338
rect 4349 49335 4401 49338
rect 4457 49335 4509 49338
rect 4565 49335 4617 49338
rect 4673 49335 4725 49338
rect 5138 49335 5190 49338
rect 5246 49335 5298 49338
rect 5354 49335 5406 49338
rect 5462 49335 5514 49338
rect 5570 49335 5622 49338
rect 5678 49335 5730 49338
rect 5786 49335 5838 49338
rect 5894 49335 5946 49338
rect 6002 49335 6054 49338
rect 6110 49335 6162 49338
rect 6218 49335 6270 49338
rect 6326 49335 6378 49338
rect 6434 49335 6486 49338
rect 6542 49335 6594 49338
rect 6650 49335 6702 49338
rect 6758 49335 6810 49338
rect 6866 49335 6918 49338
rect 6974 49335 7026 49338
rect 7082 49335 7134 49338
rect 7844 49335 7896 49338
rect 7952 49335 8004 49338
rect 8060 49335 8112 49338
rect 8168 49335 8220 49338
rect 8276 49335 8328 49338
rect 8384 49335 8436 49338
rect 8492 49335 8544 49338
rect 8600 49335 8652 49338
rect 8708 49335 8760 49338
rect 8816 49335 8868 49338
rect 8924 49335 8976 49338
rect 9032 49335 9084 49338
rect 9140 49335 9192 49338
rect 9248 49335 9300 49338
rect 9356 49335 9408 49338
rect 9464 49335 9516 49338
rect 9572 49335 9624 49338
rect 9680 49335 9732 49338
rect 9788 49335 9840 49338
rect 10253 49335 10305 49338
rect 10361 49335 10413 49338
rect 10469 49335 10521 49338
rect 10577 49335 10629 49338
rect 10685 49335 10737 49338
rect 10793 49335 10845 49338
rect 10901 49335 10953 49338
rect 11009 49335 11061 49338
rect 11117 49335 11169 49338
rect 11225 49335 11277 49338
rect 11333 49335 11385 49338
rect 11441 49335 11493 49338
rect 11549 49335 11554 49338
rect 11554 49335 11601 49338
rect 3377 49286 3429 49335
rect 3485 49286 3537 49335
rect 3593 49286 3645 49335
rect 3701 49286 3753 49335
rect 3809 49286 3861 49335
rect 3917 49286 3969 49335
rect 4025 49286 4077 49335
rect 4133 49286 4185 49335
rect 4241 49286 4293 49335
rect 4349 49286 4401 49335
rect 4457 49286 4509 49335
rect 4565 49286 4617 49335
rect 4673 49286 4725 49335
rect 5138 49286 5190 49335
rect 5246 49286 5298 49335
rect 5354 49286 5406 49335
rect 5462 49286 5514 49335
rect 5570 49286 5622 49335
rect 5678 49286 5730 49335
rect 5786 49286 5838 49335
rect 5894 49286 5946 49335
rect 6002 49286 6054 49335
rect 6110 49286 6162 49335
rect 6218 49286 6270 49335
rect 6326 49286 6378 49335
rect 6434 49286 6486 49335
rect 6542 49286 6594 49335
rect 6650 49286 6702 49335
rect 6758 49286 6810 49335
rect 6866 49286 6918 49335
rect 6974 49286 7026 49335
rect 7082 49286 7134 49335
rect 7844 49286 7896 49335
rect 7952 49286 8004 49335
rect 8060 49286 8112 49335
rect 8168 49286 8220 49335
rect 8276 49286 8328 49335
rect 8384 49286 8436 49335
rect 8492 49286 8544 49335
rect 8600 49286 8652 49335
rect 8708 49286 8760 49335
rect 8816 49286 8868 49335
rect 8924 49286 8976 49335
rect 9032 49286 9084 49335
rect 9140 49286 9192 49335
rect 9248 49286 9300 49335
rect 9356 49286 9408 49335
rect 9464 49286 9516 49335
rect 9572 49286 9624 49335
rect 9680 49286 9732 49335
rect 9788 49286 9840 49335
rect 10253 49286 10305 49335
rect 10361 49286 10413 49335
rect 10469 49286 10521 49335
rect 10577 49286 10629 49335
rect 10685 49286 10737 49335
rect 10793 49286 10845 49335
rect 10901 49286 10953 49335
rect 11009 49286 11061 49335
rect 11117 49286 11169 49335
rect 11225 49286 11277 49335
rect 11333 49286 11385 49335
rect 11441 49286 11493 49335
rect 11549 49286 11601 49335
rect 11657 49286 11709 49338
rect 11765 49286 11816 49338
rect 11816 49286 11817 49338
rect 3161 49178 3162 49230
rect 3162 49178 3213 49230
rect 3269 49178 3321 49230
rect 3377 49227 3429 49230
rect 3485 49227 3537 49230
rect 3593 49227 3645 49230
rect 3701 49227 3753 49230
rect 3809 49227 3861 49230
rect 3917 49227 3969 49230
rect 4025 49227 4077 49230
rect 4133 49227 4185 49230
rect 4241 49227 4293 49230
rect 4349 49227 4401 49230
rect 4457 49227 4509 49230
rect 4565 49227 4617 49230
rect 4673 49227 4725 49230
rect 5138 49227 5190 49230
rect 5246 49227 5298 49230
rect 5354 49227 5406 49230
rect 5462 49227 5514 49230
rect 5570 49227 5622 49230
rect 5678 49227 5730 49230
rect 5786 49227 5838 49230
rect 5894 49227 5946 49230
rect 6002 49227 6054 49230
rect 6110 49227 6162 49230
rect 6218 49227 6270 49230
rect 6326 49227 6378 49230
rect 6434 49227 6486 49230
rect 6542 49227 6594 49230
rect 6650 49227 6702 49230
rect 6758 49227 6810 49230
rect 6866 49227 6918 49230
rect 6974 49227 7026 49230
rect 7082 49227 7134 49230
rect 7844 49227 7896 49230
rect 7952 49227 8004 49230
rect 8060 49227 8112 49230
rect 8168 49227 8220 49230
rect 8276 49227 8328 49230
rect 8384 49227 8436 49230
rect 8492 49227 8544 49230
rect 8600 49227 8652 49230
rect 8708 49227 8760 49230
rect 8816 49227 8868 49230
rect 8924 49227 8976 49230
rect 9032 49227 9084 49230
rect 9140 49227 9192 49230
rect 9248 49227 9300 49230
rect 9356 49227 9408 49230
rect 9464 49227 9516 49230
rect 9572 49227 9624 49230
rect 9680 49227 9732 49230
rect 9788 49227 9840 49230
rect 10253 49227 10305 49230
rect 10361 49227 10413 49230
rect 10469 49227 10521 49230
rect 10577 49227 10629 49230
rect 10685 49227 10737 49230
rect 10793 49227 10845 49230
rect 10901 49227 10953 49230
rect 11009 49227 11061 49230
rect 11117 49227 11169 49230
rect 11225 49227 11277 49230
rect 11333 49227 11385 49230
rect 11441 49227 11493 49230
rect 11549 49227 11601 49230
rect 3377 49181 3429 49227
rect 3485 49181 3537 49227
rect 3593 49181 3645 49227
rect 3701 49181 3753 49227
rect 3809 49181 3861 49227
rect 3917 49181 3969 49227
rect 4025 49181 4077 49227
rect 4133 49181 4185 49227
rect 4241 49181 4293 49227
rect 4349 49181 4401 49227
rect 4457 49181 4509 49227
rect 4565 49181 4617 49227
rect 4673 49181 4725 49227
rect 5138 49181 5190 49227
rect 5246 49181 5298 49227
rect 5354 49181 5406 49227
rect 5462 49181 5514 49227
rect 5570 49181 5622 49227
rect 5678 49181 5730 49227
rect 5786 49181 5838 49227
rect 5894 49181 5946 49227
rect 6002 49181 6054 49227
rect 6110 49181 6162 49227
rect 6218 49181 6270 49227
rect 6326 49181 6378 49227
rect 6434 49181 6486 49227
rect 6542 49181 6594 49227
rect 6650 49181 6702 49227
rect 6758 49181 6810 49227
rect 6866 49181 6918 49227
rect 6974 49181 7026 49227
rect 7082 49181 7134 49227
rect 7844 49181 7896 49227
rect 7952 49181 8004 49227
rect 8060 49181 8112 49227
rect 8168 49181 8220 49227
rect 8276 49181 8328 49227
rect 8384 49181 8436 49227
rect 8492 49181 8544 49227
rect 8600 49181 8652 49227
rect 8708 49181 8760 49227
rect 8816 49181 8868 49227
rect 8924 49181 8976 49227
rect 9032 49181 9084 49227
rect 9140 49181 9192 49227
rect 9248 49181 9300 49227
rect 9356 49181 9408 49227
rect 9464 49181 9516 49227
rect 9572 49181 9624 49227
rect 9680 49181 9732 49227
rect 9788 49181 9840 49227
rect 10253 49181 10305 49227
rect 10361 49181 10413 49227
rect 10469 49181 10521 49227
rect 10577 49181 10629 49227
rect 10685 49181 10737 49227
rect 10793 49181 10845 49227
rect 10901 49181 10953 49227
rect 11009 49181 11061 49227
rect 11117 49181 11169 49227
rect 11225 49181 11277 49227
rect 11333 49181 11385 49227
rect 11441 49181 11493 49227
rect 11549 49181 11601 49227
rect 3377 49178 3429 49181
rect 3485 49178 3537 49181
rect 3593 49178 3645 49181
rect 3701 49178 3753 49181
rect 3809 49178 3861 49181
rect 3917 49178 3969 49181
rect 4025 49178 4077 49181
rect 4133 49178 4185 49181
rect 4241 49178 4293 49181
rect 4349 49178 4401 49181
rect 4457 49178 4509 49181
rect 4565 49178 4617 49181
rect 4673 49178 4725 49181
rect 5138 49178 5190 49181
rect 5246 49178 5298 49181
rect 5354 49178 5406 49181
rect 5462 49178 5514 49181
rect 5570 49178 5622 49181
rect 5678 49178 5730 49181
rect 5786 49178 5838 49181
rect 5894 49178 5946 49181
rect 6002 49178 6054 49181
rect 6110 49178 6162 49181
rect 6218 49178 6270 49181
rect 6326 49178 6378 49181
rect 6434 49178 6486 49181
rect 6542 49178 6594 49181
rect 6650 49178 6702 49181
rect 6758 49178 6810 49181
rect 6866 49178 6918 49181
rect 6974 49178 7026 49181
rect 7082 49178 7134 49181
rect 7844 49178 7896 49181
rect 7952 49178 8004 49181
rect 8060 49178 8112 49181
rect 8168 49178 8220 49181
rect 8276 49178 8328 49181
rect 8384 49178 8436 49181
rect 8492 49178 8544 49181
rect 8600 49178 8652 49181
rect 8708 49178 8760 49181
rect 8816 49178 8868 49181
rect 8924 49178 8976 49181
rect 9032 49178 9084 49181
rect 9140 49178 9192 49181
rect 9248 49178 9300 49181
rect 9356 49178 9408 49181
rect 9464 49178 9516 49181
rect 9572 49178 9624 49181
rect 9680 49178 9732 49181
rect 9788 49178 9840 49181
rect 10253 49178 10305 49181
rect 10361 49178 10413 49181
rect 10469 49178 10521 49181
rect 10577 49178 10629 49181
rect 10685 49178 10737 49181
rect 10793 49178 10845 49181
rect 10901 49178 10953 49181
rect 11009 49178 11061 49181
rect 11117 49178 11169 49181
rect 11225 49178 11277 49181
rect 11333 49178 11385 49181
rect 11441 49178 11493 49181
rect 11549 49178 11601 49181
rect 11657 49178 11709 49230
rect 11765 49178 11816 49230
rect 11816 49178 11817 49230
rect 3161 49070 3162 49122
rect 3162 49070 3213 49122
rect 3269 49070 3321 49122
rect 3377 49073 3429 49122
rect 3485 49073 3537 49122
rect 3593 49073 3645 49122
rect 3701 49073 3753 49122
rect 3809 49073 3861 49122
rect 3917 49073 3969 49122
rect 4025 49073 4077 49122
rect 4133 49073 4185 49122
rect 4241 49073 4293 49122
rect 4349 49073 4401 49122
rect 4457 49073 4509 49122
rect 4565 49073 4617 49122
rect 4673 49073 4725 49122
rect 5138 49073 5190 49122
rect 5246 49073 5298 49122
rect 5354 49073 5406 49122
rect 5462 49073 5514 49122
rect 5570 49073 5622 49122
rect 5678 49073 5730 49122
rect 5786 49073 5838 49122
rect 5894 49073 5946 49122
rect 6002 49073 6054 49122
rect 6110 49073 6162 49122
rect 6218 49073 6270 49122
rect 6326 49073 6378 49122
rect 6434 49073 6486 49122
rect 6542 49073 6594 49122
rect 6650 49073 6702 49122
rect 6758 49073 6810 49122
rect 6866 49073 6918 49122
rect 6974 49073 7026 49122
rect 7082 49073 7134 49122
rect 7844 49073 7896 49122
rect 7952 49073 8004 49122
rect 8060 49073 8112 49122
rect 8168 49073 8220 49122
rect 8276 49073 8328 49122
rect 8384 49073 8436 49122
rect 8492 49073 8544 49122
rect 8600 49073 8652 49122
rect 8708 49073 8760 49122
rect 8816 49073 8868 49122
rect 8924 49073 8976 49122
rect 9032 49073 9084 49122
rect 9140 49073 9192 49122
rect 9248 49073 9300 49122
rect 9356 49073 9408 49122
rect 9464 49073 9516 49122
rect 9572 49073 9624 49122
rect 9680 49073 9732 49122
rect 9788 49073 9840 49122
rect 10253 49073 10305 49122
rect 10361 49073 10413 49122
rect 10469 49073 10521 49122
rect 10577 49073 10629 49122
rect 10685 49073 10737 49122
rect 10793 49073 10845 49122
rect 10901 49073 10953 49122
rect 11009 49073 11061 49122
rect 11117 49073 11169 49122
rect 11225 49073 11277 49122
rect 11333 49073 11385 49122
rect 11441 49073 11493 49122
rect 11549 49073 11601 49122
rect 3377 49070 3424 49073
rect 3424 49070 3429 49073
rect 3485 49070 3537 49073
rect 3593 49070 3645 49073
rect 3701 49070 3753 49073
rect 3809 49070 3861 49073
rect 3917 49070 3969 49073
rect 4025 49070 4077 49073
rect 4133 49070 4185 49073
rect 4241 49070 4293 49073
rect 4349 49070 4401 49073
rect 4457 49070 4509 49073
rect 4565 49070 4617 49073
rect 4673 49070 4725 49073
rect 5138 49070 5190 49073
rect 5246 49070 5298 49073
rect 5354 49070 5406 49073
rect 5462 49070 5514 49073
rect 5570 49070 5622 49073
rect 5678 49070 5730 49073
rect 5786 49070 5838 49073
rect 5894 49070 5946 49073
rect 6002 49070 6054 49073
rect 6110 49070 6162 49073
rect 6218 49070 6270 49073
rect 6326 49070 6378 49073
rect 6434 49070 6486 49073
rect 6542 49070 6594 49073
rect 6650 49070 6702 49073
rect 6758 49070 6810 49073
rect 6866 49070 6918 49073
rect 6974 49070 7026 49073
rect 7082 49070 7134 49073
rect 7844 49070 7896 49073
rect 7952 49070 8004 49073
rect 8060 49070 8112 49073
rect 8168 49070 8220 49073
rect 8276 49070 8328 49073
rect 8384 49070 8436 49073
rect 8492 49070 8544 49073
rect 8600 49070 8652 49073
rect 8708 49070 8760 49073
rect 8816 49070 8868 49073
rect 8924 49070 8976 49073
rect 9032 49070 9084 49073
rect 9140 49070 9192 49073
rect 9248 49070 9300 49073
rect 9356 49070 9408 49073
rect 9464 49070 9516 49073
rect 9572 49070 9624 49073
rect 9680 49070 9732 49073
rect 9788 49070 9840 49073
rect 10253 49070 10305 49073
rect 10361 49070 10413 49073
rect 10469 49070 10521 49073
rect 10577 49070 10629 49073
rect 10685 49070 10737 49073
rect 10793 49070 10845 49073
rect 10901 49070 10953 49073
rect 11009 49070 11061 49073
rect 11117 49070 11169 49073
rect 11225 49070 11277 49073
rect 11333 49070 11385 49073
rect 11441 49070 11493 49073
rect 11549 49070 11554 49073
rect 11554 49070 11601 49073
rect 11657 49070 11709 49122
rect 11765 49070 11816 49122
rect 11816 49070 11817 49122
rect 4871 48778 4923 48817
rect 4979 48778 5031 48817
rect 7247 48778 7299 48817
rect 7355 48778 7407 48817
rect 7463 48778 7515 48817
rect 7571 48778 7623 48817
rect 7679 48778 7731 48817
rect 9947 48778 9999 48817
rect 10055 48778 10107 48817
rect 4871 48765 4923 48778
rect 4979 48765 5031 48778
rect 7247 48765 7299 48778
rect 7355 48765 7407 48778
rect 7463 48765 7515 48778
rect 7571 48765 7623 48778
rect 7679 48765 7731 48778
rect 9947 48765 9999 48778
rect 10055 48765 10107 48778
rect 4871 48696 4923 48709
rect 4979 48696 5031 48709
rect 7247 48696 7299 48709
rect 7355 48696 7407 48709
rect 7463 48696 7515 48709
rect 7571 48696 7623 48709
rect 7679 48696 7731 48709
rect 9947 48696 9999 48709
rect 10055 48696 10107 48709
rect 4871 48657 4923 48696
rect 4979 48657 5031 48696
rect 7247 48657 7299 48696
rect 7355 48657 7407 48696
rect 7463 48657 7515 48696
rect 7571 48657 7623 48696
rect 7679 48657 7731 48696
rect 9947 48657 9999 48696
rect 10055 48657 10107 48696
rect 3161 48376 3162 48427
rect 3162 48376 3213 48427
rect 3161 48375 3213 48376
rect 3269 48375 3321 48427
rect 3377 48401 3424 48427
rect 3424 48401 3429 48427
rect 3485 48401 3537 48427
rect 3593 48401 3645 48427
rect 3701 48401 3753 48427
rect 3809 48401 3861 48427
rect 3917 48401 3969 48427
rect 4025 48401 4077 48427
rect 4133 48401 4185 48427
rect 4241 48401 4293 48427
rect 4349 48401 4401 48427
rect 4457 48401 4509 48427
rect 4565 48401 4617 48427
rect 4673 48401 4725 48427
rect 5138 48401 5190 48427
rect 5246 48401 5298 48427
rect 5354 48401 5406 48427
rect 5462 48401 5514 48427
rect 5570 48401 5622 48427
rect 5678 48401 5730 48427
rect 5786 48401 5838 48427
rect 5894 48401 5946 48427
rect 6002 48401 6054 48427
rect 6110 48401 6162 48427
rect 6218 48401 6270 48427
rect 6326 48401 6378 48427
rect 6434 48401 6486 48427
rect 6542 48401 6594 48427
rect 6650 48401 6702 48427
rect 6758 48401 6810 48427
rect 6866 48401 6918 48427
rect 6974 48401 7026 48427
rect 7082 48401 7134 48427
rect 7844 48401 7896 48427
rect 7952 48401 8004 48427
rect 8060 48401 8112 48427
rect 8168 48401 8220 48427
rect 8276 48401 8328 48427
rect 8384 48401 8436 48427
rect 8492 48401 8544 48427
rect 8600 48401 8652 48427
rect 8708 48401 8760 48427
rect 8816 48401 8868 48427
rect 8924 48401 8976 48427
rect 9032 48401 9084 48427
rect 9140 48401 9192 48427
rect 9248 48401 9300 48427
rect 9356 48401 9408 48427
rect 9464 48401 9516 48427
rect 9572 48401 9624 48427
rect 9680 48401 9732 48427
rect 9788 48401 9840 48427
rect 10253 48401 10305 48427
rect 10361 48401 10413 48427
rect 10469 48401 10521 48427
rect 10577 48401 10629 48427
rect 10685 48401 10737 48427
rect 10793 48401 10845 48427
rect 10901 48401 10953 48427
rect 11009 48401 11061 48427
rect 11117 48401 11169 48427
rect 11225 48401 11277 48427
rect 11333 48401 11385 48427
rect 11441 48401 11493 48427
rect 11549 48401 11554 48427
rect 11554 48401 11601 48427
rect 3377 48375 3429 48401
rect 3485 48375 3537 48401
rect 3593 48375 3645 48401
rect 3701 48375 3753 48401
rect 3809 48375 3861 48401
rect 3917 48375 3969 48401
rect 4025 48375 4077 48401
rect 4133 48375 4185 48401
rect 4241 48375 4293 48401
rect 4349 48375 4401 48401
rect 4457 48375 4509 48401
rect 4565 48375 4617 48401
rect 4673 48375 4725 48401
rect 5138 48375 5190 48401
rect 5246 48375 5298 48401
rect 5354 48375 5406 48401
rect 5462 48375 5514 48401
rect 5570 48375 5622 48401
rect 5678 48375 5730 48401
rect 5786 48375 5838 48401
rect 5894 48375 5946 48401
rect 6002 48375 6054 48401
rect 6110 48375 6162 48401
rect 6218 48375 6270 48401
rect 6326 48375 6378 48401
rect 6434 48375 6486 48401
rect 6542 48375 6594 48401
rect 6650 48375 6702 48401
rect 6758 48375 6810 48401
rect 6866 48375 6918 48401
rect 6974 48375 7026 48401
rect 7082 48375 7134 48401
rect 7844 48375 7896 48401
rect 7952 48375 8004 48401
rect 8060 48375 8112 48401
rect 8168 48375 8220 48401
rect 8276 48375 8328 48401
rect 8384 48375 8436 48401
rect 8492 48375 8544 48401
rect 8600 48375 8652 48401
rect 8708 48375 8760 48401
rect 8816 48375 8868 48401
rect 8924 48375 8976 48401
rect 9032 48375 9084 48401
rect 9140 48375 9192 48401
rect 9248 48375 9300 48401
rect 9356 48375 9408 48401
rect 9464 48375 9516 48401
rect 9572 48375 9624 48401
rect 9680 48375 9732 48401
rect 9788 48375 9840 48401
rect 10253 48375 10305 48401
rect 10361 48375 10413 48401
rect 10469 48375 10521 48401
rect 10577 48375 10629 48401
rect 10685 48375 10737 48401
rect 10793 48375 10845 48401
rect 10901 48375 10953 48401
rect 11009 48375 11061 48401
rect 11117 48375 11169 48401
rect 11225 48375 11277 48401
rect 11333 48375 11385 48401
rect 11441 48375 11493 48401
rect 11549 48375 11601 48401
rect 11657 48375 11709 48427
rect 11765 48376 11816 48427
rect 11816 48376 11817 48427
rect 11765 48375 11817 48376
rect 3161 48293 3213 48319
rect 3269 48293 3321 48319
rect 3377 48293 3429 48319
rect 3485 48293 3537 48319
rect 3593 48293 3645 48319
rect 3701 48293 3753 48319
rect 3809 48293 3861 48319
rect 3917 48293 3969 48319
rect 4025 48293 4077 48319
rect 4133 48293 4185 48319
rect 4241 48293 4293 48319
rect 4349 48293 4401 48319
rect 4457 48293 4509 48319
rect 4565 48293 4617 48319
rect 4673 48293 4725 48319
rect 5138 48293 5190 48319
rect 5246 48293 5298 48319
rect 5354 48293 5406 48319
rect 5462 48293 5514 48319
rect 5570 48293 5622 48319
rect 5678 48293 5730 48319
rect 5786 48293 5838 48319
rect 5894 48293 5946 48319
rect 6002 48293 6054 48319
rect 6110 48293 6162 48319
rect 6218 48293 6270 48319
rect 6326 48293 6378 48319
rect 6434 48293 6486 48319
rect 6542 48293 6594 48319
rect 6650 48293 6702 48319
rect 6758 48293 6810 48319
rect 6866 48293 6918 48319
rect 6974 48293 7026 48319
rect 7082 48293 7134 48319
rect 7844 48293 7896 48319
rect 7952 48293 8004 48319
rect 8060 48293 8112 48319
rect 8168 48293 8220 48319
rect 8276 48293 8328 48319
rect 8384 48293 8436 48319
rect 8492 48293 8544 48319
rect 8600 48293 8652 48319
rect 8708 48293 8760 48319
rect 8816 48293 8868 48319
rect 8924 48293 8976 48319
rect 9032 48293 9084 48319
rect 9140 48293 9192 48319
rect 9248 48293 9300 48319
rect 9356 48293 9408 48319
rect 9464 48293 9516 48319
rect 9572 48293 9624 48319
rect 9680 48293 9732 48319
rect 9788 48293 9840 48319
rect 10253 48293 10305 48319
rect 10361 48293 10413 48319
rect 10469 48293 10521 48319
rect 10577 48293 10629 48319
rect 10685 48293 10737 48319
rect 10793 48293 10845 48319
rect 10901 48293 10953 48319
rect 11009 48293 11061 48319
rect 11117 48293 11169 48319
rect 11225 48293 11277 48319
rect 11333 48293 11385 48319
rect 11441 48293 11493 48319
rect 11549 48293 11601 48319
rect 11657 48293 11709 48319
rect 11765 48293 11817 48319
rect 3161 48267 3213 48293
rect 3269 48267 3321 48293
rect 3377 48267 3429 48293
rect 3485 48267 3537 48293
rect 3593 48267 3645 48293
rect 3701 48267 3753 48293
rect 3809 48267 3861 48293
rect 3917 48267 3969 48293
rect 4025 48267 4077 48293
rect 4133 48267 4185 48293
rect 4241 48267 4293 48293
rect 4349 48267 4401 48293
rect 4457 48267 4509 48293
rect 4565 48267 4617 48293
rect 4673 48267 4725 48293
rect 5138 48267 5190 48293
rect 5246 48267 5298 48293
rect 5354 48267 5406 48293
rect 5462 48267 5514 48293
rect 5570 48267 5622 48293
rect 5678 48267 5730 48293
rect 5786 48267 5838 48293
rect 5894 48267 5946 48293
rect 6002 48267 6054 48293
rect 6110 48267 6162 48293
rect 6218 48267 6270 48293
rect 6326 48267 6378 48293
rect 6434 48267 6486 48293
rect 6542 48267 6594 48293
rect 6650 48267 6702 48293
rect 6758 48267 6810 48293
rect 6866 48267 6918 48293
rect 6974 48267 7026 48293
rect 7082 48267 7134 48293
rect 7844 48267 7896 48293
rect 7952 48267 8004 48293
rect 8060 48267 8112 48293
rect 8168 48267 8220 48293
rect 8276 48267 8328 48293
rect 8384 48267 8436 48293
rect 8492 48267 8544 48293
rect 8600 48267 8652 48293
rect 8708 48267 8760 48293
rect 8816 48267 8868 48293
rect 8924 48267 8976 48293
rect 9032 48267 9084 48293
rect 9140 48267 9192 48293
rect 9248 48267 9300 48293
rect 9356 48267 9408 48293
rect 9464 48267 9516 48293
rect 9572 48267 9624 48293
rect 9680 48267 9732 48293
rect 9788 48267 9840 48293
rect 10253 48267 10305 48293
rect 10361 48267 10413 48293
rect 10469 48267 10521 48293
rect 10577 48267 10629 48293
rect 10685 48267 10737 48293
rect 10793 48267 10845 48293
rect 10901 48267 10953 48293
rect 11009 48267 11061 48293
rect 11117 48267 11169 48293
rect 11225 48267 11277 48293
rect 11333 48267 11385 48293
rect 11441 48267 11493 48293
rect 11549 48267 11601 48293
rect 11657 48267 11709 48293
rect 11765 48267 11817 48293
rect 12336 52218 12388 52270
rect 12336 52110 12388 52162
rect 12336 52002 12388 52054
rect 12336 51894 12388 51946
rect 12336 51786 12388 51838
rect 12336 51678 12388 51730
rect 12336 51570 12388 51622
rect 12336 51462 12388 51514
rect 12336 51354 12388 51406
rect 12336 51246 12388 51298
rect 12336 51138 12388 51190
rect 12336 51030 12388 51082
rect 12336 50922 12388 50974
rect 12336 50814 12388 50866
rect 12336 50706 12388 50758
rect 12336 50598 12388 50650
rect 12336 50490 12388 50542
rect 12336 50382 12388 50434
rect 12336 50274 12388 50326
rect 12336 50166 12388 50218
rect 12336 50058 12388 50110
rect 12336 49950 12388 50002
rect 12336 49842 12388 49894
rect 12336 49734 12388 49786
rect 12336 49626 12388 49678
rect 12336 49518 12388 49570
rect 12336 49410 12388 49462
rect 12336 49302 12388 49354
rect 12336 49194 12388 49246
rect 12336 49086 12388 49138
rect 12336 48978 12388 49030
rect 12336 48870 12388 48922
rect 12336 48762 12388 48814
rect 12336 48654 12388 48706
rect 12336 48546 12388 48598
rect 12336 48438 12388 48490
rect 12336 48330 12388 48382
rect 12336 48222 12388 48274
rect 12336 48114 12388 48166
rect 2590 47898 2642 47950
rect 2590 47790 2642 47842
rect 2590 47682 2642 47734
rect 4871 47920 4923 47972
rect 4979 47920 5031 47972
rect 7247 47920 7299 47972
rect 7355 47920 7407 47972
rect 7463 47920 7515 47972
rect 7571 47920 7623 47972
rect 7679 47920 7731 47972
rect 9947 47920 9999 47972
rect 10055 47920 10107 47972
rect 4871 47812 4923 47864
rect 4979 47812 5031 47864
rect 7247 47812 7299 47864
rect 7355 47812 7407 47864
rect 7463 47812 7515 47864
rect 7571 47812 7623 47864
rect 7679 47812 7731 47864
rect 9947 47812 9999 47864
rect 10055 47812 10107 47864
rect 4871 47704 4923 47756
rect 4979 47704 5031 47756
rect 7247 47704 7299 47756
rect 7355 47704 7407 47756
rect 7463 47704 7515 47756
rect 7571 47704 7623 47756
rect 7679 47704 7731 47756
rect 9947 47704 9999 47756
rect 10055 47704 10107 47756
rect 12336 48006 12388 48058
rect 12336 47898 12388 47950
rect 12336 47790 12388 47842
rect 12336 47682 12388 47734
rect 14904 52522 14956 52574
rect 14904 52414 14956 52466
rect 14904 52306 14956 52358
rect 14904 52198 14956 52250
rect 14904 52090 14956 52142
rect 14904 51982 14956 52034
rect 14904 51874 14956 51926
rect 14904 51766 14956 51818
rect 14904 51658 14956 51710
rect 14904 51550 14956 51602
rect 14904 51442 14956 51494
rect 14904 51334 14956 51386
rect 14904 51226 14956 51278
rect 14904 49322 14956 49374
rect 14904 49214 14956 49266
rect 14904 49106 14956 49158
rect 14904 48998 14956 49050
rect 14904 48890 14956 48942
rect 14904 48782 14956 48834
rect 14904 48674 14956 48726
rect 14904 48566 14956 48618
rect 14904 48458 14956 48510
rect 14904 48350 14956 48402
rect 14904 48242 14956 48294
rect 14904 48134 14956 48186
rect 14904 48026 14956 48078
rect 22 46122 74 46174
rect 22 46014 74 46066
rect 22 45906 74 45958
rect 22 45798 74 45850
rect 22 45690 74 45742
rect 22 45582 74 45634
rect 22 45474 74 45526
rect 22 45366 74 45418
rect 22 45258 74 45310
rect 22 45150 74 45202
rect 22 45042 74 45094
rect 22 44934 74 44986
rect 22 44826 74 44878
rect 14904 46122 14956 46174
rect 14904 46014 14956 46066
rect 14904 45906 14956 45958
rect 14904 45798 14956 45850
rect 14904 45690 14956 45742
rect 14904 45582 14956 45634
rect 14904 45474 14956 45526
rect 14904 45366 14956 45418
rect 14904 45258 14956 45310
rect 14904 45150 14956 45202
rect 14904 45042 14956 45094
rect 14904 44934 14956 44986
rect 14904 44826 14956 44878
rect 22 38122 74 38174
rect 22 38014 74 38066
rect 22 37906 74 37958
rect 22 37798 74 37850
rect 22 37690 74 37742
rect 22 37582 74 37634
rect 22 37474 74 37526
rect 22 37366 74 37418
rect 22 37258 74 37310
rect 22 37150 74 37202
rect 22 37042 74 37094
rect 22 36934 74 36986
rect 22 36826 74 36878
rect 22 36532 74 36584
rect 22 36424 74 36476
rect 22 36316 74 36368
rect 22 36208 74 36260
rect 22 36100 74 36152
rect 22 35992 74 36044
rect 22 35884 74 35936
rect 22 35776 74 35828
rect 22 35668 74 35720
rect 22 35560 74 35612
rect 22 35452 74 35504
rect 22 35344 74 35396
rect 22 35236 74 35288
rect 22 35128 74 35180
rect 22 35020 74 35072
rect 22 34912 74 34964
rect 22 34804 74 34856
rect 22 34696 74 34748
rect 22 34588 74 34640
rect 22 34480 74 34532
rect 22 34372 74 34424
rect 22 34264 74 34316
rect 22 34156 74 34208
rect 22 34048 74 34100
rect 22 33940 74 33992
rect 22 33832 74 33884
rect 22 33724 74 33776
rect 22 33616 74 33668
rect 22 28522 74 28574
rect 22 28414 74 28466
rect 22 28306 74 28358
rect 22 28198 74 28250
rect 22 28090 74 28142
rect 22 27982 74 28034
rect 22 27874 74 27926
rect 22 27766 74 27818
rect 22 27658 74 27710
rect 22 27550 74 27602
rect 22 27442 74 27494
rect 22 27334 74 27386
rect 22 27226 74 27278
rect 22 14122 74 14174
rect 22 14014 74 14066
rect 22 13906 74 13958
rect 22 13798 74 13850
rect 22 13690 74 13742
rect 22 13582 74 13634
rect 22 13474 74 13526
rect 22 13366 74 13418
rect 22 13258 74 13310
rect 22 13150 74 13202
rect 22 13042 74 13094
rect 22 12934 74 12986
rect 22 12826 74 12878
rect 22 10932 74 10984
rect 22 10824 74 10876
rect 22 10716 74 10768
rect 22 10608 74 10660
rect 22 10500 74 10552
rect 22 10392 74 10444
rect 22 10284 74 10336
rect 22 10176 74 10228
rect 22 10068 74 10120
rect 22 9960 74 10012
rect 22 9852 74 9904
rect 22 9744 74 9796
rect 22 9636 74 9688
rect 22 9528 74 9580
rect 22 9420 74 9472
rect 22 9312 74 9364
rect 22 9204 74 9256
rect 22 9096 74 9148
rect 22 8988 74 9040
rect 22 8880 74 8932
rect 22 8772 74 8824
rect 22 8664 74 8716
rect 22 8556 74 8608
rect 22 8448 74 8500
rect 22 8340 74 8392
rect 22 8232 74 8284
rect 22 8124 74 8176
rect 22 8016 74 8068
rect 22 7732 74 7784
rect 22 7624 74 7676
rect 22 7516 74 7568
rect 22 7408 74 7460
rect 22 7300 74 7352
rect 22 7192 74 7244
rect 22 7084 74 7136
rect 22 6976 74 7028
rect 22 6868 74 6920
rect 22 6760 74 6812
rect 22 6652 74 6704
rect 22 6544 74 6596
rect 22 6436 74 6488
rect 22 6328 74 6380
rect 22 6220 74 6272
rect 22 6112 74 6164
rect 22 6004 74 6056
rect 22 5896 74 5948
rect 22 5788 74 5840
rect 22 5680 74 5732
rect 22 5572 74 5624
rect 22 5464 74 5516
rect 22 5356 74 5408
rect 22 5248 74 5300
rect 22 5140 74 5192
rect 22 5032 74 5084
rect 22 4924 74 4976
rect 22 4816 74 4868
rect 22 4532 74 4584
rect 22 4424 74 4476
rect 22 4316 74 4368
rect 22 4208 74 4260
rect 22 4100 74 4152
rect 22 3992 74 4044
rect 22 3884 74 3936
rect 22 3776 74 3828
rect 22 3668 74 3720
rect 22 3560 74 3612
rect 22 3452 74 3504
rect 22 3344 74 3396
rect 22 3236 74 3288
rect 22 3128 74 3180
rect 22 3020 74 3072
rect 22 2912 74 2964
rect 22 2804 74 2856
rect 22 2696 74 2748
rect 22 2588 74 2640
rect 22 2480 74 2532
rect 22 2372 74 2424
rect 22 2264 74 2316
rect 22 2156 74 2208
rect 22 2048 74 2100
rect 22 1940 74 1992
rect 22 1832 74 1884
rect 22 1724 74 1776
rect 22 1616 74 1668
rect 14904 38122 14956 38174
rect 14904 38014 14956 38066
rect 14904 37906 14956 37958
rect 14904 37798 14956 37850
rect 14904 37690 14956 37742
rect 14904 37582 14956 37634
rect 14904 37474 14956 37526
rect 14904 37366 14956 37418
rect 14904 37258 14956 37310
rect 14904 37150 14956 37202
rect 14904 37042 14956 37094
rect 14904 36934 14956 36986
rect 14904 36826 14956 36878
rect 14904 36532 14956 36584
rect 14904 36424 14956 36476
rect 14904 36316 14956 36368
rect 14904 36208 14956 36260
rect 14904 36100 14956 36152
rect 14904 35992 14956 36044
rect 14904 35884 14956 35936
rect 14904 35776 14956 35828
rect 14904 35668 14956 35720
rect 14904 35560 14956 35612
rect 14904 35452 14956 35504
rect 14904 35344 14956 35396
rect 14904 35236 14956 35288
rect 14904 35128 14956 35180
rect 14904 35020 14956 35072
rect 14904 34912 14956 34964
rect 14904 34804 14956 34856
rect 14904 34696 14956 34748
rect 14904 34588 14956 34640
rect 14904 34480 14956 34532
rect 14904 34372 14956 34424
rect 14904 34264 14956 34316
rect 14904 34156 14956 34208
rect 14904 34048 14956 34100
rect 14904 33940 14956 33992
rect 14904 33832 14956 33884
rect 14904 33724 14956 33776
rect 14904 33616 14956 33668
rect 14904 28522 14956 28574
rect 14904 28414 14956 28466
rect 14904 28306 14956 28358
rect 14904 28198 14956 28250
rect 14904 28090 14956 28142
rect 14904 27982 14956 28034
rect 14904 27874 14956 27926
rect 14904 27766 14956 27818
rect 14904 27658 14956 27710
rect 14904 27550 14956 27602
rect 14904 27442 14956 27494
rect 14904 27334 14956 27386
rect 14904 27226 14956 27278
rect 14904 14122 14956 14174
rect 14904 14014 14956 14066
rect 14904 13906 14956 13958
rect 14904 13798 14956 13850
rect 14904 13690 14956 13742
rect 14904 13582 14956 13634
rect 14904 13474 14956 13526
rect 14904 13366 14956 13418
rect 14904 13258 14956 13310
rect 14904 13150 14956 13202
rect 14904 13042 14956 13094
rect 14904 12934 14956 12986
rect 14904 12826 14956 12878
rect 14904 10932 14956 10984
rect 14904 10824 14956 10876
rect 14904 10716 14956 10768
rect 14904 10608 14956 10660
rect 14904 10500 14956 10552
rect 14904 10392 14956 10444
rect 14904 10284 14956 10336
rect 14904 10176 14956 10228
rect 14904 10068 14956 10120
rect 14904 9960 14956 10012
rect 14904 9852 14956 9904
rect 14904 9744 14956 9796
rect 14904 9636 14956 9688
rect 14904 9528 14956 9580
rect 14904 9420 14956 9472
rect 14904 9312 14956 9364
rect 14904 9204 14956 9256
rect 14904 9096 14956 9148
rect 14904 8988 14956 9040
rect 14904 8880 14956 8932
rect 14904 8772 14956 8824
rect 14904 8664 14956 8716
rect 14904 8556 14956 8608
rect 14904 8448 14956 8500
rect 14904 8340 14956 8392
rect 14904 8232 14956 8284
rect 14904 8124 14956 8176
rect 14904 8016 14956 8068
rect 14904 7732 14956 7784
rect 14904 7624 14956 7676
rect 14904 7516 14956 7568
rect 14904 7408 14956 7460
rect 14904 7300 14956 7352
rect 14904 7192 14956 7244
rect 14904 7084 14956 7136
rect 14904 6976 14956 7028
rect 14904 6868 14956 6920
rect 14904 6760 14956 6812
rect 14904 6652 14956 6704
rect 14904 6544 14956 6596
rect 14904 6436 14956 6488
rect 14904 6328 14956 6380
rect 14904 6220 14956 6272
rect 14904 6112 14956 6164
rect 14904 6004 14956 6056
rect 14904 5896 14956 5948
rect 14904 5788 14956 5840
rect 14904 5680 14956 5732
rect 14904 5572 14956 5624
rect 14904 5464 14956 5516
rect 14904 5356 14956 5408
rect 14904 5248 14956 5300
rect 14904 5140 14956 5192
rect 14904 5032 14956 5084
rect 14904 4924 14956 4976
rect 14904 4816 14956 4868
rect 14904 4532 14956 4584
rect 14904 4424 14956 4476
rect 14904 4316 14956 4368
rect 14904 4208 14956 4260
rect 14904 4100 14956 4152
rect 14904 3992 14956 4044
rect 14904 3884 14956 3936
rect 14904 3776 14956 3828
rect 14904 3668 14956 3720
rect 14904 3560 14956 3612
rect 14904 3452 14956 3504
rect 14904 3344 14956 3396
rect 14904 3236 14956 3288
rect 14904 3128 14956 3180
rect 14904 3020 14956 3072
rect 14904 2912 14956 2964
rect 14904 2804 14956 2856
rect 14904 2696 14956 2748
rect 14904 2588 14956 2640
rect 14904 2480 14956 2532
rect 14904 2372 14956 2424
rect 14904 2264 14956 2316
rect 14904 2156 14956 2208
rect 14904 2048 14956 2100
rect 14904 1940 14956 1992
rect 14904 1832 14956 1884
rect 14904 1724 14956 1776
rect 14904 1616 14956 1668
<< metal2 >>
rect -11 57259 86 57271
rect -11 57207 22 57259
rect 74 57207 86 57259
rect -11 57151 86 57207
rect -11 57099 22 57151
rect 74 57099 86 57151
rect -11 57043 86 57099
rect -11 56991 22 57043
rect 74 56991 86 57043
rect -11 56935 86 56991
rect -11 56883 22 56935
rect 74 56883 86 56935
rect -11 56827 86 56883
rect -11 56775 22 56827
rect 74 56775 86 56827
rect -11 56719 86 56775
rect -11 56667 22 56719
rect 74 56667 86 56719
rect -11 56611 86 56667
rect -11 56559 22 56611
rect 74 56559 86 56611
rect -11 56503 86 56559
rect -11 56451 22 56503
rect 74 56451 86 56503
rect -11 56395 86 56451
rect -11 56343 22 56395
rect 74 56343 86 56395
rect -11 56287 86 56343
rect -11 56235 22 56287
rect 74 56235 86 56287
rect -11 56179 86 56235
rect -11 56127 22 56179
rect 74 56127 86 56179
rect -11 56071 86 56127
rect -11 56019 22 56071
rect 74 56019 86 56071
rect -11 54174 86 56019
rect -11 54122 22 54174
rect 74 54122 86 54174
rect -11 54066 86 54122
rect -11 54014 22 54066
rect 74 54014 86 54066
rect -11 53958 86 54014
rect -11 53906 22 53958
rect 74 53906 86 53958
rect -11 53850 86 53906
rect -11 53798 22 53850
rect 74 53798 86 53850
rect -11 53742 86 53798
rect -11 53690 22 53742
rect 74 53690 86 53742
rect -11 53634 86 53690
rect -11 53582 22 53634
rect 74 53582 86 53634
rect -11 53526 86 53582
rect -11 53474 22 53526
rect 74 53474 86 53526
rect -11 53418 86 53474
rect -11 53366 22 53418
rect 74 53366 86 53418
rect -11 53310 86 53366
rect -11 53258 22 53310
rect 74 53258 86 53310
rect -11 53202 86 53258
rect -11 53150 22 53202
rect 74 53150 86 53202
rect -11 53094 86 53150
rect -11 53042 22 53094
rect 74 53042 86 53094
rect -11 52986 86 53042
rect -11 52934 22 52986
rect 74 52934 86 52986
rect -11 52878 86 52934
rect -11 52826 22 52878
rect 74 52826 86 52878
rect -11 52576 86 52826
rect -11 51224 20 52576
rect 76 51224 86 52576
rect -11 49374 86 51224
rect -11 49322 22 49374
rect 74 49322 86 49374
rect -11 49266 86 49322
rect -11 49214 22 49266
rect 74 49214 86 49266
rect -11 49158 86 49214
rect -11 49106 22 49158
rect 74 49106 86 49158
rect -11 49050 86 49106
rect -11 48998 22 49050
rect 74 48998 86 49050
rect -11 48942 86 48998
rect -11 48890 22 48942
rect 74 48890 86 48942
rect -11 48834 86 48890
rect -11 48782 22 48834
rect 74 48782 86 48834
rect -11 48726 86 48782
rect -11 48674 22 48726
rect 74 48674 86 48726
rect -11 48618 86 48674
rect -11 48566 22 48618
rect 74 48566 86 48618
rect -11 48510 86 48566
rect -11 48458 22 48510
rect 74 48458 86 48510
rect -11 48402 86 48458
rect -11 48350 22 48402
rect 74 48350 86 48402
rect -11 48294 86 48350
rect -11 48242 22 48294
rect 74 48242 86 48294
rect -11 48186 86 48242
rect -11 48134 22 48186
rect 74 48134 86 48186
rect -11 48078 86 48134
rect -11 48026 22 48078
rect 74 48026 86 48078
rect -11 46174 86 48026
rect 261 57104 2161 57600
rect 261 57052 375 57104
rect 427 57052 483 57104
rect 535 57052 591 57104
rect 643 57052 699 57104
rect 751 57052 807 57104
rect 859 57052 915 57104
rect 967 57052 1023 57104
rect 1075 57052 1131 57104
rect 1183 57052 1239 57104
rect 1291 57052 1347 57104
rect 1399 57052 1455 57104
rect 1507 57052 1563 57104
rect 1615 57052 1671 57104
rect 1723 57052 1779 57104
rect 1831 57052 1887 57104
rect 1939 57052 1995 57104
rect 2047 57052 2161 57104
rect 261 56643 2161 57052
rect 261 56591 369 56643
rect 421 56591 493 56643
rect 545 56591 617 56643
rect 669 56591 741 56643
rect 793 56591 2161 56643
rect 261 56519 2161 56591
rect 261 56467 369 56519
rect 421 56467 493 56519
rect 545 56467 617 56519
rect 669 56467 741 56519
rect 793 56467 2161 56519
rect 261 56395 2161 56467
rect 261 56343 369 56395
rect 421 56343 493 56395
rect 545 56343 617 56395
rect 669 56343 741 56395
rect 793 56343 2161 56395
rect 261 56271 2161 56343
rect 261 56219 369 56271
rect 421 56219 493 56271
rect 545 56219 617 56271
rect 669 56219 741 56271
rect 793 56219 2161 56271
rect 261 56147 2161 56219
rect 261 56095 369 56147
rect 421 56095 493 56147
rect 545 56095 617 56147
rect 669 56095 741 56147
rect 793 56095 2161 56147
rect 261 56023 2161 56095
rect 261 55971 369 56023
rect 421 55971 493 56023
rect 545 55971 617 56023
rect 669 55971 741 56023
rect 793 55971 2161 56023
rect 261 55899 2161 55971
rect 261 55847 369 55899
rect 421 55847 493 55899
rect 545 55847 617 55899
rect 669 55847 741 55899
rect 793 55847 2161 55899
rect 261 55775 2161 55847
rect 261 55723 369 55775
rect 421 55723 493 55775
rect 545 55723 617 55775
rect 669 55723 741 55775
rect 793 55723 2161 55775
rect 261 55651 2161 55723
rect 261 55599 369 55651
rect 421 55599 493 55651
rect 545 55599 617 55651
rect 669 55599 741 55651
rect 793 55599 2161 55651
rect 261 55527 2161 55599
rect 261 55475 369 55527
rect 421 55475 493 55527
rect 545 55475 617 55527
rect 669 55475 741 55527
rect 793 55475 2161 55527
rect 261 55403 2161 55475
rect 261 55351 369 55403
rect 421 55351 493 55403
rect 545 55351 617 55403
rect 669 55351 741 55403
rect 793 55351 2161 55403
rect 261 55279 2161 55351
rect 261 55227 369 55279
rect 421 55227 493 55279
rect 545 55227 617 55279
rect 669 55227 741 55279
rect 793 55227 2161 55279
rect 261 55155 2161 55227
rect 261 55103 369 55155
rect 421 55103 493 55155
rect 545 55103 617 55155
rect 669 55103 741 55155
rect 793 55103 2161 55155
rect 261 55031 2161 55103
rect 261 54979 369 55031
rect 421 54979 493 55031
rect 545 54979 617 55031
rect 669 54979 741 55031
rect 793 54979 2161 55031
rect 261 54907 2161 54979
rect 261 54855 369 54907
rect 421 54855 493 54907
rect 545 54855 617 54907
rect 669 54855 741 54907
rect 793 54855 2161 54907
rect 261 54783 2161 54855
rect 261 54731 369 54783
rect 421 54731 493 54783
rect 545 54731 617 54783
rect 669 54731 741 54783
rect 793 54731 2161 54783
rect 261 54659 2161 54731
rect 261 54607 369 54659
rect 421 54607 493 54659
rect 545 54607 617 54659
rect 669 54607 741 54659
rect 793 54607 2161 54659
rect 261 54535 2161 54607
rect 261 54483 369 54535
rect 421 54483 493 54535
rect 545 54483 617 54535
rect 669 54483 741 54535
rect 793 54483 2161 54535
rect 261 54411 2161 54483
rect 261 54359 369 54411
rect 421 54359 493 54411
rect 545 54359 617 54411
rect 669 54359 741 54411
rect 793 54359 2161 54411
rect 261 54287 2161 54359
rect 261 54235 369 54287
rect 421 54235 493 54287
rect 545 54235 617 54287
rect 669 54235 741 54287
rect 793 54235 2161 54287
rect 261 54163 2161 54235
rect 261 54111 369 54163
rect 421 54111 493 54163
rect 545 54111 617 54163
rect 669 54111 741 54163
rect 793 54111 2161 54163
rect 261 54039 2161 54111
rect 261 53987 369 54039
rect 421 53987 493 54039
rect 545 53987 617 54039
rect 669 53987 741 54039
rect 793 53987 2161 54039
rect 261 53915 2161 53987
rect 261 53863 369 53915
rect 421 53863 493 53915
rect 545 53863 617 53915
rect 669 53863 741 53915
rect 793 53863 2161 53915
rect 261 53791 2161 53863
rect 261 53739 369 53791
rect 421 53739 493 53791
rect 545 53739 617 53791
rect 669 53739 741 53791
rect 793 53739 2161 53791
rect 261 53667 2161 53739
rect 261 53615 369 53667
rect 421 53615 493 53667
rect 545 53615 617 53667
rect 669 53615 741 53667
rect 793 53615 2161 53667
rect 261 53543 2161 53615
rect 261 53491 369 53543
rect 421 53491 493 53543
rect 545 53491 617 53543
rect 669 53491 741 53543
rect 793 53491 2161 53543
rect 261 53483 2161 53491
rect 261 53431 869 53483
rect 921 53431 977 53483
rect 1029 53431 1085 53483
rect 1137 53431 1193 53483
rect 1245 53431 1301 53483
rect 1353 53431 1409 53483
rect 1461 53431 1517 53483
rect 1569 53431 1625 53483
rect 1677 53431 1733 53483
rect 1785 53431 1841 53483
rect 1893 53431 1949 53483
rect 2001 53431 2057 53483
rect 2109 53431 2161 53483
rect 261 53419 2161 53431
rect 261 53367 369 53419
rect 421 53367 493 53419
rect 545 53367 617 53419
rect 669 53367 741 53419
rect 793 53375 2161 53419
rect 793 53367 869 53375
rect 261 53323 869 53367
rect 921 53323 977 53375
rect 1029 53323 1085 53375
rect 1137 53323 1193 53375
rect 1245 53323 1301 53375
rect 1353 53323 1409 53375
rect 1461 53323 1517 53375
rect 1569 53323 1625 53375
rect 1677 53323 1733 53375
rect 1785 53323 1841 53375
rect 1893 53323 1949 53375
rect 2001 53323 2057 53375
rect 2109 53323 2161 53375
rect 261 53295 2161 53323
rect 261 53243 369 53295
rect 421 53243 493 53295
rect 545 53243 617 53295
rect 669 53243 741 53295
rect 793 53267 2161 53295
rect 793 53243 869 53267
rect 261 53215 869 53243
rect 921 53215 977 53267
rect 1029 53215 1085 53267
rect 1137 53215 1193 53267
rect 1245 53215 1301 53267
rect 1353 53215 1409 53267
rect 1461 53215 1517 53267
rect 1569 53215 1625 53267
rect 1677 53215 1733 53267
rect 1785 53215 1841 53267
rect 1893 53215 1949 53267
rect 2001 53215 2057 53267
rect 2109 53215 2161 53267
rect 261 52548 2161 53215
rect 261 52492 315 52548
rect 371 52492 439 52548
rect 495 52492 563 52548
rect 619 52492 687 52548
rect 743 52492 811 52548
rect 867 52492 935 52548
rect 991 52492 1059 52548
rect 1115 52492 1183 52548
rect 1239 52492 1307 52548
rect 1363 52492 1431 52548
rect 1487 52492 1555 52548
rect 1611 52492 1679 52548
rect 1735 52492 1803 52548
rect 1859 52492 1927 52548
rect 1983 52492 2051 52548
rect 2107 52492 2161 52548
rect 261 52424 2161 52492
rect 261 52368 315 52424
rect 371 52368 439 52424
rect 495 52368 563 52424
rect 619 52368 687 52424
rect 743 52368 811 52424
rect 867 52368 935 52424
rect 991 52368 1059 52424
rect 1115 52368 1183 52424
rect 1239 52368 1307 52424
rect 1363 52368 1431 52424
rect 1487 52368 1555 52424
rect 1611 52368 1679 52424
rect 1735 52368 1803 52424
rect 1859 52368 1927 52424
rect 1983 52368 2051 52424
rect 2107 52368 2161 52424
rect 261 52300 2161 52368
rect 261 52244 315 52300
rect 371 52244 439 52300
rect 495 52244 563 52300
rect 619 52244 687 52300
rect 743 52244 811 52300
rect 867 52244 935 52300
rect 991 52244 1059 52300
rect 1115 52244 1183 52300
rect 1239 52244 1307 52300
rect 1363 52244 1431 52300
rect 1487 52244 1555 52300
rect 1611 52244 1679 52300
rect 1735 52244 1803 52300
rect 1859 52244 1927 52300
rect 1983 52244 2051 52300
rect 2107 52244 2161 52300
rect 261 52176 2161 52244
rect 261 52120 315 52176
rect 371 52120 439 52176
rect 495 52120 563 52176
rect 619 52120 687 52176
rect 743 52120 811 52176
rect 867 52120 935 52176
rect 991 52120 1059 52176
rect 1115 52120 1183 52176
rect 1239 52120 1307 52176
rect 1363 52120 1431 52176
rect 1487 52120 1555 52176
rect 1611 52120 1679 52176
rect 1735 52120 1803 52176
rect 1859 52120 1927 52176
rect 1983 52120 2051 52176
rect 2107 52120 2161 52176
rect 261 52052 2161 52120
rect 261 51996 315 52052
rect 371 51996 439 52052
rect 495 51996 563 52052
rect 619 51996 687 52052
rect 743 51996 811 52052
rect 867 51996 935 52052
rect 991 51996 1059 52052
rect 1115 51996 1183 52052
rect 1239 51996 1307 52052
rect 1363 51996 1431 52052
rect 1487 51996 1555 52052
rect 1611 51996 1679 52052
rect 1735 51996 1803 52052
rect 1859 51996 1927 52052
rect 1983 51996 2051 52052
rect 2107 51996 2161 52052
rect 261 51928 2161 51996
rect 261 51872 315 51928
rect 371 51872 439 51928
rect 495 51872 563 51928
rect 619 51872 687 51928
rect 743 51872 811 51928
rect 867 51872 935 51928
rect 991 51872 1059 51928
rect 1115 51872 1183 51928
rect 1239 51872 1307 51928
rect 1363 51872 1431 51928
rect 1487 51872 1555 51928
rect 1611 51872 1679 51928
rect 1735 51872 1803 51928
rect 1859 51872 1927 51928
rect 1983 51872 2051 51928
rect 2107 51872 2161 51928
rect 261 51804 2161 51872
rect 261 51748 315 51804
rect 371 51748 439 51804
rect 495 51748 563 51804
rect 619 51748 687 51804
rect 743 51748 811 51804
rect 867 51748 935 51804
rect 991 51748 1059 51804
rect 1115 51748 1183 51804
rect 1239 51748 1307 51804
rect 1363 51748 1431 51804
rect 1487 51748 1555 51804
rect 1611 51748 1679 51804
rect 1735 51748 1803 51804
rect 1859 51748 1927 51804
rect 1983 51748 2051 51804
rect 2107 51748 2161 51804
rect 261 51680 2161 51748
rect 261 51624 315 51680
rect 371 51624 439 51680
rect 495 51624 563 51680
rect 619 51624 687 51680
rect 743 51624 811 51680
rect 867 51624 935 51680
rect 991 51624 1059 51680
rect 1115 51624 1183 51680
rect 1239 51624 1307 51680
rect 1363 51624 1431 51680
rect 1487 51624 1555 51680
rect 1611 51624 1679 51680
rect 1735 51624 1803 51680
rect 1859 51624 1927 51680
rect 1983 51624 2051 51680
rect 2107 51624 2161 51680
rect 261 51556 2161 51624
rect 261 51500 315 51556
rect 371 51500 439 51556
rect 495 51500 563 51556
rect 619 51500 687 51556
rect 743 51500 811 51556
rect 867 51500 935 51556
rect 991 51500 1059 51556
rect 1115 51500 1183 51556
rect 1239 51500 1307 51556
rect 1363 51500 1431 51556
rect 1487 51500 1555 51556
rect 1611 51500 1679 51556
rect 1735 51500 1803 51556
rect 1859 51500 1927 51556
rect 1983 51500 2051 51556
rect 2107 51500 2161 51556
rect 261 51432 2161 51500
rect 261 51376 315 51432
rect 371 51376 439 51432
rect 495 51376 563 51432
rect 619 51376 687 51432
rect 743 51376 811 51432
rect 867 51376 935 51432
rect 991 51376 1059 51432
rect 1115 51376 1183 51432
rect 1239 51376 1307 51432
rect 1363 51376 1431 51432
rect 1487 51376 1555 51432
rect 1611 51376 1679 51432
rect 1735 51376 1803 51432
rect 1859 51376 1927 51432
rect 1983 51376 2051 51432
rect 2107 51376 2161 51432
rect 261 51308 2161 51376
rect 261 51252 315 51308
rect 371 51252 439 51308
rect 495 51252 563 51308
rect 619 51252 687 51308
rect 743 51252 811 51308
rect 867 51252 935 51308
rect 991 51252 1059 51308
rect 1115 51252 1183 51308
rect 1239 51252 1307 51308
rect 1363 51252 1431 51308
rect 1487 51252 1555 51308
rect 1611 51252 1679 51308
rect 1735 51252 1803 51308
rect 1859 51252 1927 51308
rect 1983 51252 2051 51308
rect 2107 51252 2161 51308
rect 261 47163 2161 51252
rect 2481 56741 2681 57278
rect 2481 56689 2501 56741
rect 2553 56689 2609 56741
rect 2661 56689 2681 56741
rect 2481 53621 2681 56689
rect 2481 53569 2501 53621
rect 2553 53569 2609 53621
rect 2661 53569 2681 53621
rect 2481 52594 2681 53569
rect 2481 52542 2590 52594
rect 2642 52542 2681 52594
rect 2481 52486 2681 52542
rect 2481 52434 2590 52486
rect 2642 52434 2681 52486
rect 2481 52378 2681 52434
rect 2481 52326 2590 52378
rect 2642 52326 2681 52378
rect 2481 52270 2681 52326
rect 2481 52218 2590 52270
rect 2642 52218 2681 52270
rect 2481 52162 2681 52218
rect 2481 52110 2590 52162
rect 2642 52110 2681 52162
rect 2481 52054 2681 52110
rect 2481 52002 2590 52054
rect 2642 52002 2681 52054
rect 2481 51946 2681 52002
rect 2481 51894 2590 51946
rect 2642 51894 2681 51946
rect 2481 51838 2681 51894
rect 2481 51786 2590 51838
rect 2642 51786 2681 51838
rect 2481 51730 2681 51786
rect 2481 51678 2590 51730
rect 2642 51678 2681 51730
rect 2481 51622 2681 51678
rect 2481 51570 2590 51622
rect 2642 51570 2681 51622
rect 2481 51514 2681 51570
rect 2481 51462 2590 51514
rect 2642 51462 2681 51514
rect 2481 51406 2681 51462
rect 2481 51354 2590 51406
rect 2642 51354 2681 51406
rect 2481 51298 2681 51354
rect 2481 51246 2590 51298
rect 2642 51246 2681 51298
rect 2481 51190 2681 51246
rect 2481 51138 2590 51190
rect 2642 51138 2681 51190
rect 2481 51082 2681 51138
rect 2481 51030 2590 51082
rect 2642 51030 2681 51082
rect 2292 50926 2368 51000
rect 2292 50870 2302 50926
rect 2358 50870 2368 50926
rect 2292 50794 2368 50870
rect 2292 50738 2302 50794
rect 2358 50738 2368 50794
rect 2292 50662 2368 50738
rect 2292 50606 2302 50662
rect 2358 50606 2368 50662
rect 2292 50530 2368 50606
rect 2292 50474 2302 50530
rect 2358 50474 2368 50530
rect 2292 50398 2368 50474
rect 2292 50342 2302 50398
rect 2358 50342 2368 50398
rect 2292 50266 2368 50342
rect 2292 50210 2302 50266
rect 2358 50210 2368 50266
rect 2292 50134 2368 50210
rect 2292 50078 2302 50134
rect 2358 50078 2368 50134
rect 2292 50002 2368 50078
rect 2292 49946 2302 50002
rect 2358 49946 2368 50002
rect 2292 49870 2368 49946
rect 2292 49814 2302 49870
rect 2358 49814 2368 49870
rect 2292 49738 2368 49814
rect 2292 49682 2302 49738
rect 2358 49682 2368 49738
rect -11 46122 22 46174
rect 74 46122 86 46174
rect -11 46066 86 46122
rect -11 46014 22 46066
rect 74 46014 86 46066
rect -11 45958 86 46014
rect -11 45906 22 45958
rect 74 45906 86 45958
rect -11 45850 86 45906
rect -11 45798 22 45850
rect 74 45798 86 45850
rect -11 45742 86 45798
rect -11 45690 22 45742
rect 74 45690 86 45742
rect -11 45634 86 45690
rect -11 45582 22 45634
rect 74 45582 86 45634
rect -11 45526 86 45582
rect -11 45474 22 45526
rect 74 45474 86 45526
rect -11 45418 86 45474
rect -11 45366 22 45418
rect 74 45366 86 45418
rect -11 45310 86 45366
rect -11 45258 22 45310
rect 74 45258 86 45310
rect -11 45202 86 45258
rect -11 45150 22 45202
rect 74 45150 86 45202
rect -11 45094 86 45150
rect -11 45042 22 45094
rect 74 45042 86 45094
rect -11 44986 86 45042
rect -11 44934 22 44986
rect 74 44934 86 44986
rect -11 44878 86 44934
rect -11 44826 22 44878
rect 74 44826 86 44878
rect 305 44842 2117 46158
rect -11 38176 86 44826
rect 2292 39727 2368 49682
rect 2481 50974 2681 51030
rect 2481 50948 2590 50974
rect 2642 50948 2681 50974
rect 2481 50892 2491 50948
rect 2547 50922 2590 50948
rect 2547 50892 2615 50922
rect 2671 50892 2681 50948
rect 2481 50866 2681 50892
rect 2481 50824 2590 50866
rect 2642 50824 2681 50866
rect 2481 50768 2491 50824
rect 2547 50814 2590 50824
rect 2547 50768 2615 50814
rect 2671 50768 2681 50824
rect 2481 50758 2681 50768
rect 2481 50706 2590 50758
rect 2642 50706 2681 50758
rect 2481 50700 2681 50706
rect 2481 50644 2491 50700
rect 2547 50650 2615 50700
rect 2547 50644 2590 50650
rect 2671 50644 2681 50700
rect 2481 50598 2590 50644
rect 2642 50598 2681 50644
rect 2481 50576 2681 50598
rect 2481 50520 2491 50576
rect 2547 50542 2615 50576
rect 2547 50520 2590 50542
rect 2671 50520 2681 50576
rect 2481 50490 2590 50520
rect 2642 50490 2681 50520
rect 2481 50452 2681 50490
rect 2481 50396 2491 50452
rect 2547 50434 2615 50452
rect 2547 50396 2590 50434
rect 2671 50396 2681 50452
rect 2481 50382 2590 50396
rect 2642 50382 2681 50396
rect 2481 50328 2681 50382
rect 2481 50272 2491 50328
rect 2547 50326 2615 50328
rect 2547 50274 2590 50326
rect 2547 50272 2615 50274
rect 2671 50272 2681 50328
rect 2481 50218 2681 50272
rect 2481 50204 2590 50218
rect 2642 50204 2681 50218
rect 2481 50148 2491 50204
rect 2547 50166 2590 50204
rect 2547 50148 2615 50166
rect 2671 50148 2681 50204
rect 2481 50110 2681 50148
rect 2481 50080 2590 50110
rect 2642 50080 2681 50110
rect 2481 50024 2491 50080
rect 2547 50058 2590 50080
rect 2547 50024 2615 50058
rect 2671 50024 2681 50080
rect 2481 50002 2681 50024
rect 2481 49956 2590 50002
rect 2642 49956 2681 50002
rect 2481 49900 2491 49956
rect 2547 49950 2590 49956
rect 2547 49900 2615 49950
rect 2671 49900 2681 49956
rect 2481 49894 2681 49900
rect 2481 49842 2590 49894
rect 2642 49842 2681 49894
rect 2481 49832 2681 49842
rect 2481 49776 2491 49832
rect 2547 49786 2615 49832
rect 2547 49776 2590 49786
rect 2671 49776 2681 49832
rect 2481 49734 2590 49776
rect 2642 49734 2681 49776
rect 2481 49708 2681 49734
rect 2481 49652 2491 49708
rect 2547 49678 2615 49708
rect 2547 49652 2590 49678
rect 2671 49652 2681 49708
rect 2481 49626 2590 49652
rect 2642 49626 2681 49652
rect 2481 49570 2681 49626
rect 2481 49518 2590 49570
rect 2642 49518 2681 49570
rect 2481 49462 2681 49518
rect 2481 49410 2590 49462
rect 2642 49410 2681 49462
rect 2481 49354 2681 49410
rect 2481 49302 2590 49354
rect 2642 49302 2681 49354
rect 2481 49246 2681 49302
rect 2481 49194 2590 49246
rect 2642 49194 2681 49246
rect 2481 49138 2681 49194
rect 2481 49086 2590 49138
rect 2642 49086 2681 49138
rect 2481 49030 2681 49086
rect 2481 48978 2590 49030
rect 2642 48978 2681 49030
rect 2481 48922 2681 48978
rect 2481 48870 2590 48922
rect 2642 48870 2681 48922
rect 2481 48814 2681 48870
rect 2481 48762 2590 48814
rect 2642 48762 2681 48814
rect 2481 48706 2681 48762
rect 2481 48654 2590 48706
rect 2642 48654 2681 48706
rect 2481 48598 2681 48654
rect 2481 48546 2590 48598
rect 2642 48546 2681 48598
rect 2481 48490 2681 48546
rect 2481 48438 2590 48490
rect 2642 48438 2681 48490
rect 2481 48382 2681 48438
rect 2481 48330 2590 48382
rect 2642 48330 2681 48382
rect 2481 48274 2681 48330
rect 2481 48222 2590 48274
rect 2642 48222 2681 48274
rect 2481 48166 2681 48222
rect 2481 48114 2590 48166
rect 2642 48114 2681 48166
rect 2481 48058 2681 48114
rect 2481 48006 2590 48058
rect 2642 48006 2681 48058
rect 2481 47950 2681 48006
rect 2481 47898 2590 47950
rect 2642 47898 2681 47950
rect 2481 47842 2681 47898
rect 2481 47790 2590 47842
rect 2642 47790 2681 47842
rect 2481 47734 2681 47790
rect 2481 47682 2590 47734
rect 2642 47682 2681 47734
rect 2481 46442 2681 47682
rect 2741 57104 4791 57600
rect 2741 57052 2768 57104
rect 2820 57052 2876 57104
rect 2928 57052 2984 57104
rect 3036 57052 3092 57104
rect 3144 57052 3200 57104
rect 3252 57052 3308 57104
rect 3360 57052 3416 57104
rect 3468 57052 3524 57104
rect 3576 57052 3632 57104
rect 3684 57052 3740 57104
rect 3792 57052 3848 57104
rect 3900 57052 3956 57104
rect 4008 57052 4064 57104
rect 4116 57052 4172 57104
rect 4224 57052 4280 57104
rect 4332 57052 4388 57104
rect 4440 57052 4496 57104
rect 4548 57052 4604 57104
rect 4656 57052 4712 57104
rect 4764 57052 4791 57104
rect 2741 56643 4791 57052
rect 2741 56591 3903 56643
rect 3955 56591 4027 56643
rect 4079 56591 4151 56643
rect 4203 56591 4791 56643
rect 2741 56519 4791 56591
rect 2741 56467 3903 56519
rect 3955 56467 4027 56519
rect 4079 56467 4151 56519
rect 4203 56467 4791 56519
rect 2741 56395 4791 56467
rect 2741 56343 3903 56395
rect 3955 56343 4027 56395
rect 4079 56343 4151 56395
rect 4203 56343 4791 56395
rect 2741 56271 4791 56343
rect 2741 56219 3903 56271
rect 3955 56219 4027 56271
rect 4079 56219 4151 56271
rect 4203 56219 4791 56271
rect 2741 56147 4791 56219
rect 2741 56095 3903 56147
rect 3955 56095 4027 56147
rect 4079 56095 4151 56147
rect 4203 56095 4791 56147
rect 2741 56023 4791 56095
rect 2741 55971 3903 56023
rect 3955 55971 4027 56023
rect 4079 55971 4151 56023
rect 4203 55971 4791 56023
rect 2741 55899 4791 55971
rect 2741 55847 3903 55899
rect 3955 55847 4027 55899
rect 4079 55847 4151 55899
rect 4203 55847 4791 55899
rect 2741 55775 4791 55847
rect 2741 55723 3903 55775
rect 3955 55723 4027 55775
rect 4079 55723 4151 55775
rect 4203 55723 4791 55775
rect 2741 55651 4791 55723
rect 2741 55599 3903 55651
rect 3955 55599 4027 55651
rect 4079 55599 4151 55651
rect 4203 55599 4791 55651
rect 2741 55527 4791 55599
rect 2741 55475 3903 55527
rect 3955 55475 4027 55527
rect 4079 55475 4151 55527
rect 4203 55475 4791 55527
rect 2741 55403 4791 55475
rect 2741 55351 3903 55403
rect 3955 55351 4027 55403
rect 4079 55351 4151 55403
rect 4203 55351 4791 55403
rect 2741 55279 4791 55351
rect 2741 55227 3903 55279
rect 3955 55227 4027 55279
rect 4079 55227 4151 55279
rect 4203 55227 4791 55279
rect 2741 55155 4791 55227
rect 2741 55103 3903 55155
rect 3955 55103 4027 55155
rect 4079 55103 4151 55155
rect 4203 55103 4791 55155
rect 2741 55031 4791 55103
rect 2741 54979 3903 55031
rect 3955 54979 4027 55031
rect 4079 54979 4151 55031
rect 4203 54979 4791 55031
rect 2741 54907 4791 54979
rect 2741 54855 3903 54907
rect 3955 54855 4027 54907
rect 4079 54855 4151 54907
rect 4203 54855 4791 54907
rect 2741 54783 4791 54855
rect 2741 54731 3903 54783
rect 3955 54731 4027 54783
rect 4079 54731 4151 54783
rect 4203 54731 4791 54783
rect 2741 54659 4791 54731
rect 2741 54607 3903 54659
rect 3955 54607 4027 54659
rect 4079 54607 4151 54659
rect 4203 54607 4791 54659
rect 2741 54535 4791 54607
rect 2741 54483 3903 54535
rect 3955 54483 4027 54535
rect 4079 54483 4151 54535
rect 4203 54483 4791 54535
rect 2741 54411 4791 54483
rect 2741 54359 3903 54411
rect 3955 54359 4027 54411
rect 4079 54359 4151 54411
rect 4203 54359 4791 54411
rect 2741 54287 4791 54359
rect 2741 54235 3903 54287
rect 3955 54235 4027 54287
rect 4079 54235 4151 54287
rect 4203 54235 4791 54287
rect 2741 54163 4791 54235
rect 2741 54111 3903 54163
rect 3955 54111 4027 54163
rect 4079 54111 4151 54163
rect 4203 54111 4791 54163
rect 2741 54039 4791 54111
rect 2741 53987 3903 54039
rect 3955 53987 4027 54039
rect 4079 53987 4151 54039
rect 4203 53987 4791 54039
rect 2741 53915 4791 53987
rect 2741 53863 3903 53915
rect 3955 53863 4027 53915
rect 4079 53863 4151 53915
rect 4203 53863 4791 53915
rect 2741 53791 4791 53863
rect 2741 53739 3903 53791
rect 3955 53739 4027 53791
rect 4079 53739 4151 53791
rect 4203 53739 4791 53791
rect 2741 53667 4791 53739
rect 2741 53615 3903 53667
rect 3955 53615 4027 53667
rect 4079 53615 4151 53667
rect 4203 53615 4791 53667
rect 2741 53543 4791 53615
rect 2741 53491 3903 53543
rect 3955 53491 4027 53543
rect 4079 53491 4151 53543
rect 4203 53491 4791 53543
rect 2741 53483 4791 53491
rect 2741 53431 2763 53483
rect 2815 53431 2871 53483
rect 2923 53431 2979 53483
rect 3031 53431 3087 53483
rect 3139 53431 3195 53483
rect 3247 53431 3303 53483
rect 3355 53431 3411 53483
rect 3463 53431 3519 53483
rect 3571 53431 3627 53483
rect 3679 53431 3735 53483
rect 3787 53431 4791 53483
rect 2741 53419 4791 53431
rect 2741 53375 3903 53419
rect 2741 53323 2763 53375
rect 2815 53323 2871 53375
rect 2923 53323 2979 53375
rect 3031 53323 3087 53375
rect 3139 53323 3195 53375
rect 3247 53323 3303 53375
rect 3355 53323 3411 53375
rect 3463 53323 3519 53375
rect 3571 53323 3627 53375
rect 3679 53323 3735 53375
rect 3787 53367 3903 53375
rect 3955 53367 4027 53419
rect 4079 53367 4151 53419
rect 4203 53367 4791 53419
rect 3787 53323 4791 53367
rect 2741 53295 4791 53323
rect 2741 53267 3903 53295
rect 2741 53215 2763 53267
rect 2815 53215 2871 53267
rect 2923 53215 2979 53267
rect 3031 53215 3087 53267
rect 3139 53215 3195 53267
rect 3247 53215 3303 53267
rect 3355 53215 3411 53267
rect 3463 53215 3519 53267
rect 3571 53215 3627 53267
rect 3679 53215 3735 53267
rect 3787 53243 3903 53267
rect 3955 53243 4027 53295
rect 4079 53243 4151 53295
rect 4203 53243 4791 53295
rect 3787 53215 4791 53243
rect 2741 52548 4791 53215
rect 2741 52492 2808 52548
rect 2864 52492 2932 52548
rect 2988 52492 3056 52548
rect 3112 52492 3180 52548
rect 3236 52492 3304 52548
rect 3360 52492 3428 52548
rect 3484 52492 3552 52548
rect 3608 52492 3676 52548
rect 3732 52492 3800 52548
rect 3856 52492 3924 52548
rect 3980 52492 4048 52548
rect 4104 52492 4172 52548
rect 4228 52492 4296 52548
rect 4352 52492 4420 52548
rect 4476 52492 4544 52548
rect 4600 52492 4668 52548
rect 4724 52492 4791 52548
rect 2741 52424 4791 52492
rect 2741 52368 2808 52424
rect 2864 52368 2932 52424
rect 2988 52368 3056 52424
rect 3112 52368 3180 52424
rect 3236 52368 3304 52424
rect 3360 52368 3428 52424
rect 3484 52368 3552 52424
rect 3608 52368 3676 52424
rect 3732 52368 3800 52424
rect 3856 52368 3924 52424
rect 3980 52368 4048 52424
rect 4104 52368 4172 52424
rect 4228 52368 4296 52424
rect 4352 52368 4420 52424
rect 4476 52368 4544 52424
rect 4600 52368 4668 52424
rect 4724 52368 4791 52424
rect 2741 52300 4791 52368
rect 2741 52244 2808 52300
rect 2864 52244 2932 52300
rect 2988 52244 3056 52300
rect 3112 52244 3180 52300
rect 3236 52244 3304 52300
rect 3360 52244 3428 52300
rect 3484 52244 3552 52300
rect 3608 52244 3676 52300
rect 3732 52244 3800 52300
rect 3856 52244 3924 52300
rect 3980 52244 4048 52300
rect 4104 52244 4172 52300
rect 4228 52244 4296 52300
rect 4352 52244 4420 52300
rect 4476 52244 4544 52300
rect 4600 52244 4668 52300
rect 4724 52244 4791 52300
rect 2741 52176 4791 52244
rect 2741 52120 2808 52176
rect 2864 52120 2932 52176
rect 2988 52120 3056 52176
rect 3112 52120 3180 52176
rect 3236 52120 3304 52176
rect 3360 52120 3428 52176
rect 3484 52120 3552 52176
rect 3608 52120 3676 52176
rect 3732 52120 3800 52176
rect 3856 52120 3924 52176
rect 3980 52120 4048 52176
rect 4104 52120 4172 52176
rect 4228 52120 4296 52176
rect 4352 52120 4420 52176
rect 4476 52120 4544 52176
rect 4600 52120 4668 52176
rect 4724 52120 4791 52176
rect 2741 52052 4791 52120
rect 2741 51996 2808 52052
rect 2864 51996 2932 52052
rect 2988 51996 3056 52052
rect 3112 52009 3180 52052
rect 3236 52009 3304 52052
rect 3360 52009 3428 52052
rect 3484 52009 3552 52052
rect 3608 52009 3676 52052
rect 3732 52009 3800 52052
rect 3856 52009 3924 52052
rect 3980 52009 4048 52052
rect 4104 52009 4172 52052
rect 4228 52009 4296 52052
rect 4352 52009 4420 52052
rect 4476 52009 4544 52052
rect 4600 52009 4668 52052
rect 4724 52009 4791 52052
rect 3112 51996 3161 52009
rect 3236 51996 3269 52009
rect 3360 51996 3377 52009
rect 3484 51996 3485 52009
rect 2741 51957 3161 51996
rect 3213 51957 3269 51996
rect 3321 51957 3377 51996
rect 3429 51957 3485 51996
rect 3537 51996 3552 52009
rect 3645 51996 3676 52009
rect 3753 51996 3800 52009
rect 3537 51957 3593 51996
rect 3645 51957 3701 51996
rect 3753 51957 3809 51996
rect 3861 51957 3917 52009
rect 3980 51996 4025 52009
rect 4104 51996 4133 52009
rect 4228 51996 4241 52009
rect 3969 51957 4025 51996
rect 4077 51957 4133 51996
rect 4185 51957 4241 51996
rect 4293 51996 4296 52009
rect 4401 51996 4420 52009
rect 4509 51996 4544 52009
rect 4617 51996 4668 52009
rect 4293 51957 4349 51996
rect 4401 51957 4457 51996
rect 4509 51957 4565 51996
rect 4617 51957 4673 51996
rect 4725 51957 4791 52009
rect 2741 51928 4791 51957
rect 2741 51872 2808 51928
rect 2864 51872 2932 51928
rect 2988 51872 3056 51928
rect 3112 51901 3180 51928
rect 3236 51901 3304 51928
rect 3360 51901 3428 51928
rect 3484 51901 3552 51928
rect 3608 51901 3676 51928
rect 3732 51901 3800 51928
rect 3856 51901 3924 51928
rect 3980 51901 4048 51928
rect 4104 51901 4172 51928
rect 4228 51901 4296 51928
rect 4352 51901 4420 51928
rect 4476 51901 4544 51928
rect 4600 51901 4668 51928
rect 4724 51901 4791 51928
rect 3112 51872 3161 51901
rect 3236 51872 3269 51901
rect 3360 51872 3377 51901
rect 3484 51872 3485 51901
rect 2741 51849 3161 51872
rect 3213 51849 3269 51872
rect 3321 51849 3377 51872
rect 3429 51849 3485 51872
rect 3537 51872 3552 51901
rect 3645 51872 3676 51901
rect 3753 51872 3800 51901
rect 3537 51849 3593 51872
rect 3645 51849 3701 51872
rect 3753 51849 3809 51872
rect 3861 51849 3917 51901
rect 3980 51872 4025 51901
rect 4104 51872 4133 51901
rect 4228 51872 4241 51901
rect 3969 51849 4025 51872
rect 4077 51849 4133 51872
rect 4185 51849 4241 51872
rect 4293 51872 4296 51901
rect 4401 51872 4420 51901
rect 4509 51872 4544 51901
rect 4617 51872 4668 51901
rect 4293 51849 4349 51872
rect 4401 51849 4457 51872
rect 4509 51849 4565 51872
rect 4617 51849 4673 51872
rect 4725 51849 4791 51901
rect 2741 51804 4791 51849
rect 2741 51748 2808 51804
rect 2864 51748 2932 51804
rect 2988 51748 3056 51804
rect 3112 51748 3180 51804
rect 3236 51748 3304 51804
rect 3360 51748 3428 51804
rect 3484 51748 3552 51804
rect 3608 51748 3676 51804
rect 3732 51748 3800 51804
rect 3856 51748 3924 51804
rect 3980 51748 4048 51804
rect 4104 51748 4172 51804
rect 4228 51748 4296 51804
rect 4352 51748 4420 51804
rect 4476 51748 4544 51804
rect 4600 51748 4668 51804
rect 4724 51748 4791 51804
rect 2741 51680 4791 51748
rect 2741 51624 2808 51680
rect 2864 51624 2932 51680
rect 2988 51624 3056 51680
rect 3112 51624 3180 51680
rect 3236 51624 3304 51680
rect 3360 51624 3428 51680
rect 3484 51624 3552 51680
rect 3608 51624 3676 51680
rect 3732 51624 3800 51680
rect 3856 51624 3924 51680
rect 3980 51624 4048 51680
rect 4104 51624 4172 51680
rect 4228 51624 4296 51680
rect 4352 51624 4420 51680
rect 4476 51624 4544 51680
rect 4600 51624 4668 51680
rect 4724 51624 4791 51680
rect 2741 51556 4791 51624
rect 2741 51500 2808 51556
rect 2864 51500 2932 51556
rect 2988 51500 3056 51556
rect 3112 51500 3180 51556
rect 3236 51500 3304 51556
rect 3360 51500 3428 51556
rect 3484 51500 3552 51556
rect 3608 51500 3676 51556
rect 3732 51500 3800 51556
rect 3856 51500 3924 51556
rect 3980 51500 4048 51556
rect 4104 51500 4172 51556
rect 4228 51500 4296 51556
rect 4352 51500 4420 51556
rect 4476 51500 4544 51556
rect 4600 51500 4668 51556
rect 4724 51500 4791 51556
rect 2741 51432 4791 51500
rect 2741 51376 2808 51432
rect 2864 51376 2932 51432
rect 2988 51376 3056 51432
rect 3112 51376 3180 51432
rect 3236 51376 3304 51432
rect 3360 51376 3428 51432
rect 3484 51376 3552 51432
rect 3608 51376 3676 51432
rect 3732 51376 3800 51432
rect 3856 51376 3924 51432
rect 3980 51376 4048 51432
rect 4104 51376 4172 51432
rect 4228 51376 4296 51432
rect 4352 51376 4420 51432
rect 4476 51376 4544 51432
rect 4600 51376 4668 51432
rect 4724 51376 4791 51432
rect 2741 51308 4791 51376
rect 2741 51252 2808 51308
rect 2864 51252 2932 51308
rect 2988 51252 3056 51308
rect 3112 51252 3180 51308
rect 3236 51252 3304 51308
rect 3360 51252 3428 51308
rect 3484 51252 3552 51308
rect 3608 51252 3676 51308
rect 3732 51252 3800 51308
rect 3856 51252 3924 51308
rect 3980 51252 4048 51308
rect 4104 51252 4172 51308
rect 4228 51252 4296 51308
rect 4352 51252 4420 51308
rect 4476 51252 4544 51308
rect 4600 51252 4668 51308
rect 4724 51252 4791 51308
rect 2741 51206 4791 51252
rect 2741 51154 3161 51206
rect 3213 51154 3269 51206
rect 3321 51154 3377 51206
rect 3429 51154 3485 51206
rect 3537 51154 3593 51206
rect 3645 51154 3701 51206
rect 3753 51154 3809 51206
rect 3861 51154 3917 51206
rect 3969 51154 4025 51206
rect 4077 51154 4133 51206
rect 4185 51154 4241 51206
rect 4293 51154 4349 51206
rect 4401 51154 4457 51206
rect 4509 51154 4565 51206
rect 4617 51154 4673 51206
rect 4725 51154 4791 51206
rect 2741 51098 4791 51154
rect 2741 51046 3161 51098
rect 3213 51046 3269 51098
rect 3321 51046 3377 51098
rect 3429 51046 3485 51098
rect 3537 51046 3593 51098
rect 3645 51046 3701 51098
rect 3753 51046 3809 51098
rect 3861 51046 3917 51098
rect 3969 51046 4025 51098
rect 4077 51046 4133 51098
rect 4185 51046 4241 51098
rect 4293 51046 4349 51098
rect 4401 51046 4457 51098
rect 4509 51046 4565 51098
rect 4617 51046 4673 51098
rect 4725 51046 4791 51098
rect 2741 50990 4791 51046
rect 2741 50938 3161 50990
rect 3213 50938 3269 50990
rect 3321 50938 3377 50990
rect 3429 50938 3485 50990
rect 3537 50938 3593 50990
rect 3645 50938 3701 50990
rect 3753 50938 3809 50990
rect 3861 50938 3917 50990
rect 3969 50938 4025 50990
rect 4077 50938 4133 50990
rect 4185 50938 4241 50990
rect 4293 50938 4349 50990
rect 4401 50938 4457 50990
rect 4509 50938 4565 50990
rect 4617 50938 4673 50990
rect 4725 50938 4791 50990
rect 2741 50272 4791 50938
rect 2741 50220 3161 50272
rect 3213 50220 3269 50272
rect 3321 50220 3377 50272
rect 3429 50220 3485 50272
rect 3537 50220 3593 50272
rect 3645 50220 3701 50272
rect 3753 50220 3809 50272
rect 3861 50220 3917 50272
rect 3969 50220 4025 50272
rect 4077 50220 4133 50272
rect 4185 50220 4241 50272
rect 4293 50220 4349 50272
rect 4401 50220 4457 50272
rect 4509 50220 4565 50272
rect 4617 50220 4673 50272
rect 4725 50220 4791 50272
rect 2741 50164 4791 50220
rect 2741 50112 3161 50164
rect 3213 50112 3269 50164
rect 3321 50112 3377 50164
rect 3429 50112 3485 50164
rect 3537 50112 3593 50164
rect 3645 50112 3701 50164
rect 3753 50112 3809 50164
rect 3861 50112 3917 50164
rect 3969 50112 4025 50164
rect 4077 50112 4133 50164
rect 4185 50112 4241 50164
rect 4293 50112 4349 50164
rect 4401 50112 4457 50164
rect 4509 50112 4565 50164
rect 4617 50112 4673 50164
rect 4725 50112 4791 50164
rect 2741 50056 4791 50112
rect 2741 50004 3161 50056
rect 3213 50004 3269 50056
rect 3321 50004 3377 50056
rect 3429 50004 3485 50056
rect 3537 50004 3593 50056
rect 3645 50004 3701 50056
rect 3753 50004 3809 50056
rect 3861 50004 3917 50056
rect 3969 50004 4025 50056
rect 4077 50004 4133 50056
rect 4185 50004 4241 50056
rect 4293 50004 4349 50056
rect 4401 50004 4457 50056
rect 4509 50004 4565 50056
rect 4617 50004 4673 50056
rect 4725 50004 4791 50056
rect 2741 49338 4791 50004
rect 2741 49286 3161 49338
rect 3213 49286 3269 49338
rect 3321 49286 3377 49338
rect 3429 49286 3485 49338
rect 3537 49286 3593 49338
rect 3645 49286 3701 49338
rect 3753 49286 3809 49338
rect 3861 49286 3917 49338
rect 3969 49286 4025 49338
rect 4077 49286 4133 49338
rect 4185 49286 4241 49338
rect 4293 49286 4349 49338
rect 4401 49286 4457 49338
rect 4509 49286 4565 49338
rect 4617 49286 4673 49338
rect 4725 49286 4791 49338
rect 2741 49230 4791 49286
rect 2741 49178 3161 49230
rect 3213 49178 3269 49230
rect 3321 49178 3377 49230
rect 3429 49178 3485 49230
rect 3537 49178 3593 49230
rect 3645 49178 3701 49230
rect 3753 49178 3809 49230
rect 3861 49178 3917 49230
rect 3969 49178 4025 49230
rect 4077 49178 4133 49230
rect 4185 49178 4241 49230
rect 4293 49178 4349 49230
rect 4401 49178 4457 49230
rect 4509 49178 4565 49230
rect 4617 49178 4673 49230
rect 4725 49178 4791 49230
rect 2741 49122 4791 49178
rect 2741 49070 3161 49122
rect 3213 49070 3269 49122
rect 3321 49070 3377 49122
rect 3429 49070 3485 49122
rect 3537 49070 3593 49122
rect 3645 49070 3701 49122
rect 3753 49070 3809 49122
rect 3861 49070 3917 49122
rect 3969 49070 4025 49122
rect 4077 49070 4133 49122
rect 4185 49070 4241 49122
rect 4293 49070 4349 49122
rect 4401 49070 4457 49122
rect 4509 49070 4565 49122
rect 4617 49070 4673 49122
rect 4725 49070 4791 49122
rect 2741 48427 4791 49070
rect 2741 48375 3161 48427
rect 3213 48375 3269 48427
rect 3321 48375 3377 48427
rect 3429 48375 3485 48427
rect 3537 48375 3593 48427
rect 3645 48375 3701 48427
rect 3753 48375 3809 48427
rect 3861 48375 3917 48427
rect 3969 48375 4025 48427
rect 4077 48375 4133 48427
rect 4185 48375 4241 48427
rect 4293 48375 4349 48427
rect 4401 48375 4457 48427
rect 4509 48375 4565 48427
rect 4617 48375 4673 48427
rect 4725 48375 4791 48427
rect 2741 48319 4791 48375
rect 2741 48267 3161 48319
rect 3213 48267 3269 48319
rect 3321 48267 3377 48319
rect 3429 48267 3485 48319
rect 3537 48267 3593 48319
rect 3645 48267 3701 48319
rect 3753 48267 3809 48319
rect 3861 48267 3917 48319
rect 3969 48267 4025 48319
rect 4077 48267 4133 48319
rect 4185 48267 4241 48319
rect 4293 48267 4349 48319
rect 4401 48267 4457 48319
rect 4509 48267 4565 48319
rect 4617 48267 4673 48319
rect 4725 48267 4791 48319
rect 2741 47163 4791 48267
rect 4851 56693 5051 57278
rect 4851 56641 4871 56693
rect 4923 56641 4979 56693
rect 5031 56641 5051 56693
rect 4851 56585 5051 56641
rect 4851 56533 4871 56585
rect 4923 56533 4979 56585
rect 5031 56533 5051 56585
rect 4851 56477 5051 56533
rect 4851 56425 4871 56477
rect 4923 56425 4979 56477
rect 5031 56425 5051 56477
rect 4851 56369 5051 56425
rect 4851 56317 4871 56369
rect 4923 56317 4979 56369
rect 5031 56317 5051 56369
rect 4851 56261 5051 56317
rect 4851 56209 4871 56261
rect 4923 56209 4979 56261
rect 5031 56209 5051 56261
rect 4851 56153 5051 56209
rect 4851 56101 4871 56153
rect 4923 56101 4979 56153
rect 5031 56101 5051 56153
rect 4851 56045 5051 56101
rect 4851 55993 4871 56045
rect 4923 55993 4979 56045
rect 5031 55993 5051 56045
rect 4851 55937 5051 55993
rect 4851 55885 4871 55937
rect 4923 55885 4979 55937
rect 5031 55885 5051 55937
rect 4851 55829 5051 55885
rect 4851 55777 4871 55829
rect 4923 55777 4979 55829
rect 5031 55777 5051 55829
rect 4851 55721 5051 55777
rect 4851 55669 4871 55721
rect 4923 55669 4979 55721
rect 5031 55669 5051 55721
rect 4851 55613 5051 55669
rect 4851 55561 4871 55613
rect 4923 55561 4979 55613
rect 5031 55561 5051 55613
rect 4851 55505 5051 55561
rect 4851 55453 4871 55505
rect 4923 55453 4979 55505
rect 5031 55453 5051 55505
rect 4851 55397 5051 55453
rect 4851 55345 4871 55397
rect 4923 55345 4979 55397
rect 5031 55345 5051 55397
rect 4851 55289 5051 55345
rect 4851 55237 4871 55289
rect 4923 55237 4979 55289
rect 5031 55237 5051 55289
rect 4851 55181 5051 55237
rect 4851 55129 4871 55181
rect 4923 55129 4979 55181
rect 5031 55129 5051 55181
rect 4851 55073 5051 55129
rect 4851 55021 4871 55073
rect 4923 55021 4979 55073
rect 5031 55021 5051 55073
rect 4851 54965 5051 55021
rect 4851 54913 4871 54965
rect 4923 54913 4979 54965
rect 5031 54913 5051 54965
rect 4851 54857 5051 54913
rect 4851 54805 4871 54857
rect 4923 54805 4979 54857
rect 5031 54805 5051 54857
rect 4851 54749 5051 54805
rect 4851 54697 4871 54749
rect 4923 54697 4979 54749
rect 5031 54697 5051 54749
rect 4851 54641 5051 54697
rect 4851 54589 4871 54641
rect 4923 54589 4979 54641
rect 5031 54589 5051 54641
rect 4851 54533 5051 54589
rect 4851 54481 4871 54533
rect 4923 54481 4979 54533
rect 5031 54481 5051 54533
rect 4851 54425 5051 54481
rect 4851 54373 4871 54425
rect 4923 54373 4979 54425
rect 5031 54373 5051 54425
rect 4851 54317 5051 54373
rect 4851 54265 4871 54317
rect 4923 54265 4979 54317
rect 5031 54265 5051 54317
rect 4851 54209 5051 54265
rect 4851 54157 4871 54209
rect 4923 54157 4979 54209
rect 5031 54157 5051 54209
rect 4851 54101 5051 54157
rect 4851 54049 4871 54101
rect 4923 54049 4979 54101
rect 5031 54049 5051 54101
rect 4851 53993 5051 54049
rect 4851 53941 4871 53993
rect 4923 53941 4979 53993
rect 5031 53941 5051 53993
rect 4851 53885 5051 53941
rect 4851 53833 4871 53885
rect 4923 53833 4979 53885
rect 5031 53833 5051 53885
rect 4851 53777 5051 53833
rect 4851 53725 4871 53777
rect 4923 53725 4979 53777
rect 5031 53725 5051 53777
rect 4851 53669 5051 53725
rect 4851 53617 4871 53669
rect 4923 53617 4979 53669
rect 5031 53617 5051 53669
rect 4851 52572 5051 53617
rect 4851 52520 4871 52572
rect 4923 52520 4979 52572
rect 5031 52520 5051 52572
rect 4851 52464 5051 52520
rect 4851 52412 4871 52464
rect 4923 52412 4979 52464
rect 5031 52412 5051 52464
rect 4851 52356 5051 52412
rect 4851 52304 4871 52356
rect 4923 52304 4979 52356
rect 5031 52304 5051 52356
rect 4851 51619 5051 52304
rect 4851 51567 4871 51619
rect 4923 51567 4979 51619
rect 5031 51567 5051 51619
rect 4851 51511 5051 51567
rect 4851 51459 4871 51511
rect 4923 51459 4979 51511
rect 5031 51459 5051 51511
rect 4851 50948 5051 51459
rect 4851 50892 4861 50948
rect 4917 50892 4985 50948
rect 5041 50892 5051 50948
rect 4851 50824 5051 50892
rect 4851 50768 4861 50824
rect 4917 50768 4985 50824
rect 5041 50768 5051 50824
rect 4851 50700 5051 50768
rect 4851 50644 4861 50700
rect 4917 50685 4985 50700
rect 4851 50633 4871 50644
rect 4923 50633 4979 50685
rect 5041 50644 5051 50700
rect 5031 50633 5051 50644
rect 4851 50577 5051 50633
rect 4851 50576 4871 50577
rect 4851 50520 4861 50576
rect 4923 50525 4979 50577
rect 5031 50576 5051 50577
rect 4917 50520 4985 50525
rect 5041 50520 5051 50576
rect 4851 50452 5051 50520
rect 4851 50396 4861 50452
rect 4917 50396 4985 50452
rect 5041 50396 5051 50452
rect 4851 50328 5051 50396
rect 4851 50272 4861 50328
rect 4917 50272 4985 50328
rect 5041 50272 5051 50328
rect 4851 50204 5051 50272
rect 4851 50148 4861 50204
rect 4917 50148 4985 50204
rect 5041 50148 5051 50204
rect 4851 50080 5051 50148
rect 4851 50024 4861 50080
rect 4917 50024 4985 50080
rect 5041 50024 5051 50080
rect 4851 49956 5051 50024
rect 4851 49900 4861 49956
rect 4917 49900 4985 49956
rect 5041 49900 5051 49956
rect 4851 49832 5051 49900
rect 4851 49776 4861 49832
rect 4917 49776 4985 49832
rect 5041 49776 5051 49832
rect 4851 49751 5051 49776
rect 4851 49708 4871 49751
rect 4851 49652 4861 49708
rect 4923 49699 4979 49751
rect 5031 49708 5051 49751
rect 4917 49652 4985 49699
rect 5041 49652 5051 49708
rect 4851 49643 5051 49652
rect 4851 49591 4871 49643
rect 4923 49591 4979 49643
rect 5031 49591 5051 49643
rect 4851 48817 5051 49591
rect 4851 48765 4871 48817
rect 4923 48765 4979 48817
rect 5031 48765 5051 48817
rect 4851 48709 5051 48765
rect 4851 48657 4871 48709
rect 4923 48657 4979 48709
rect 5031 48657 5051 48709
rect 4851 47972 5051 48657
rect 4851 47920 4871 47972
rect 4923 47920 4979 47972
rect 5031 47920 5051 47972
rect 4851 47864 5051 47920
rect 4851 47812 4871 47864
rect 4923 47812 4979 47864
rect 5031 47812 5051 47864
rect 4851 47756 5051 47812
rect 4851 47704 4871 47756
rect 4923 47704 4979 47756
rect 5031 47704 5051 47756
rect 4851 46442 5051 47704
rect 5111 57104 7161 57600
rect 5111 57052 5138 57104
rect 5190 57052 5246 57104
rect 5298 57052 5354 57104
rect 5406 57052 5462 57104
rect 5514 57052 5570 57104
rect 5622 57052 5678 57104
rect 5730 57052 5786 57104
rect 5838 57052 5894 57104
rect 5946 57052 6002 57104
rect 6054 57052 6110 57104
rect 6162 57052 6218 57104
rect 6270 57052 6326 57104
rect 6378 57052 6434 57104
rect 6486 57052 6542 57104
rect 6594 57052 6650 57104
rect 6702 57052 6758 57104
rect 6810 57052 6866 57104
rect 6918 57052 6974 57104
rect 7026 57052 7082 57104
rect 7134 57052 7161 57104
rect 5111 53483 7161 57052
rect 5111 53431 5138 53483
rect 5190 53431 5246 53483
rect 5298 53431 5354 53483
rect 5406 53431 5462 53483
rect 5514 53431 5570 53483
rect 5622 53431 5678 53483
rect 5730 53431 5786 53483
rect 5838 53431 5894 53483
rect 5946 53431 6002 53483
rect 6054 53431 6110 53483
rect 6162 53431 6218 53483
rect 6270 53431 6326 53483
rect 6378 53431 6434 53483
rect 6486 53431 6542 53483
rect 6594 53431 6650 53483
rect 6702 53431 6758 53483
rect 6810 53431 6866 53483
rect 6918 53431 6974 53483
rect 7026 53431 7082 53483
rect 7134 53431 7161 53483
rect 5111 53375 7161 53431
rect 5111 53323 5138 53375
rect 5190 53323 5246 53375
rect 5298 53323 5354 53375
rect 5406 53323 5462 53375
rect 5514 53323 5570 53375
rect 5622 53323 5678 53375
rect 5730 53323 5786 53375
rect 5838 53323 5894 53375
rect 5946 53323 6002 53375
rect 6054 53323 6110 53375
rect 6162 53323 6218 53375
rect 6270 53323 6326 53375
rect 6378 53323 6434 53375
rect 6486 53323 6542 53375
rect 6594 53323 6650 53375
rect 6702 53323 6758 53375
rect 6810 53323 6866 53375
rect 6918 53323 6974 53375
rect 7026 53323 7082 53375
rect 7134 53323 7161 53375
rect 5111 53267 7161 53323
rect 5111 53215 5138 53267
rect 5190 53215 5246 53267
rect 5298 53215 5354 53267
rect 5406 53215 5462 53267
rect 5514 53215 5570 53267
rect 5622 53215 5678 53267
rect 5730 53215 5786 53267
rect 5838 53215 5894 53267
rect 5946 53215 6002 53267
rect 6054 53215 6110 53267
rect 6162 53215 6218 53267
rect 6270 53215 6326 53267
rect 6378 53215 6434 53267
rect 6486 53215 6542 53267
rect 6594 53215 6650 53267
rect 6702 53215 6758 53267
rect 6810 53215 6866 53267
rect 6918 53215 6974 53267
rect 7026 53215 7082 53267
rect 7134 53215 7161 53267
rect 5111 52548 7161 53215
rect 5111 52492 5178 52548
rect 5234 52492 5302 52548
rect 5358 52492 5426 52548
rect 5482 52492 5550 52548
rect 5606 52492 5674 52548
rect 5730 52492 5798 52548
rect 5854 52492 5922 52548
rect 5978 52492 6046 52548
rect 6102 52492 6170 52548
rect 6226 52492 6294 52548
rect 6350 52492 6418 52548
rect 6474 52492 6542 52548
rect 6598 52492 6666 52548
rect 6722 52492 6790 52548
rect 6846 52492 6914 52548
rect 6970 52492 7038 52548
rect 7094 52492 7161 52548
rect 5111 52424 7161 52492
rect 5111 52368 5178 52424
rect 5234 52368 5302 52424
rect 5358 52368 5426 52424
rect 5482 52368 5550 52424
rect 5606 52368 5674 52424
rect 5730 52368 5798 52424
rect 5854 52368 5922 52424
rect 5978 52368 6046 52424
rect 6102 52368 6170 52424
rect 6226 52368 6294 52424
rect 6350 52368 6418 52424
rect 6474 52368 6542 52424
rect 6598 52368 6666 52424
rect 6722 52368 6790 52424
rect 6846 52368 6914 52424
rect 6970 52368 7038 52424
rect 7094 52368 7161 52424
rect 5111 52300 7161 52368
rect 5111 52244 5178 52300
rect 5234 52244 5302 52300
rect 5358 52244 5426 52300
rect 5482 52244 5550 52300
rect 5606 52244 5674 52300
rect 5730 52244 5798 52300
rect 5854 52244 5922 52300
rect 5978 52244 6046 52300
rect 6102 52244 6170 52300
rect 6226 52244 6294 52300
rect 6350 52244 6418 52300
rect 6474 52244 6542 52300
rect 6598 52244 6666 52300
rect 6722 52244 6790 52300
rect 6846 52244 6914 52300
rect 6970 52244 7038 52300
rect 7094 52244 7161 52300
rect 5111 52176 7161 52244
rect 5111 52120 5178 52176
rect 5234 52120 5302 52176
rect 5358 52120 5426 52176
rect 5482 52120 5550 52176
rect 5606 52120 5674 52176
rect 5730 52120 5798 52176
rect 5854 52120 5922 52176
rect 5978 52120 6046 52176
rect 6102 52120 6170 52176
rect 6226 52120 6294 52176
rect 6350 52120 6418 52176
rect 6474 52120 6542 52176
rect 6598 52120 6666 52176
rect 6722 52120 6790 52176
rect 6846 52120 6914 52176
rect 6970 52120 7038 52176
rect 7094 52120 7161 52176
rect 5111 52052 7161 52120
rect 5111 52009 5178 52052
rect 5234 52009 5302 52052
rect 5358 52009 5426 52052
rect 5482 52009 5550 52052
rect 5606 52009 5674 52052
rect 5730 52009 5798 52052
rect 5854 52009 5922 52052
rect 5978 52009 6046 52052
rect 6102 52009 6170 52052
rect 6226 52009 6294 52052
rect 6350 52009 6418 52052
rect 6474 52009 6542 52052
rect 6598 52009 6666 52052
rect 6722 52009 6790 52052
rect 6846 52009 6914 52052
rect 6970 52009 7038 52052
rect 7094 52009 7161 52052
rect 5111 51957 5138 52009
rect 5234 51996 5246 52009
rect 5190 51957 5246 51996
rect 5298 51996 5302 52009
rect 5406 51996 5426 52009
rect 5514 51996 5550 52009
rect 5622 51996 5674 52009
rect 5298 51957 5354 51996
rect 5406 51957 5462 51996
rect 5514 51957 5570 51996
rect 5622 51957 5678 51996
rect 5730 51957 5786 52009
rect 5854 51996 5894 52009
rect 5978 51996 6002 52009
rect 6102 51996 6110 52009
rect 5838 51957 5894 51996
rect 5946 51957 6002 51996
rect 6054 51957 6110 51996
rect 6162 51996 6170 52009
rect 6270 51996 6294 52009
rect 6378 51996 6418 52009
rect 6162 51957 6218 51996
rect 6270 51957 6326 51996
rect 6378 51957 6434 51996
rect 6486 51957 6542 52009
rect 6598 51996 6650 52009
rect 6722 51996 6758 52009
rect 6846 51996 6866 52009
rect 6970 51996 6974 52009
rect 6594 51957 6650 51996
rect 6702 51957 6758 51996
rect 6810 51957 6866 51996
rect 6918 51957 6974 51996
rect 7026 51996 7038 52009
rect 7026 51957 7082 51996
rect 7134 51957 7161 52009
rect 5111 51928 7161 51957
rect 5111 51901 5178 51928
rect 5234 51901 5302 51928
rect 5358 51901 5426 51928
rect 5482 51901 5550 51928
rect 5606 51901 5674 51928
rect 5730 51901 5798 51928
rect 5854 51901 5922 51928
rect 5978 51901 6046 51928
rect 6102 51901 6170 51928
rect 6226 51901 6294 51928
rect 6350 51901 6418 51928
rect 6474 51901 6542 51928
rect 6598 51901 6666 51928
rect 6722 51901 6790 51928
rect 6846 51901 6914 51928
rect 6970 51901 7038 51928
rect 7094 51901 7161 51928
rect 5111 51849 5138 51901
rect 5234 51872 5246 51901
rect 5190 51849 5246 51872
rect 5298 51872 5302 51901
rect 5406 51872 5426 51901
rect 5514 51872 5550 51901
rect 5622 51872 5674 51901
rect 5298 51849 5354 51872
rect 5406 51849 5462 51872
rect 5514 51849 5570 51872
rect 5622 51849 5678 51872
rect 5730 51849 5786 51901
rect 5854 51872 5894 51901
rect 5978 51872 6002 51901
rect 6102 51872 6110 51901
rect 5838 51849 5894 51872
rect 5946 51849 6002 51872
rect 6054 51849 6110 51872
rect 6162 51872 6170 51901
rect 6270 51872 6294 51901
rect 6378 51872 6418 51901
rect 6162 51849 6218 51872
rect 6270 51849 6326 51872
rect 6378 51849 6434 51872
rect 6486 51849 6542 51901
rect 6598 51872 6650 51901
rect 6722 51872 6758 51901
rect 6846 51872 6866 51901
rect 6970 51872 6974 51901
rect 6594 51849 6650 51872
rect 6702 51849 6758 51872
rect 6810 51849 6866 51872
rect 6918 51849 6974 51872
rect 7026 51872 7038 51901
rect 7026 51849 7082 51872
rect 7134 51849 7161 51901
rect 5111 51804 7161 51849
rect 5111 51748 5178 51804
rect 5234 51748 5302 51804
rect 5358 51748 5426 51804
rect 5482 51748 5550 51804
rect 5606 51748 5674 51804
rect 5730 51748 5798 51804
rect 5854 51748 5922 51804
rect 5978 51748 6046 51804
rect 6102 51748 6170 51804
rect 6226 51748 6294 51804
rect 6350 51748 6418 51804
rect 6474 51748 6542 51804
rect 6598 51748 6666 51804
rect 6722 51748 6790 51804
rect 6846 51748 6914 51804
rect 6970 51748 7038 51804
rect 7094 51748 7161 51804
rect 5111 51680 7161 51748
rect 5111 51624 5178 51680
rect 5234 51624 5302 51680
rect 5358 51624 5426 51680
rect 5482 51624 5550 51680
rect 5606 51624 5674 51680
rect 5730 51624 5798 51680
rect 5854 51624 5922 51680
rect 5978 51624 6046 51680
rect 6102 51624 6170 51680
rect 6226 51624 6294 51680
rect 6350 51624 6418 51680
rect 6474 51624 6542 51680
rect 6598 51624 6666 51680
rect 6722 51624 6790 51680
rect 6846 51624 6914 51680
rect 6970 51624 7038 51680
rect 7094 51624 7161 51680
rect 5111 51556 7161 51624
rect 5111 51500 5178 51556
rect 5234 51500 5302 51556
rect 5358 51500 5426 51556
rect 5482 51500 5550 51556
rect 5606 51500 5674 51556
rect 5730 51500 5798 51556
rect 5854 51500 5922 51556
rect 5978 51500 6046 51556
rect 6102 51500 6170 51556
rect 6226 51500 6294 51556
rect 6350 51500 6418 51556
rect 6474 51500 6542 51556
rect 6598 51500 6666 51556
rect 6722 51500 6790 51556
rect 6846 51500 6914 51556
rect 6970 51500 7038 51556
rect 7094 51500 7161 51556
rect 5111 51432 7161 51500
rect 5111 51376 5178 51432
rect 5234 51376 5302 51432
rect 5358 51376 5426 51432
rect 5482 51376 5550 51432
rect 5606 51376 5674 51432
rect 5730 51376 5798 51432
rect 5854 51376 5922 51432
rect 5978 51376 6046 51432
rect 6102 51376 6170 51432
rect 6226 51376 6294 51432
rect 6350 51376 6418 51432
rect 6474 51376 6542 51432
rect 6598 51376 6666 51432
rect 6722 51376 6790 51432
rect 6846 51376 6914 51432
rect 6970 51376 7038 51432
rect 7094 51376 7161 51432
rect 5111 51308 7161 51376
rect 5111 51252 5178 51308
rect 5234 51252 5302 51308
rect 5358 51252 5426 51308
rect 5482 51252 5550 51308
rect 5606 51252 5674 51308
rect 5730 51252 5798 51308
rect 5854 51252 5922 51308
rect 5978 51252 6046 51308
rect 6102 51252 6170 51308
rect 6226 51252 6294 51308
rect 6350 51252 6418 51308
rect 6474 51252 6542 51308
rect 6598 51252 6666 51308
rect 6722 51252 6790 51308
rect 6846 51252 6914 51308
rect 6970 51252 7038 51308
rect 7094 51252 7161 51308
rect 5111 51206 7161 51252
rect 5111 51154 5138 51206
rect 5190 51154 5246 51206
rect 5298 51154 5354 51206
rect 5406 51154 5462 51206
rect 5514 51154 5570 51206
rect 5622 51154 5678 51206
rect 5730 51154 5786 51206
rect 5838 51154 5894 51206
rect 5946 51154 6002 51206
rect 6054 51154 6110 51206
rect 6162 51154 6218 51206
rect 6270 51154 6326 51206
rect 6378 51154 6434 51206
rect 6486 51154 6542 51206
rect 6594 51154 6650 51206
rect 6702 51154 6758 51206
rect 6810 51154 6866 51206
rect 6918 51154 6974 51206
rect 7026 51154 7082 51206
rect 7134 51154 7161 51206
rect 5111 51098 7161 51154
rect 5111 51046 5138 51098
rect 5190 51046 5246 51098
rect 5298 51046 5354 51098
rect 5406 51046 5462 51098
rect 5514 51046 5570 51098
rect 5622 51046 5678 51098
rect 5730 51046 5786 51098
rect 5838 51046 5894 51098
rect 5946 51046 6002 51098
rect 6054 51046 6110 51098
rect 6162 51046 6218 51098
rect 6270 51046 6326 51098
rect 6378 51046 6434 51098
rect 6486 51046 6542 51098
rect 6594 51046 6650 51098
rect 6702 51046 6758 51098
rect 6810 51046 6866 51098
rect 6918 51046 6974 51098
rect 7026 51046 7082 51098
rect 7134 51046 7161 51098
rect 5111 50990 7161 51046
rect 5111 50938 5138 50990
rect 5190 50938 5246 50990
rect 5298 50938 5354 50990
rect 5406 50938 5462 50990
rect 5514 50938 5570 50990
rect 5622 50938 5678 50990
rect 5730 50938 5786 50990
rect 5838 50938 5894 50990
rect 5946 50938 6002 50990
rect 6054 50938 6110 50990
rect 6162 50938 6218 50990
rect 6270 50938 6326 50990
rect 6378 50938 6434 50990
rect 6486 50938 6542 50990
rect 6594 50938 6650 50990
rect 6702 50938 6758 50990
rect 6810 50938 6866 50990
rect 6918 50938 6974 50990
rect 7026 50938 7082 50990
rect 7134 50938 7161 50990
rect 5111 50272 7161 50938
rect 5111 50220 5138 50272
rect 5190 50220 5246 50272
rect 5298 50220 5354 50272
rect 5406 50220 5462 50272
rect 5514 50220 5570 50272
rect 5622 50220 5678 50272
rect 5730 50220 5786 50272
rect 5838 50220 5894 50272
rect 5946 50220 6002 50272
rect 6054 50220 6110 50272
rect 6162 50220 6218 50272
rect 6270 50220 6326 50272
rect 6378 50220 6434 50272
rect 6486 50220 6542 50272
rect 6594 50220 6650 50272
rect 6702 50220 6758 50272
rect 6810 50220 6866 50272
rect 6918 50220 6974 50272
rect 7026 50220 7082 50272
rect 7134 50220 7161 50272
rect 5111 50164 7161 50220
rect 5111 50112 5138 50164
rect 5190 50112 5246 50164
rect 5298 50112 5354 50164
rect 5406 50112 5462 50164
rect 5514 50112 5570 50164
rect 5622 50112 5678 50164
rect 5730 50112 5786 50164
rect 5838 50112 5894 50164
rect 5946 50112 6002 50164
rect 6054 50112 6110 50164
rect 6162 50112 6218 50164
rect 6270 50112 6326 50164
rect 6378 50112 6434 50164
rect 6486 50112 6542 50164
rect 6594 50112 6650 50164
rect 6702 50112 6758 50164
rect 6810 50112 6866 50164
rect 6918 50112 6974 50164
rect 7026 50112 7082 50164
rect 7134 50112 7161 50164
rect 5111 50056 7161 50112
rect 5111 50004 5138 50056
rect 5190 50004 5246 50056
rect 5298 50004 5354 50056
rect 5406 50004 5462 50056
rect 5514 50004 5570 50056
rect 5622 50004 5678 50056
rect 5730 50004 5786 50056
rect 5838 50004 5894 50056
rect 5946 50004 6002 50056
rect 6054 50004 6110 50056
rect 6162 50004 6218 50056
rect 6270 50004 6326 50056
rect 6378 50004 6434 50056
rect 6486 50004 6542 50056
rect 6594 50004 6650 50056
rect 6702 50004 6758 50056
rect 6810 50004 6866 50056
rect 6918 50004 6974 50056
rect 7026 50004 7082 50056
rect 7134 50004 7161 50056
rect 5111 49338 7161 50004
rect 5111 49286 5138 49338
rect 5190 49286 5246 49338
rect 5298 49286 5354 49338
rect 5406 49286 5462 49338
rect 5514 49286 5570 49338
rect 5622 49286 5678 49338
rect 5730 49286 5786 49338
rect 5838 49286 5894 49338
rect 5946 49286 6002 49338
rect 6054 49286 6110 49338
rect 6162 49286 6218 49338
rect 6270 49286 6326 49338
rect 6378 49286 6434 49338
rect 6486 49286 6542 49338
rect 6594 49286 6650 49338
rect 6702 49286 6758 49338
rect 6810 49286 6866 49338
rect 6918 49286 6974 49338
rect 7026 49286 7082 49338
rect 7134 49286 7161 49338
rect 5111 49230 7161 49286
rect 5111 49178 5138 49230
rect 5190 49178 5246 49230
rect 5298 49178 5354 49230
rect 5406 49178 5462 49230
rect 5514 49178 5570 49230
rect 5622 49178 5678 49230
rect 5730 49178 5786 49230
rect 5838 49178 5894 49230
rect 5946 49178 6002 49230
rect 6054 49178 6110 49230
rect 6162 49178 6218 49230
rect 6270 49178 6326 49230
rect 6378 49178 6434 49230
rect 6486 49178 6542 49230
rect 6594 49178 6650 49230
rect 6702 49178 6758 49230
rect 6810 49178 6866 49230
rect 6918 49178 6974 49230
rect 7026 49178 7082 49230
rect 7134 49178 7161 49230
rect 5111 49122 7161 49178
rect 5111 49070 5138 49122
rect 5190 49070 5246 49122
rect 5298 49070 5354 49122
rect 5406 49070 5462 49122
rect 5514 49070 5570 49122
rect 5622 49070 5678 49122
rect 5730 49070 5786 49122
rect 5838 49070 5894 49122
rect 5946 49070 6002 49122
rect 6054 49070 6110 49122
rect 6162 49070 6218 49122
rect 6270 49070 6326 49122
rect 6378 49070 6434 49122
rect 6486 49070 6542 49122
rect 6594 49070 6650 49122
rect 6702 49070 6758 49122
rect 6810 49070 6866 49122
rect 6918 49070 6974 49122
rect 7026 49070 7082 49122
rect 7134 49070 7161 49122
rect 5111 48427 7161 49070
rect 5111 48375 5138 48427
rect 5190 48375 5246 48427
rect 5298 48375 5354 48427
rect 5406 48375 5462 48427
rect 5514 48375 5570 48427
rect 5622 48375 5678 48427
rect 5730 48375 5786 48427
rect 5838 48375 5894 48427
rect 5946 48375 6002 48427
rect 6054 48375 6110 48427
rect 6162 48375 6218 48427
rect 6270 48375 6326 48427
rect 6378 48375 6434 48427
rect 6486 48375 6542 48427
rect 6594 48375 6650 48427
rect 6702 48375 6758 48427
rect 6810 48375 6866 48427
rect 6918 48375 6974 48427
rect 7026 48375 7082 48427
rect 7134 48375 7161 48427
rect 5111 48319 7161 48375
rect 5111 48267 5138 48319
rect 5190 48267 5246 48319
rect 5298 48267 5354 48319
rect 5406 48267 5462 48319
rect 5514 48267 5570 48319
rect 5622 48267 5678 48319
rect 5730 48267 5786 48319
rect 5838 48267 5894 48319
rect 5946 48267 6002 48319
rect 6054 48267 6110 48319
rect 6162 48267 6218 48319
rect 6270 48267 6326 48319
rect 6378 48267 6434 48319
rect 6486 48267 6542 48319
rect 6594 48267 6650 48319
rect 6702 48267 6758 48319
rect 6810 48267 6866 48319
rect 6918 48267 6974 48319
rect 7026 48267 7082 48319
rect 7134 48267 7161 48319
rect 5111 47163 7161 48267
rect 7221 52572 7757 57278
rect 7221 52520 7247 52572
rect 7299 52520 7355 52572
rect 7407 52520 7463 52572
rect 7515 52520 7571 52572
rect 7623 52520 7679 52572
rect 7731 52520 7757 52572
rect 7221 52464 7757 52520
rect 7221 52412 7247 52464
rect 7299 52412 7355 52464
rect 7407 52412 7463 52464
rect 7515 52412 7571 52464
rect 7623 52412 7679 52464
rect 7731 52412 7757 52464
rect 7221 52356 7757 52412
rect 7221 52304 7247 52356
rect 7299 52304 7355 52356
rect 7407 52304 7463 52356
rect 7515 52304 7571 52356
rect 7623 52304 7679 52356
rect 7731 52304 7757 52356
rect 7221 51619 7757 52304
rect 7221 51567 7247 51619
rect 7299 51567 7355 51619
rect 7407 51567 7463 51619
rect 7515 51567 7571 51619
rect 7623 51567 7679 51619
rect 7731 51567 7757 51619
rect 7221 51511 7757 51567
rect 7221 51459 7247 51511
rect 7299 51459 7355 51511
rect 7407 51459 7463 51511
rect 7515 51459 7571 51511
rect 7623 51459 7679 51511
rect 7731 51459 7757 51511
rect 7221 50948 7757 51459
rect 7221 50892 7275 50948
rect 7331 50892 7399 50948
rect 7455 50892 7523 50948
rect 7579 50892 7647 50948
rect 7703 50892 7757 50948
rect 7221 50824 7757 50892
rect 7221 50768 7275 50824
rect 7331 50768 7399 50824
rect 7455 50768 7523 50824
rect 7579 50768 7647 50824
rect 7703 50768 7757 50824
rect 7221 50700 7757 50768
rect 7221 50685 7275 50700
rect 7331 50685 7399 50700
rect 7455 50685 7523 50700
rect 7579 50685 7647 50700
rect 7703 50685 7757 50700
rect 7221 50633 7247 50685
rect 7331 50644 7355 50685
rect 7455 50644 7463 50685
rect 7299 50633 7355 50644
rect 7407 50633 7463 50644
rect 7515 50644 7523 50685
rect 7623 50644 7647 50685
rect 7515 50633 7571 50644
rect 7623 50633 7679 50644
rect 7731 50633 7757 50685
rect 7221 50577 7757 50633
rect 7221 50525 7247 50577
rect 7299 50576 7355 50577
rect 7407 50576 7463 50577
rect 7331 50525 7355 50576
rect 7455 50525 7463 50576
rect 7515 50576 7571 50577
rect 7623 50576 7679 50577
rect 7515 50525 7523 50576
rect 7623 50525 7647 50576
rect 7731 50525 7757 50577
rect 7221 50520 7275 50525
rect 7331 50520 7399 50525
rect 7455 50520 7523 50525
rect 7579 50520 7647 50525
rect 7703 50520 7757 50525
rect 7221 50452 7757 50520
rect 7221 50396 7275 50452
rect 7331 50396 7399 50452
rect 7455 50396 7523 50452
rect 7579 50396 7647 50452
rect 7703 50396 7757 50452
rect 7221 50328 7757 50396
rect 7221 50272 7275 50328
rect 7331 50272 7399 50328
rect 7455 50272 7523 50328
rect 7579 50272 7647 50328
rect 7703 50272 7757 50328
rect 7221 50204 7757 50272
rect 7221 50148 7275 50204
rect 7331 50148 7399 50204
rect 7455 50148 7523 50204
rect 7579 50148 7647 50204
rect 7703 50148 7757 50204
rect 7221 50080 7757 50148
rect 7221 50024 7275 50080
rect 7331 50024 7399 50080
rect 7455 50024 7523 50080
rect 7579 50024 7647 50080
rect 7703 50024 7757 50080
rect 7221 49956 7757 50024
rect 7221 49900 7275 49956
rect 7331 49900 7399 49956
rect 7455 49900 7523 49956
rect 7579 49900 7647 49956
rect 7703 49900 7757 49956
rect 7221 49832 7757 49900
rect 7221 49776 7275 49832
rect 7331 49776 7399 49832
rect 7455 49776 7523 49832
rect 7579 49776 7647 49832
rect 7703 49776 7757 49832
rect 7221 49751 7757 49776
rect 7221 49699 7247 49751
rect 7299 49708 7355 49751
rect 7407 49708 7463 49751
rect 7331 49699 7355 49708
rect 7455 49699 7463 49708
rect 7515 49708 7571 49751
rect 7623 49708 7679 49751
rect 7515 49699 7523 49708
rect 7623 49699 7647 49708
rect 7731 49699 7757 49751
rect 7221 49652 7275 49699
rect 7331 49652 7399 49699
rect 7455 49652 7523 49699
rect 7579 49652 7647 49699
rect 7703 49652 7757 49699
rect 7221 49643 7757 49652
rect 7221 49591 7247 49643
rect 7299 49591 7355 49643
rect 7407 49591 7463 49643
rect 7515 49591 7571 49643
rect 7623 49591 7679 49643
rect 7731 49591 7757 49643
rect 7221 48817 7757 49591
rect 7221 48765 7247 48817
rect 7299 48765 7355 48817
rect 7407 48765 7463 48817
rect 7515 48765 7571 48817
rect 7623 48765 7679 48817
rect 7731 48765 7757 48817
rect 7221 48709 7757 48765
rect 7221 48657 7247 48709
rect 7299 48657 7355 48709
rect 7407 48657 7463 48709
rect 7515 48657 7571 48709
rect 7623 48657 7679 48709
rect 7731 48657 7757 48709
rect 7221 47972 7757 48657
rect 7221 47920 7247 47972
rect 7299 47920 7355 47972
rect 7407 47920 7463 47972
rect 7515 47920 7571 47972
rect 7623 47920 7679 47972
rect 7731 47920 7757 47972
rect 7221 47864 7757 47920
rect 7221 47812 7247 47864
rect 7299 47812 7355 47864
rect 7407 47812 7463 47864
rect 7515 47812 7571 47864
rect 7623 47812 7679 47864
rect 7731 47812 7757 47864
rect 7221 47756 7757 47812
rect 7221 47704 7247 47756
rect 7299 47704 7355 47756
rect 7407 47704 7463 47756
rect 7515 47704 7571 47756
rect 7623 47704 7679 47756
rect 7731 47704 7757 47756
rect 7221 47163 7757 47704
rect 7817 57104 9867 57600
rect 7817 57052 7844 57104
rect 7896 57052 7952 57104
rect 8004 57052 8060 57104
rect 8112 57052 8168 57104
rect 8220 57052 8276 57104
rect 8328 57052 8384 57104
rect 8436 57052 8492 57104
rect 8544 57052 8600 57104
rect 8652 57052 8708 57104
rect 8760 57052 8816 57104
rect 8868 57052 8924 57104
rect 8976 57052 9032 57104
rect 9084 57052 9140 57104
rect 9192 57052 9248 57104
rect 9300 57052 9356 57104
rect 9408 57052 9464 57104
rect 9516 57052 9572 57104
rect 9624 57052 9680 57104
rect 9732 57052 9788 57104
rect 9840 57052 9867 57104
rect 7817 53483 9867 57052
rect 7817 53431 7844 53483
rect 7896 53431 7952 53483
rect 8004 53431 8060 53483
rect 8112 53431 8168 53483
rect 8220 53431 8276 53483
rect 8328 53431 8384 53483
rect 8436 53431 8492 53483
rect 8544 53431 8600 53483
rect 8652 53431 8708 53483
rect 8760 53431 8816 53483
rect 8868 53431 8924 53483
rect 8976 53431 9032 53483
rect 9084 53431 9140 53483
rect 9192 53431 9248 53483
rect 9300 53431 9356 53483
rect 9408 53431 9464 53483
rect 9516 53431 9572 53483
rect 9624 53431 9680 53483
rect 9732 53431 9788 53483
rect 9840 53431 9867 53483
rect 7817 53375 9867 53431
rect 7817 53323 7844 53375
rect 7896 53323 7952 53375
rect 8004 53323 8060 53375
rect 8112 53323 8168 53375
rect 8220 53323 8276 53375
rect 8328 53323 8384 53375
rect 8436 53323 8492 53375
rect 8544 53323 8600 53375
rect 8652 53323 8708 53375
rect 8760 53323 8816 53375
rect 8868 53323 8924 53375
rect 8976 53323 9032 53375
rect 9084 53323 9140 53375
rect 9192 53323 9248 53375
rect 9300 53323 9356 53375
rect 9408 53323 9464 53375
rect 9516 53323 9572 53375
rect 9624 53323 9680 53375
rect 9732 53323 9788 53375
rect 9840 53323 9867 53375
rect 7817 53267 9867 53323
rect 7817 53215 7844 53267
rect 7896 53215 7952 53267
rect 8004 53215 8060 53267
rect 8112 53215 8168 53267
rect 8220 53215 8276 53267
rect 8328 53215 8384 53267
rect 8436 53215 8492 53267
rect 8544 53215 8600 53267
rect 8652 53215 8708 53267
rect 8760 53215 8816 53267
rect 8868 53215 8924 53267
rect 8976 53215 9032 53267
rect 9084 53215 9140 53267
rect 9192 53215 9248 53267
rect 9300 53215 9356 53267
rect 9408 53215 9464 53267
rect 9516 53215 9572 53267
rect 9624 53215 9680 53267
rect 9732 53215 9788 53267
rect 9840 53215 9867 53267
rect 7817 52548 9867 53215
rect 7817 52492 7884 52548
rect 7940 52492 8008 52548
rect 8064 52492 8132 52548
rect 8188 52492 8256 52548
rect 8312 52492 8380 52548
rect 8436 52492 8504 52548
rect 8560 52492 8628 52548
rect 8684 52492 8752 52548
rect 8808 52492 8876 52548
rect 8932 52492 9000 52548
rect 9056 52492 9124 52548
rect 9180 52492 9248 52548
rect 9304 52492 9372 52548
rect 9428 52492 9496 52548
rect 9552 52492 9620 52548
rect 9676 52492 9744 52548
rect 9800 52492 9867 52548
rect 7817 52424 9867 52492
rect 7817 52368 7884 52424
rect 7940 52368 8008 52424
rect 8064 52368 8132 52424
rect 8188 52368 8256 52424
rect 8312 52368 8380 52424
rect 8436 52368 8504 52424
rect 8560 52368 8628 52424
rect 8684 52368 8752 52424
rect 8808 52368 8876 52424
rect 8932 52368 9000 52424
rect 9056 52368 9124 52424
rect 9180 52368 9248 52424
rect 9304 52368 9372 52424
rect 9428 52368 9496 52424
rect 9552 52368 9620 52424
rect 9676 52368 9744 52424
rect 9800 52368 9867 52424
rect 7817 52300 9867 52368
rect 7817 52244 7884 52300
rect 7940 52244 8008 52300
rect 8064 52244 8132 52300
rect 8188 52244 8256 52300
rect 8312 52244 8380 52300
rect 8436 52244 8504 52300
rect 8560 52244 8628 52300
rect 8684 52244 8752 52300
rect 8808 52244 8876 52300
rect 8932 52244 9000 52300
rect 9056 52244 9124 52300
rect 9180 52244 9248 52300
rect 9304 52244 9372 52300
rect 9428 52244 9496 52300
rect 9552 52244 9620 52300
rect 9676 52244 9744 52300
rect 9800 52244 9867 52300
rect 7817 52176 9867 52244
rect 7817 52120 7884 52176
rect 7940 52120 8008 52176
rect 8064 52120 8132 52176
rect 8188 52120 8256 52176
rect 8312 52120 8380 52176
rect 8436 52120 8504 52176
rect 8560 52120 8628 52176
rect 8684 52120 8752 52176
rect 8808 52120 8876 52176
rect 8932 52120 9000 52176
rect 9056 52120 9124 52176
rect 9180 52120 9248 52176
rect 9304 52120 9372 52176
rect 9428 52120 9496 52176
rect 9552 52120 9620 52176
rect 9676 52120 9744 52176
rect 9800 52120 9867 52176
rect 7817 52052 9867 52120
rect 7817 52009 7884 52052
rect 7940 52009 8008 52052
rect 8064 52009 8132 52052
rect 8188 52009 8256 52052
rect 8312 52009 8380 52052
rect 8436 52009 8504 52052
rect 8560 52009 8628 52052
rect 8684 52009 8752 52052
rect 8808 52009 8876 52052
rect 8932 52009 9000 52052
rect 9056 52009 9124 52052
rect 9180 52009 9248 52052
rect 9304 52009 9372 52052
rect 9428 52009 9496 52052
rect 9552 52009 9620 52052
rect 9676 52009 9744 52052
rect 9800 52009 9867 52052
rect 7817 51957 7844 52009
rect 7940 51996 7952 52009
rect 7896 51957 7952 51996
rect 8004 51996 8008 52009
rect 8112 51996 8132 52009
rect 8220 51996 8256 52009
rect 8328 51996 8380 52009
rect 8004 51957 8060 51996
rect 8112 51957 8168 51996
rect 8220 51957 8276 51996
rect 8328 51957 8384 51996
rect 8436 51957 8492 52009
rect 8560 51996 8600 52009
rect 8684 51996 8708 52009
rect 8808 51996 8816 52009
rect 8544 51957 8600 51996
rect 8652 51957 8708 51996
rect 8760 51957 8816 51996
rect 8868 51996 8876 52009
rect 8976 51996 9000 52009
rect 9084 51996 9124 52009
rect 8868 51957 8924 51996
rect 8976 51957 9032 51996
rect 9084 51957 9140 51996
rect 9192 51957 9248 52009
rect 9304 51996 9356 52009
rect 9428 51996 9464 52009
rect 9552 51996 9572 52009
rect 9676 51996 9680 52009
rect 9300 51957 9356 51996
rect 9408 51957 9464 51996
rect 9516 51957 9572 51996
rect 9624 51957 9680 51996
rect 9732 51996 9744 52009
rect 9732 51957 9788 51996
rect 9840 51957 9867 52009
rect 7817 51928 9867 51957
rect 7817 51901 7884 51928
rect 7940 51901 8008 51928
rect 8064 51901 8132 51928
rect 8188 51901 8256 51928
rect 8312 51901 8380 51928
rect 8436 51901 8504 51928
rect 8560 51901 8628 51928
rect 8684 51901 8752 51928
rect 8808 51901 8876 51928
rect 8932 51901 9000 51928
rect 9056 51901 9124 51928
rect 9180 51901 9248 51928
rect 9304 51901 9372 51928
rect 9428 51901 9496 51928
rect 9552 51901 9620 51928
rect 9676 51901 9744 51928
rect 9800 51901 9867 51928
rect 7817 51849 7844 51901
rect 7940 51872 7952 51901
rect 7896 51849 7952 51872
rect 8004 51872 8008 51901
rect 8112 51872 8132 51901
rect 8220 51872 8256 51901
rect 8328 51872 8380 51901
rect 8004 51849 8060 51872
rect 8112 51849 8168 51872
rect 8220 51849 8276 51872
rect 8328 51849 8384 51872
rect 8436 51849 8492 51901
rect 8560 51872 8600 51901
rect 8684 51872 8708 51901
rect 8808 51872 8816 51901
rect 8544 51849 8600 51872
rect 8652 51849 8708 51872
rect 8760 51849 8816 51872
rect 8868 51872 8876 51901
rect 8976 51872 9000 51901
rect 9084 51872 9124 51901
rect 8868 51849 8924 51872
rect 8976 51849 9032 51872
rect 9084 51849 9140 51872
rect 9192 51849 9248 51901
rect 9304 51872 9356 51901
rect 9428 51872 9464 51901
rect 9552 51872 9572 51901
rect 9676 51872 9680 51901
rect 9300 51849 9356 51872
rect 9408 51849 9464 51872
rect 9516 51849 9572 51872
rect 9624 51849 9680 51872
rect 9732 51872 9744 51901
rect 9732 51849 9788 51872
rect 9840 51849 9867 51901
rect 7817 51804 9867 51849
rect 7817 51748 7884 51804
rect 7940 51748 8008 51804
rect 8064 51748 8132 51804
rect 8188 51748 8256 51804
rect 8312 51748 8380 51804
rect 8436 51748 8504 51804
rect 8560 51748 8628 51804
rect 8684 51748 8752 51804
rect 8808 51748 8876 51804
rect 8932 51748 9000 51804
rect 9056 51748 9124 51804
rect 9180 51748 9248 51804
rect 9304 51748 9372 51804
rect 9428 51748 9496 51804
rect 9552 51748 9620 51804
rect 9676 51748 9744 51804
rect 9800 51748 9867 51804
rect 7817 51680 9867 51748
rect 7817 51624 7884 51680
rect 7940 51624 8008 51680
rect 8064 51624 8132 51680
rect 8188 51624 8256 51680
rect 8312 51624 8380 51680
rect 8436 51624 8504 51680
rect 8560 51624 8628 51680
rect 8684 51624 8752 51680
rect 8808 51624 8876 51680
rect 8932 51624 9000 51680
rect 9056 51624 9124 51680
rect 9180 51624 9248 51680
rect 9304 51624 9372 51680
rect 9428 51624 9496 51680
rect 9552 51624 9620 51680
rect 9676 51624 9744 51680
rect 9800 51624 9867 51680
rect 7817 51556 9867 51624
rect 7817 51500 7884 51556
rect 7940 51500 8008 51556
rect 8064 51500 8132 51556
rect 8188 51500 8256 51556
rect 8312 51500 8380 51556
rect 8436 51500 8504 51556
rect 8560 51500 8628 51556
rect 8684 51500 8752 51556
rect 8808 51500 8876 51556
rect 8932 51500 9000 51556
rect 9056 51500 9124 51556
rect 9180 51500 9248 51556
rect 9304 51500 9372 51556
rect 9428 51500 9496 51556
rect 9552 51500 9620 51556
rect 9676 51500 9744 51556
rect 9800 51500 9867 51556
rect 7817 51432 9867 51500
rect 7817 51376 7884 51432
rect 7940 51376 8008 51432
rect 8064 51376 8132 51432
rect 8188 51376 8256 51432
rect 8312 51376 8380 51432
rect 8436 51376 8504 51432
rect 8560 51376 8628 51432
rect 8684 51376 8752 51432
rect 8808 51376 8876 51432
rect 8932 51376 9000 51432
rect 9056 51376 9124 51432
rect 9180 51376 9248 51432
rect 9304 51376 9372 51432
rect 9428 51376 9496 51432
rect 9552 51376 9620 51432
rect 9676 51376 9744 51432
rect 9800 51376 9867 51432
rect 7817 51308 9867 51376
rect 7817 51252 7884 51308
rect 7940 51252 8008 51308
rect 8064 51252 8132 51308
rect 8188 51252 8256 51308
rect 8312 51252 8380 51308
rect 8436 51252 8504 51308
rect 8560 51252 8628 51308
rect 8684 51252 8752 51308
rect 8808 51252 8876 51308
rect 8932 51252 9000 51308
rect 9056 51252 9124 51308
rect 9180 51252 9248 51308
rect 9304 51252 9372 51308
rect 9428 51252 9496 51308
rect 9552 51252 9620 51308
rect 9676 51252 9744 51308
rect 9800 51252 9867 51308
rect 7817 51206 9867 51252
rect 7817 51154 7844 51206
rect 7896 51154 7952 51206
rect 8004 51154 8060 51206
rect 8112 51154 8168 51206
rect 8220 51154 8276 51206
rect 8328 51154 8384 51206
rect 8436 51154 8492 51206
rect 8544 51154 8600 51206
rect 8652 51154 8708 51206
rect 8760 51154 8816 51206
rect 8868 51154 8924 51206
rect 8976 51154 9032 51206
rect 9084 51154 9140 51206
rect 9192 51154 9248 51206
rect 9300 51154 9356 51206
rect 9408 51154 9464 51206
rect 9516 51154 9572 51206
rect 9624 51154 9680 51206
rect 9732 51154 9788 51206
rect 9840 51154 9867 51206
rect 7817 51098 9867 51154
rect 7817 51046 7844 51098
rect 7896 51046 7952 51098
rect 8004 51046 8060 51098
rect 8112 51046 8168 51098
rect 8220 51046 8276 51098
rect 8328 51046 8384 51098
rect 8436 51046 8492 51098
rect 8544 51046 8600 51098
rect 8652 51046 8708 51098
rect 8760 51046 8816 51098
rect 8868 51046 8924 51098
rect 8976 51046 9032 51098
rect 9084 51046 9140 51098
rect 9192 51046 9248 51098
rect 9300 51046 9356 51098
rect 9408 51046 9464 51098
rect 9516 51046 9572 51098
rect 9624 51046 9680 51098
rect 9732 51046 9788 51098
rect 9840 51046 9867 51098
rect 7817 50990 9867 51046
rect 7817 50938 7844 50990
rect 7896 50938 7952 50990
rect 8004 50938 8060 50990
rect 8112 50938 8168 50990
rect 8220 50938 8276 50990
rect 8328 50938 8384 50990
rect 8436 50938 8492 50990
rect 8544 50938 8600 50990
rect 8652 50938 8708 50990
rect 8760 50938 8816 50990
rect 8868 50938 8924 50990
rect 8976 50938 9032 50990
rect 9084 50938 9140 50990
rect 9192 50938 9248 50990
rect 9300 50938 9356 50990
rect 9408 50938 9464 50990
rect 9516 50938 9572 50990
rect 9624 50938 9680 50990
rect 9732 50938 9788 50990
rect 9840 50938 9867 50990
rect 7817 50272 9867 50938
rect 7817 50220 7844 50272
rect 7896 50220 7952 50272
rect 8004 50220 8060 50272
rect 8112 50220 8168 50272
rect 8220 50220 8276 50272
rect 8328 50220 8384 50272
rect 8436 50220 8492 50272
rect 8544 50220 8600 50272
rect 8652 50220 8708 50272
rect 8760 50220 8816 50272
rect 8868 50220 8924 50272
rect 8976 50220 9032 50272
rect 9084 50220 9140 50272
rect 9192 50220 9248 50272
rect 9300 50220 9356 50272
rect 9408 50220 9464 50272
rect 9516 50220 9572 50272
rect 9624 50220 9680 50272
rect 9732 50220 9788 50272
rect 9840 50220 9867 50272
rect 7817 50164 9867 50220
rect 7817 50112 7844 50164
rect 7896 50112 7952 50164
rect 8004 50112 8060 50164
rect 8112 50112 8168 50164
rect 8220 50112 8276 50164
rect 8328 50112 8384 50164
rect 8436 50112 8492 50164
rect 8544 50112 8600 50164
rect 8652 50112 8708 50164
rect 8760 50112 8816 50164
rect 8868 50112 8924 50164
rect 8976 50112 9032 50164
rect 9084 50112 9140 50164
rect 9192 50112 9248 50164
rect 9300 50112 9356 50164
rect 9408 50112 9464 50164
rect 9516 50112 9572 50164
rect 9624 50112 9680 50164
rect 9732 50112 9788 50164
rect 9840 50112 9867 50164
rect 7817 50056 9867 50112
rect 7817 50004 7844 50056
rect 7896 50004 7952 50056
rect 8004 50004 8060 50056
rect 8112 50004 8168 50056
rect 8220 50004 8276 50056
rect 8328 50004 8384 50056
rect 8436 50004 8492 50056
rect 8544 50004 8600 50056
rect 8652 50004 8708 50056
rect 8760 50004 8816 50056
rect 8868 50004 8924 50056
rect 8976 50004 9032 50056
rect 9084 50004 9140 50056
rect 9192 50004 9248 50056
rect 9300 50004 9356 50056
rect 9408 50004 9464 50056
rect 9516 50004 9572 50056
rect 9624 50004 9680 50056
rect 9732 50004 9788 50056
rect 9840 50004 9867 50056
rect 7817 49338 9867 50004
rect 7817 49286 7844 49338
rect 7896 49286 7952 49338
rect 8004 49286 8060 49338
rect 8112 49286 8168 49338
rect 8220 49286 8276 49338
rect 8328 49286 8384 49338
rect 8436 49286 8492 49338
rect 8544 49286 8600 49338
rect 8652 49286 8708 49338
rect 8760 49286 8816 49338
rect 8868 49286 8924 49338
rect 8976 49286 9032 49338
rect 9084 49286 9140 49338
rect 9192 49286 9248 49338
rect 9300 49286 9356 49338
rect 9408 49286 9464 49338
rect 9516 49286 9572 49338
rect 9624 49286 9680 49338
rect 9732 49286 9788 49338
rect 9840 49286 9867 49338
rect 7817 49230 9867 49286
rect 7817 49178 7844 49230
rect 7896 49178 7952 49230
rect 8004 49178 8060 49230
rect 8112 49178 8168 49230
rect 8220 49178 8276 49230
rect 8328 49178 8384 49230
rect 8436 49178 8492 49230
rect 8544 49178 8600 49230
rect 8652 49178 8708 49230
rect 8760 49178 8816 49230
rect 8868 49178 8924 49230
rect 8976 49178 9032 49230
rect 9084 49178 9140 49230
rect 9192 49178 9248 49230
rect 9300 49178 9356 49230
rect 9408 49178 9464 49230
rect 9516 49178 9572 49230
rect 9624 49178 9680 49230
rect 9732 49178 9788 49230
rect 9840 49178 9867 49230
rect 7817 49122 9867 49178
rect 7817 49070 7844 49122
rect 7896 49070 7952 49122
rect 8004 49070 8060 49122
rect 8112 49070 8168 49122
rect 8220 49070 8276 49122
rect 8328 49070 8384 49122
rect 8436 49070 8492 49122
rect 8544 49070 8600 49122
rect 8652 49070 8708 49122
rect 8760 49070 8816 49122
rect 8868 49070 8924 49122
rect 8976 49070 9032 49122
rect 9084 49070 9140 49122
rect 9192 49070 9248 49122
rect 9300 49070 9356 49122
rect 9408 49070 9464 49122
rect 9516 49070 9572 49122
rect 9624 49070 9680 49122
rect 9732 49070 9788 49122
rect 9840 49070 9867 49122
rect 7817 48427 9867 49070
rect 7817 48375 7844 48427
rect 7896 48375 7952 48427
rect 8004 48375 8060 48427
rect 8112 48375 8168 48427
rect 8220 48375 8276 48427
rect 8328 48375 8384 48427
rect 8436 48375 8492 48427
rect 8544 48375 8600 48427
rect 8652 48375 8708 48427
rect 8760 48375 8816 48427
rect 8868 48375 8924 48427
rect 8976 48375 9032 48427
rect 9084 48375 9140 48427
rect 9192 48375 9248 48427
rect 9300 48375 9356 48427
rect 9408 48375 9464 48427
rect 9516 48375 9572 48427
rect 9624 48375 9680 48427
rect 9732 48375 9788 48427
rect 9840 48375 9867 48427
rect 7817 48319 9867 48375
rect 7817 48267 7844 48319
rect 7896 48267 7952 48319
rect 8004 48267 8060 48319
rect 8112 48267 8168 48319
rect 8220 48267 8276 48319
rect 8328 48267 8384 48319
rect 8436 48267 8492 48319
rect 8544 48267 8600 48319
rect 8652 48267 8708 48319
rect 8760 48267 8816 48319
rect 8868 48267 8924 48319
rect 8976 48267 9032 48319
rect 9084 48267 9140 48319
rect 9192 48267 9248 48319
rect 9300 48267 9356 48319
rect 9408 48267 9464 48319
rect 9516 48267 9572 48319
rect 9624 48267 9680 48319
rect 9732 48267 9788 48319
rect 9840 48267 9867 48319
rect 7817 47163 9867 48267
rect 9927 56693 10127 57278
rect 9927 56641 9947 56693
rect 9999 56641 10055 56693
rect 10107 56641 10127 56693
rect 9927 56585 10127 56641
rect 9927 56533 9947 56585
rect 9999 56533 10055 56585
rect 10107 56533 10127 56585
rect 9927 56477 10127 56533
rect 9927 56425 9947 56477
rect 9999 56425 10055 56477
rect 10107 56425 10127 56477
rect 9927 56369 10127 56425
rect 9927 56317 9947 56369
rect 9999 56317 10055 56369
rect 10107 56317 10127 56369
rect 9927 56261 10127 56317
rect 9927 56209 9947 56261
rect 9999 56209 10055 56261
rect 10107 56209 10127 56261
rect 9927 56153 10127 56209
rect 9927 56101 9947 56153
rect 9999 56101 10055 56153
rect 10107 56101 10127 56153
rect 9927 56045 10127 56101
rect 9927 55993 9947 56045
rect 9999 55993 10055 56045
rect 10107 55993 10127 56045
rect 9927 55937 10127 55993
rect 9927 55885 9947 55937
rect 9999 55885 10055 55937
rect 10107 55885 10127 55937
rect 9927 55829 10127 55885
rect 9927 55777 9947 55829
rect 9999 55777 10055 55829
rect 10107 55777 10127 55829
rect 9927 55721 10127 55777
rect 9927 55669 9947 55721
rect 9999 55669 10055 55721
rect 10107 55669 10127 55721
rect 9927 55613 10127 55669
rect 9927 55561 9947 55613
rect 9999 55561 10055 55613
rect 10107 55561 10127 55613
rect 9927 55505 10127 55561
rect 9927 55453 9947 55505
rect 9999 55453 10055 55505
rect 10107 55453 10127 55505
rect 9927 55397 10127 55453
rect 9927 55345 9947 55397
rect 9999 55345 10055 55397
rect 10107 55345 10127 55397
rect 9927 55289 10127 55345
rect 9927 55237 9947 55289
rect 9999 55237 10055 55289
rect 10107 55237 10127 55289
rect 9927 55181 10127 55237
rect 9927 55129 9947 55181
rect 9999 55129 10055 55181
rect 10107 55129 10127 55181
rect 9927 55073 10127 55129
rect 9927 55021 9947 55073
rect 9999 55021 10055 55073
rect 10107 55021 10127 55073
rect 9927 54965 10127 55021
rect 9927 54913 9947 54965
rect 9999 54913 10055 54965
rect 10107 54913 10127 54965
rect 9927 54857 10127 54913
rect 9927 54805 9947 54857
rect 9999 54805 10055 54857
rect 10107 54805 10127 54857
rect 9927 54749 10127 54805
rect 9927 54697 9947 54749
rect 9999 54697 10055 54749
rect 10107 54697 10127 54749
rect 9927 54641 10127 54697
rect 9927 54589 9947 54641
rect 9999 54589 10055 54641
rect 10107 54589 10127 54641
rect 9927 54533 10127 54589
rect 9927 54481 9947 54533
rect 9999 54481 10055 54533
rect 10107 54481 10127 54533
rect 9927 54425 10127 54481
rect 9927 54373 9947 54425
rect 9999 54373 10055 54425
rect 10107 54373 10127 54425
rect 9927 54317 10127 54373
rect 9927 54265 9947 54317
rect 9999 54265 10055 54317
rect 10107 54265 10127 54317
rect 9927 54209 10127 54265
rect 9927 54157 9947 54209
rect 9999 54157 10055 54209
rect 10107 54157 10127 54209
rect 9927 54101 10127 54157
rect 9927 54049 9947 54101
rect 9999 54049 10055 54101
rect 10107 54049 10127 54101
rect 9927 53993 10127 54049
rect 9927 53941 9947 53993
rect 9999 53941 10055 53993
rect 10107 53941 10127 53993
rect 9927 53885 10127 53941
rect 9927 53833 9947 53885
rect 9999 53833 10055 53885
rect 10107 53833 10127 53885
rect 9927 53777 10127 53833
rect 9927 53725 9947 53777
rect 9999 53725 10055 53777
rect 10107 53725 10127 53777
rect 9927 53669 10127 53725
rect 9927 53617 9947 53669
rect 9999 53617 10055 53669
rect 10107 53617 10127 53669
rect 9927 52572 10127 53617
rect 9927 52520 9947 52572
rect 9999 52520 10055 52572
rect 10107 52520 10127 52572
rect 9927 52464 10127 52520
rect 9927 52412 9947 52464
rect 9999 52412 10055 52464
rect 10107 52412 10127 52464
rect 9927 52356 10127 52412
rect 9927 52304 9947 52356
rect 9999 52304 10055 52356
rect 10107 52304 10127 52356
rect 9927 51619 10127 52304
rect 9927 51567 9947 51619
rect 9999 51567 10055 51619
rect 10107 51567 10127 51619
rect 9927 51511 10127 51567
rect 9927 51459 9947 51511
rect 9999 51459 10055 51511
rect 10107 51459 10127 51511
rect 9927 50948 10127 51459
rect 9927 50892 9937 50948
rect 9993 50892 10061 50948
rect 10117 50892 10127 50948
rect 9927 50824 10127 50892
rect 9927 50768 9937 50824
rect 9993 50768 10061 50824
rect 10117 50768 10127 50824
rect 9927 50700 10127 50768
rect 9927 50644 9937 50700
rect 9993 50685 10061 50700
rect 9927 50633 9947 50644
rect 9999 50633 10055 50685
rect 10117 50644 10127 50700
rect 10107 50633 10127 50644
rect 9927 50577 10127 50633
rect 9927 50576 9947 50577
rect 9927 50520 9937 50576
rect 9999 50525 10055 50577
rect 10107 50576 10127 50577
rect 9993 50520 10061 50525
rect 10117 50520 10127 50576
rect 9927 50452 10127 50520
rect 9927 50396 9937 50452
rect 9993 50396 10061 50452
rect 10117 50396 10127 50452
rect 9927 50328 10127 50396
rect 9927 50272 9937 50328
rect 9993 50272 10061 50328
rect 10117 50272 10127 50328
rect 9927 50204 10127 50272
rect 9927 50148 9937 50204
rect 9993 50148 10061 50204
rect 10117 50148 10127 50204
rect 9927 50080 10127 50148
rect 9927 50024 9937 50080
rect 9993 50024 10061 50080
rect 10117 50024 10127 50080
rect 9927 49956 10127 50024
rect 9927 49900 9937 49956
rect 9993 49900 10061 49956
rect 10117 49900 10127 49956
rect 9927 49832 10127 49900
rect 9927 49776 9937 49832
rect 9993 49776 10061 49832
rect 10117 49776 10127 49832
rect 9927 49751 10127 49776
rect 9927 49708 9947 49751
rect 9927 49652 9937 49708
rect 9999 49699 10055 49751
rect 10107 49708 10127 49751
rect 9993 49652 10061 49699
rect 10117 49652 10127 49708
rect 9927 49643 10127 49652
rect 9927 49591 9947 49643
rect 9999 49591 10055 49643
rect 10107 49591 10127 49643
rect 9927 48817 10127 49591
rect 9927 48765 9947 48817
rect 9999 48765 10055 48817
rect 10107 48765 10127 48817
rect 9927 48709 10127 48765
rect 9927 48657 9947 48709
rect 9999 48657 10055 48709
rect 10107 48657 10127 48709
rect 9927 47972 10127 48657
rect 9927 47920 9947 47972
rect 9999 47920 10055 47972
rect 10107 47920 10127 47972
rect 9927 47864 10127 47920
rect 9927 47812 9947 47864
rect 9999 47812 10055 47864
rect 10107 47812 10127 47864
rect 9927 47756 10127 47812
rect 9927 47704 9947 47756
rect 9999 47704 10055 47756
rect 10107 47704 10127 47756
rect 7265 46442 7713 47163
rect 9927 46442 10127 47704
rect 10187 57104 12237 57600
rect 10187 57052 10214 57104
rect 10266 57052 10322 57104
rect 10374 57052 10430 57104
rect 10482 57052 10538 57104
rect 10590 57052 10646 57104
rect 10698 57052 10754 57104
rect 10806 57052 10862 57104
rect 10914 57052 10970 57104
rect 11022 57052 11078 57104
rect 11130 57052 11186 57104
rect 11238 57052 11294 57104
rect 11346 57052 11402 57104
rect 11454 57052 11510 57104
rect 11562 57052 11618 57104
rect 11670 57052 11726 57104
rect 11778 57052 11834 57104
rect 11886 57052 11942 57104
rect 11994 57052 12050 57104
rect 12102 57052 12158 57104
rect 12210 57052 12237 57104
rect 10187 56643 12237 57052
rect 10187 56591 10775 56643
rect 10827 56591 10899 56643
rect 10951 56591 11023 56643
rect 11075 56591 12237 56643
rect 10187 56519 12237 56591
rect 10187 56467 10775 56519
rect 10827 56467 10899 56519
rect 10951 56467 11023 56519
rect 11075 56467 12237 56519
rect 10187 56395 12237 56467
rect 10187 56343 10775 56395
rect 10827 56343 10899 56395
rect 10951 56343 11023 56395
rect 11075 56343 12237 56395
rect 10187 56271 12237 56343
rect 10187 56219 10775 56271
rect 10827 56219 10899 56271
rect 10951 56219 11023 56271
rect 11075 56219 12237 56271
rect 10187 56147 12237 56219
rect 10187 56095 10775 56147
rect 10827 56095 10899 56147
rect 10951 56095 11023 56147
rect 11075 56095 12237 56147
rect 10187 56023 12237 56095
rect 10187 55971 10775 56023
rect 10827 55971 10899 56023
rect 10951 55971 11023 56023
rect 11075 55971 12237 56023
rect 10187 55899 12237 55971
rect 10187 55847 10775 55899
rect 10827 55847 10899 55899
rect 10951 55847 11023 55899
rect 11075 55847 12237 55899
rect 10187 55775 12237 55847
rect 10187 55723 10775 55775
rect 10827 55723 10899 55775
rect 10951 55723 11023 55775
rect 11075 55723 12237 55775
rect 10187 55651 12237 55723
rect 10187 55599 10775 55651
rect 10827 55599 10899 55651
rect 10951 55599 11023 55651
rect 11075 55599 12237 55651
rect 10187 55527 12237 55599
rect 10187 55475 10775 55527
rect 10827 55475 10899 55527
rect 10951 55475 11023 55527
rect 11075 55475 12237 55527
rect 10187 55403 12237 55475
rect 10187 55351 10775 55403
rect 10827 55351 10899 55403
rect 10951 55351 11023 55403
rect 11075 55351 12237 55403
rect 10187 55279 12237 55351
rect 10187 55227 10775 55279
rect 10827 55227 10899 55279
rect 10951 55227 11023 55279
rect 11075 55227 12237 55279
rect 10187 55155 12237 55227
rect 10187 55103 10775 55155
rect 10827 55103 10899 55155
rect 10951 55103 11023 55155
rect 11075 55103 12237 55155
rect 10187 55031 12237 55103
rect 10187 54979 10775 55031
rect 10827 54979 10899 55031
rect 10951 54979 11023 55031
rect 11075 54979 12237 55031
rect 10187 54907 12237 54979
rect 10187 54855 10775 54907
rect 10827 54855 10899 54907
rect 10951 54855 11023 54907
rect 11075 54855 12237 54907
rect 10187 54783 12237 54855
rect 10187 54731 10775 54783
rect 10827 54731 10899 54783
rect 10951 54731 11023 54783
rect 11075 54731 12237 54783
rect 10187 54659 12237 54731
rect 10187 54607 10775 54659
rect 10827 54607 10899 54659
rect 10951 54607 11023 54659
rect 11075 54607 12237 54659
rect 10187 54535 12237 54607
rect 10187 54483 10775 54535
rect 10827 54483 10899 54535
rect 10951 54483 11023 54535
rect 11075 54483 12237 54535
rect 10187 54411 12237 54483
rect 10187 54359 10775 54411
rect 10827 54359 10899 54411
rect 10951 54359 11023 54411
rect 11075 54359 12237 54411
rect 10187 54287 12237 54359
rect 10187 54235 10775 54287
rect 10827 54235 10899 54287
rect 10951 54235 11023 54287
rect 11075 54235 12237 54287
rect 10187 54163 12237 54235
rect 10187 54111 10775 54163
rect 10827 54111 10899 54163
rect 10951 54111 11023 54163
rect 11075 54111 12237 54163
rect 10187 54039 12237 54111
rect 10187 53987 10775 54039
rect 10827 53987 10899 54039
rect 10951 53987 11023 54039
rect 11075 53987 12237 54039
rect 10187 53915 12237 53987
rect 10187 53863 10775 53915
rect 10827 53863 10899 53915
rect 10951 53863 11023 53915
rect 11075 53863 12237 53915
rect 10187 53791 12237 53863
rect 10187 53739 10775 53791
rect 10827 53739 10899 53791
rect 10951 53739 11023 53791
rect 11075 53739 12237 53791
rect 10187 53667 12237 53739
rect 10187 53615 10775 53667
rect 10827 53615 10899 53667
rect 10951 53615 11023 53667
rect 11075 53615 12237 53667
rect 10187 53543 12237 53615
rect 10187 53491 10775 53543
rect 10827 53491 10899 53543
rect 10951 53491 11023 53543
rect 11075 53491 12237 53543
rect 10187 53483 12237 53491
rect 10187 53431 11191 53483
rect 11243 53431 11299 53483
rect 11351 53431 11407 53483
rect 11459 53431 11515 53483
rect 11567 53431 11623 53483
rect 11675 53431 11731 53483
rect 11783 53431 11839 53483
rect 11891 53431 11947 53483
rect 11999 53431 12055 53483
rect 12107 53431 12163 53483
rect 12215 53431 12237 53483
rect 10187 53419 12237 53431
rect 10187 53367 10775 53419
rect 10827 53367 10899 53419
rect 10951 53367 11023 53419
rect 11075 53375 12237 53419
rect 11075 53367 11191 53375
rect 10187 53323 11191 53367
rect 11243 53323 11299 53375
rect 11351 53323 11407 53375
rect 11459 53323 11515 53375
rect 11567 53323 11623 53375
rect 11675 53323 11731 53375
rect 11783 53323 11839 53375
rect 11891 53323 11947 53375
rect 11999 53323 12055 53375
rect 12107 53323 12163 53375
rect 12215 53323 12237 53375
rect 10187 53295 12237 53323
rect 10187 53243 10775 53295
rect 10827 53243 10899 53295
rect 10951 53243 11023 53295
rect 11075 53267 12237 53295
rect 11075 53243 11191 53267
rect 10187 53215 11191 53243
rect 11243 53215 11299 53267
rect 11351 53215 11407 53267
rect 11459 53215 11515 53267
rect 11567 53215 11623 53267
rect 11675 53215 11731 53267
rect 11783 53215 11839 53267
rect 11891 53215 11947 53267
rect 11999 53215 12055 53267
rect 12107 53215 12163 53267
rect 12215 53215 12237 53267
rect 10187 52548 12237 53215
rect 10187 52492 10254 52548
rect 10310 52492 10378 52548
rect 10434 52492 10502 52548
rect 10558 52492 10626 52548
rect 10682 52492 10750 52548
rect 10806 52492 10874 52548
rect 10930 52492 10998 52548
rect 11054 52492 11122 52548
rect 11178 52492 11246 52548
rect 11302 52492 11370 52548
rect 11426 52492 11494 52548
rect 11550 52492 11618 52548
rect 11674 52492 11742 52548
rect 11798 52492 11866 52548
rect 11922 52492 11990 52548
rect 12046 52492 12114 52548
rect 12170 52492 12237 52548
rect 10187 52424 12237 52492
rect 10187 52368 10254 52424
rect 10310 52368 10378 52424
rect 10434 52368 10502 52424
rect 10558 52368 10626 52424
rect 10682 52368 10750 52424
rect 10806 52368 10874 52424
rect 10930 52368 10998 52424
rect 11054 52368 11122 52424
rect 11178 52368 11246 52424
rect 11302 52368 11370 52424
rect 11426 52368 11494 52424
rect 11550 52368 11618 52424
rect 11674 52368 11742 52424
rect 11798 52368 11866 52424
rect 11922 52368 11990 52424
rect 12046 52368 12114 52424
rect 12170 52368 12237 52424
rect 10187 52300 12237 52368
rect 10187 52244 10254 52300
rect 10310 52244 10378 52300
rect 10434 52244 10502 52300
rect 10558 52244 10626 52300
rect 10682 52244 10750 52300
rect 10806 52244 10874 52300
rect 10930 52244 10998 52300
rect 11054 52244 11122 52300
rect 11178 52244 11246 52300
rect 11302 52244 11370 52300
rect 11426 52244 11494 52300
rect 11550 52244 11618 52300
rect 11674 52244 11742 52300
rect 11798 52244 11866 52300
rect 11922 52244 11990 52300
rect 12046 52244 12114 52300
rect 12170 52244 12237 52300
rect 10187 52176 12237 52244
rect 10187 52120 10254 52176
rect 10310 52120 10378 52176
rect 10434 52120 10502 52176
rect 10558 52120 10626 52176
rect 10682 52120 10750 52176
rect 10806 52120 10874 52176
rect 10930 52120 10998 52176
rect 11054 52120 11122 52176
rect 11178 52120 11246 52176
rect 11302 52120 11370 52176
rect 11426 52120 11494 52176
rect 11550 52120 11618 52176
rect 11674 52120 11742 52176
rect 11798 52120 11866 52176
rect 11922 52120 11990 52176
rect 12046 52120 12114 52176
rect 12170 52120 12237 52176
rect 10187 52052 12237 52120
rect 10187 52009 10254 52052
rect 10310 52009 10378 52052
rect 10434 52009 10502 52052
rect 10558 52009 10626 52052
rect 10682 52009 10750 52052
rect 10806 52009 10874 52052
rect 10930 52009 10998 52052
rect 11054 52009 11122 52052
rect 11178 52009 11246 52052
rect 11302 52009 11370 52052
rect 11426 52009 11494 52052
rect 11550 52009 11618 52052
rect 11674 52009 11742 52052
rect 11798 52009 11866 52052
rect 10187 51957 10253 52009
rect 10310 51996 10361 52009
rect 10434 51996 10469 52009
rect 10558 51996 10577 52009
rect 10682 51996 10685 52009
rect 10305 51957 10361 51996
rect 10413 51957 10469 51996
rect 10521 51957 10577 51996
rect 10629 51957 10685 51996
rect 10737 51996 10750 52009
rect 10845 51996 10874 52009
rect 10953 51996 10998 52009
rect 10737 51957 10793 51996
rect 10845 51957 10901 51996
rect 10953 51957 11009 51996
rect 11061 51957 11117 52009
rect 11178 51996 11225 52009
rect 11302 51996 11333 52009
rect 11426 51996 11441 52009
rect 11169 51957 11225 51996
rect 11277 51957 11333 51996
rect 11385 51957 11441 51996
rect 11493 51996 11494 52009
rect 11601 51996 11618 52009
rect 11709 51996 11742 52009
rect 11817 51996 11866 52009
rect 11922 51996 11990 52052
rect 12046 51996 12114 52052
rect 12170 51996 12237 52052
rect 11493 51957 11549 51996
rect 11601 51957 11657 51996
rect 11709 51957 11765 51996
rect 11817 51957 12237 51996
rect 10187 51928 12237 51957
rect 10187 51901 10254 51928
rect 10310 51901 10378 51928
rect 10434 51901 10502 51928
rect 10558 51901 10626 51928
rect 10682 51901 10750 51928
rect 10806 51901 10874 51928
rect 10930 51901 10998 51928
rect 11054 51901 11122 51928
rect 11178 51901 11246 51928
rect 11302 51901 11370 51928
rect 11426 51901 11494 51928
rect 11550 51901 11618 51928
rect 11674 51901 11742 51928
rect 11798 51901 11866 51928
rect 10187 51849 10253 51901
rect 10310 51872 10361 51901
rect 10434 51872 10469 51901
rect 10558 51872 10577 51901
rect 10682 51872 10685 51901
rect 10305 51849 10361 51872
rect 10413 51849 10469 51872
rect 10521 51849 10577 51872
rect 10629 51849 10685 51872
rect 10737 51872 10750 51901
rect 10845 51872 10874 51901
rect 10953 51872 10998 51901
rect 10737 51849 10793 51872
rect 10845 51849 10901 51872
rect 10953 51849 11009 51872
rect 11061 51849 11117 51901
rect 11178 51872 11225 51901
rect 11302 51872 11333 51901
rect 11426 51872 11441 51901
rect 11169 51849 11225 51872
rect 11277 51849 11333 51872
rect 11385 51849 11441 51872
rect 11493 51872 11494 51901
rect 11601 51872 11618 51901
rect 11709 51872 11742 51901
rect 11817 51872 11866 51901
rect 11922 51872 11990 51928
rect 12046 51872 12114 51928
rect 12170 51872 12237 51928
rect 11493 51849 11549 51872
rect 11601 51849 11657 51872
rect 11709 51849 11765 51872
rect 11817 51849 12237 51872
rect 10187 51804 12237 51849
rect 10187 51748 10254 51804
rect 10310 51748 10378 51804
rect 10434 51748 10502 51804
rect 10558 51748 10626 51804
rect 10682 51748 10750 51804
rect 10806 51748 10874 51804
rect 10930 51748 10998 51804
rect 11054 51748 11122 51804
rect 11178 51748 11246 51804
rect 11302 51748 11370 51804
rect 11426 51748 11494 51804
rect 11550 51748 11618 51804
rect 11674 51748 11742 51804
rect 11798 51748 11866 51804
rect 11922 51748 11990 51804
rect 12046 51748 12114 51804
rect 12170 51748 12237 51804
rect 10187 51680 12237 51748
rect 10187 51624 10254 51680
rect 10310 51624 10378 51680
rect 10434 51624 10502 51680
rect 10558 51624 10626 51680
rect 10682 51624 10750 51680
rect 10806 51624 10874 51680
rect 10930 51624 10998 51680
rect 11054 51624 11122 51680
rect 11178 51624 11246 51680
rect 11302 51624 11370 51680
rect 11426 51624 11494 51680
rect 11550 51624 11618 51680
rect 11674 51624 11742 51680
rect 11798 51624 11866 51680
rect 11922 51624 11990 51680
rect 12046 51624 12114 51680
rect 12170 51624 12237 51680
rect 10187 51556 12237 51624
rect 10187 51500 10254 51556
rect 10310 51500 10378 51556
rect 10434 51500 10502 51556
rect 10558 51500 10626 51556
rect 10682 51500 10750 51556
rect 10806 51500 10874 51556
rect 10930 51500 10998 51556
rect 11054 51500 11122 51556
rect 11178 51500 11246 51556
rect 11302 51500 11370 51556
rect 11426 51500 11494 51556
rect 11550 51500 11618 51556
rect 11674 51500 11742 51556
rect 11798 51500 11866 51556
rect 11922 51500 11990 51556
rect 12046 51500 12114 51556
rect 12170 51500 12237 51556
rect 10187 51432 12237 51500
rect 10187 51376 10254 51432
rect 10310 51376 10378 51432
rect 10434 51376 10502 51432
rect 10558 51376 10626 51432
rect 10682 51376 10750 51432
rect 10806 51376 10874 51432
rect 10930 51376 10998 51432
rect 11054 51376 11122 51432
rect 11178 51376 11246 51432
rect 11302 51376 11370 51432
rect 11426 51376 11494 51432
rect 11550 51376 11618 51432
rect 11674 51376 11742 51432
rect 11798 51376 11866 51432
rect 11922 51376 11990 51432
rect 12046 51376 12114 51432
rect 12170 51376 12237 51432
rect 10187 51308 12237 51376
rect 10187 51252 10254 51308
rect 10310 51252 10378 51308
rect 10434 51252 10502 51308
rect 10558 51252 10626 51308
rect 10682 51252 10750 51308
rect 10806 51252 10874 51308
rect 10930 51252 10998 51308
rect 11054 51252 11122 51308
rect 11178 51252 11246 51308
rect 11302 51252 11370 51308
rect 11426 51252 11494 51308
rect 11550 51252 11618 51308
rect 11674 51252 11742 51308
rect 11798 51252 11866 51308
rect 11922 51252 11990 51308
rect 12046 51252 12114 51308
rect 12170 51252 12237 51308
rect 10187 51206 12237 51252
rect 10187 51154 10253 51206
rect 10305 51154 10361 51206
rect 10413 51154 10469 51206
rect 10521 51154 10577 51206
rect 10629 51154 10685 51206
rect 10737 51154 10793 51206
rect 10845 51154 10901 51206
rect 10953 51154 11009 51206
rect 11061 51154 11117 51206
rect 11169 51154 11225 51206
rect 11277 51154 11333 51206
rect 11385 51154 11441 51206
rect 11493 51154 11549 51206
rect 11601 51154 11657 51206
rect 11709 51154 11765 51206
rect 11817 51154 12237 51206
rect 10187 51098 12237 51154
rect 10187 51046 10253 51098
rect 10305 51046 10361 51098
rect 10413 51046 10469 51098
rect 10521 51046 10577 51098
rect 10629 51046 10685 51098
rect 10737 51046 10793 51098
rect 10845 51046 10901 51098
rect 10953 51046 11009 51098
rect 11061 51046 11117 51098
rect 11169 51046 11225 51098
rect 11277 51046 11333 51098
rect 11385 51046 11441 51098
rect 11493 51046 11549 51098
rect 11601 51046 11657 51098
rect 11709 51046 11765 51098
rect 11817 51046 12237 51098
rect 10187 50990 12237 51046
rect 10187 50938 10253 50990
rect 10305 50938 10361 50990
rect 10413 50938 10469 50990
rect 10521 50938 10577 50990
rect 10629 50938 10685 50990
rect 10737 50938 10793 50990
rect 10845 50938 10901 50990
rect 10953 50938 11009 50990
rect 11061 50938 11117 50990
rect 11169 50938 11225 50990
rect 11277 50938 11333 50990
rect 11385 50938 11441 50990
rect 11493 50938 11549 50990
rect 11601 50938 11657 50990
rect 11709 50938 11765 50990
rect 11817 50938 12237 50990
rect 10187 50272 12237 50938
rect 10187 50220 10253 50272
rect 10305 50220 10361 50272
rect 10413 50220 10469 50272
rect 10521 50220 10577 50272
rect 10629 50220 10685 50272
rect 10737 50220 10793 50272
rect 10845 50220 10901 50272
rect 10953 50220 11009 50272
rect 11061 50220 11117 50272
rect 11169 50220 11225 50272
rect 11277 50220 11333 50272
rect 11385 50220 11441 50272
rect 11493 50220 11549 50272
rect 11601 50220 11657 50272
rect 11709 50220 11765 50272
rect 11817 50220 12237 50272
rect 10187 50164 12237 50220
rect 10187 50112 10253 50164
rect 10305 50112 10361 50164
rect 10413 50112 10469 50164
rect 10521 50112 10577 50164
rect 10629 50112 10685 50164
rect 10737 50112 10793 50164
rect 10845 50112 10901 50164
rect 10953 50112 11009 50164
rect 11061 50112 11117 50164
rect 11169 50112 11225 50164
rect 11277 50112 11333 50164
rect 11385 50112 11441 50164
rect 11493 50112 11549 50164
rect 11601 50112 11657 50164
rect 11709 50112 11765 50164
rect 11817 50112 12237 50164
rect 10187 50056 12237 50112
rect 10187 50004 10253 50056
rect 10305 50004 10361 50056
rect 10413 50004 10469 50056
rect 10521 50004 10577 50056
rect 10629 50004 10685 50056
rect 10737 50004 10793 50056
rect 10845 50004 10901 50056
rect 10953 50004 11009 50056
rect 11061 50004 11117 50056
rect 11169 50004 11225 50056
rect 11277 50004 11333 50056
rect 11385 50004 11441 50056
rect 11493 50004 11549 50056
rect 11601 50004 11657 50056
rect 11709 50004 11765 50056
rect 11817 50004 12237 50056
rect 10187 49338 12237 50004
rect 10187 49286 10253 49338
rect 10305 49286 10361 49338
rect 10413 49286 10469 49338
rect 10521 49286 10577 49338
rect 10629 49286 10685 49338
rect 10737 49286 10793 49338
rect 10845 49286 10901 49338
rect 10953 49286 11009 49338
rect 11061 49286 11117 49338
rect 11169 49286 11225 49338
rect 11277 49286 11333 49338
rect 11385 49286 11441 49338
rect 11493 49286 11549 49338
rect 11601 49286 11657 49338
rect 11709 49286 11765 49338
rect 11817 49286 12237 49338
rect 10187 49230 12237 49286
rect 10187 49178 10253 49230
rect 10305 49178 10361 49230
rect 10413 49178 10469 49230
rect 10521 49178 10577 49230
rect 10629 49178 10685 49230
rect 10737 49178 10793 49230
rect 10845 49178 10901 49230
rect 10953 49178 11009 49230
rect 11061 49178 11117 49230
rect 11169 49178 11225 49230
rect 11277 49178 11333 49230
rect 11385 49178 11441 49230
rect 11493 49178 11549 49230
rect 11601 49178 11657 49230
rect 11709 49178 11765 49230
rect 11817 49178 12237 49230
rect 10187 49122 12237 49178
rect 10187 49070 10253 49122
rect 10305 49070 10361 49122
rect 10413 49070 10469 49122
rect 10521 49070 10577 49122
rect 10629 49070 10685 49122
rect 10737 49070 10793 49122
rect 10845 49070 10901 49122
rect 10953 49070 11009 49122
rect 11061 49070 11117 49122
rect 11169 49070 11225 49122
rect 11277 49070 11333 49122
rect 11385 49070 11441 49122
rect 11493 49070 11549 49122
rect 11601 49070 11657 49122
rect 11709 49070 11765 49122
rect 11817 49070 12237 49122
rect 10187 48427 12237 49070
rect 10187 48375 10253 48427
rect 10305 48375 10361 48427
rect 10413 48375 10469 48427
rect 10521 48375 10577 48427
rect 10629 48375 10685 48427
rect 10737 48375 10793 48427
rect 10845 48375 10901 48427
rect 10953 48375 11009 48427
rect 11061 48375 11117 48427
rect 11169 48375 11225 48427
rect 11277 48375 11333 48427
rect 11385 48375 11441 48427
rect 11493 48375 11549 48427
rect 11601 48375 11657 48427
rect 11709 48375 11765 48427
rect 11817 48375 12237 48427
rect 10187 48319 12237 48375
rect 10187 48267 10253 48319
rect 10305 48267 10361 48319
rect 10413 48267 10469 48319
rect 10521 48267 10577 48319
rect 10629 48267 10685 48319
rect 10737 48267 10793 48319
rect 10845 48267 10901 48319
rect 10953 48267 11009 48319
rect 11061 48267 11117 48319
rect 11169 48267 11225 48319
rect 11277 48267 11333 48319
rect 11385 48267 11441 48319
rect 11493 48267 11549 48319
rect 11601 48267 11657 48319
rect 11709 48267 11765 48319
rect 11817 48267 12237 48319
rect 10187 47163 12237 48267
rect 12297 56741 12497 57278
rect 12297 56689 12317 56741
rect 12369 56689 12425 56741
rect 12477 56689 12497 56741
rect 12297 53621 12497 56689
rect 12297 53569 12317 53621
rect 12369 53569 12425 53621
rect 12477 53569 12497 53621
rect 12297 52594 12497 53569
rect 12297 52542 12336 52594
rect 12388 52542 12497 52594
rect 12297 52486 12497 52542
rect 12297 52434 12336 52486
rect 12388 52434 12497 52486
rect 12297 52378 12497 52434
rect 12297 52326 12336 52378
rect 12388 52326 12497 52378
rect 12297 52270 12497 52326
rect 12297 52218 12336 52270
rect 12388 52218 12497 52270
rect 12297 52162 12497 52218
rect 12297 52110 12336 52162
rect 12388 52110 12497 52162
rect 12297 52054 12497 52110
rect 12297 52002 12336 52054
rect 12388 52002 12497 52054
rect 12297 51946 12497 52002
rect 12297 51894 12336 51946
rect 12388 51894 12497 51946
rect 12297 51838 12497 51894
rect 12297 51786 12336 51838
rect 12388 51786 12497 51838
rect 12297 51730 12497 51786
rect 12297 51678 12336 51730
rect 12388 51678 12497 51730
rect 12297 51622 12497 51678
rect 12297 51570 12336 51622
rect 12388 51570 12497 51622
rect 12297 51514 12497 51570
rect 12297 51462 12336 51514
rect 12388 51462 12497 51514
rect 12297 51406 12497 51462
rect 12297 51354 12336 51406
rect 12388 51354 12497 51406
rect 12297 51298 12497 51354
rect 12297 51246 12336 51298
rect 12388 51246 12497 51298
rect 12297 51190 12497 51246
rect 12297 51138 12336 51190
rect 12388 51138 12497 51190
rect 12297 51082 12497 51138
rect 12297 51030 12336 51082
rect 12388 51030 12497 51082
rect 12297 50974 12497 51030
rect 12297 50948 12336 50974
rect 12388 50948 12497 50974
rect 12297 50892 12307 50948
rect 12388 50922 12431 50948
rect 12363 50892 12431 50922
rect 12487 50892 12497 50948
rect 12297 50866 12497 50892
rect 12297 50824 12336 50866
rect 12388 50824 12497 50866
rect 12297 50768 12307 50824
rect 12388 50814 12431 50824
rect 12363 50768 12431 50814
rect 12487 50768 12497 50824
rect 12297 50758 12497 50768
rect 12297 50706 12336 50758
rect 12388 50706 12497 50758
rect 12297 50700 12497 50706
rect 12297 50644 12307 50700
rect 12363 50650 12431 50700
rect 12388 50644 12431 50650
rect 12487 50644 12497 50700
rect 12297 50598 12336 50644
rect 12388 50598 12497 50644
rect 12297 50576 12497 50598
rect 12297 50520 12307 50576
rect 12363 50542 12431 50576
rect 12388 50520 12431 50542
rect 12487 50520 12497 50576
rect 12297 50490 12336 50520
rect 12388 50490 12497 50520
rect 12297 50452 12497 50490
rect 12297 50396 12307 50452
rect 12363 50434 12431 50452
rect 12388 50396 12431 50434
rect 12487 50396 12497 50452
rect 12297 50382 12336 50396
rect 12388 50382 12497 50396
rect 12297 50328 12497 50382
rect 12297 50272 12307 50328
rect 12363 50326 12431 50328
rect 12388 50274 12431 50326
rect 12363 50272 12431 50274
rect 12487 50272 12497 50328
rect 12297 50218 12497 50272
rect 12297 50204 12336 50218
rect 12388 50204 12497 50218
rect 12297 50148 12307 50204
rect 12388 50166 12431 50204
rect 12363 50148 12431 50166
rect 12487 50148 12497 50204
rect 12297 50110 12497 50148
rect 12297 50080 12336 50110
rect 12388 50080 12497 50110
rect 12297 50024 12307 50080
rect 12388 50058 12431 50080
rect 12363 50024 12431 50058
rect 12487 50024 12497 50080
rect 12297 50002 12497 50024
rect 12297 49956 12336 50002
rect 12388 49956 12497 50002
rect 12297 49900 12307 49956
rect 12388 49950 12431 49956
rect 12363 49900 12431 49950
rect 12487 49900 12497 49956
rect 12297 49894 12497 49900
rect 12297 49842 12336 49894
rect 12388 49842 12497 49894
rect 12297 49832 12497 49842
rect 12297 49776 12307 49832
rect 12363 49786 12431 49832
rect 12388 49776 12431 49786
rect 12487 49776 12497 49832
rect 12297 49734 12336 49776
rect 12388 49734 12497 49776
rect 12297 49708 12497 49734
rect 12297 49652 12307 49708
rect 12363 49678 12431 49708
rect 12388 49652 12431 49678
rect 12487 49652 12497 49708
rect 12297 49626 12336 49652
rect 12388 49626 12497 49652
rect 12297 49570 12497 49626
rect 12297 49518 12336 49570
rect 12388 49518 12497 49570
rect 12297 49462 12497 49518
rect 12297 49410 12336 49462
rect 12388 49410 12497 49462
rect 12297 49354 12497 49410
rect 12297 49302 12336 49354
rect 12388 49302 12497 49354
rect 12297 49246 12497 49302
rect 12297 49194 12336 49246
rect 12388 49194 12497 49246
rect 12297 49138 12497 49194
rect 12297 49086 12336 49138
rect 12388 49086 12497 49138
rect 12297 49030 12497 49086
rect 12297 48978 12336 49030
rect 12388 48978 12497 49030
rect 12297 48922 12497 48978
rect 12297 48870 12336 48922
rect 12388 48870 12497 48922
rect 12297 48814 12497 48870
rect 12297 48762 12336 48814
rect 12388 48762 12497 48814
rect 12297 48706 12497 48762
rect 12297 48654 12336 48706
rect 12388 48654 12497 48706
rect 12297 48598 12497 48654
rect 12297 48546 12336 48598
rect 12388 48546 12497 48598
rect 12297 48490 12497 48546
rect 12297 48438 12336 48490
rect 12388 48438 12497 48490
rect 12297 48382 12497 48438
rect 12297 48330 12336 48382
rect 12388 48330 12497 48382
rect 12297 48274 12497 48330
rect 12297 48222 12336 48274
rect 12388 48222 12497 48274
rect 12297 48166 12497 48222
rect 12297 48114 12336 48166
rect 12388 48114 12497 48166
rect 12297 48058 12497 48114
rect 12297 48006 12336 48058
rect 12388 48006 12497 48058
rect 12297 47950 12497 48006
rect 12297 47898 12336 47950
rect 12388 47898 12497 47950
rect 12297 47842 12497 47898
rect 12297 47790 12336 47842
rect 12388 47790 12497 47842
rect 12297 47734 12497 47790
rect 12297 47682 12336 47734
rect 12388 47682 12497 47734
rect 12297 46442 12497 47682
rect 12817 57104 14717 57600
rect 12817 57052 12931 57104
rect 12983 57052 13039 57104
rect 13091 57052 13147 57104
rect 13199 57052 13255 57104
rect 13307 57052 13363 57104
rect 13415 57052 13471 57104
rect 13523 57052 13579 57104
rect 13631 57052 13687 57104
rect 13739 57052 13795 57104
rect 13847 57052 13903 57104
rect 13955 57052 14011 57104
rect 14063 57052 14119 57104
rect 14171 57052 14227 57104
rect 14279 57052 14335 57104
rect 14387 57052 14443 57104
rect 14495 57052 14551 57104
rect 14603 57052 14717 57104
rect 12817 56643 14717 57052
rect 12817 56591 14185 56643
rect 14237 56591 14309 56643
rect 14361 56591 14433 56643
rect 14485 56591 14557 56643
rect 14609 56591 14717 56643
rect 12817 56519 14717 56591
rect 12817 56467 14185 56519
rect 14237 56467 14309 56519
rect 14361 56467 14433 56519
rect 14485 56467 14557 56519
rect 14609 56467 14717 56519
rect 12817 56395 14717 56467
rect 12817 56343 14185 56395
rect 14237 56343 14309 56395
rect 14361 56343 14433 56395
rect 14485 56343 14557 56395
rect 14609 56343 14717 56395
rect 12817 56271 14717 56343
rect 12817 56219 14185 56271
rect 14237 56219 14309 56271
rect 14361 56219 14433 56271
rect 14485 56219 14557 56271
rect 14609 56219 14717 56271
rect 12817 56147 14717 56219
rect 12817 56095 14185 56147
rect 14237 56095 14309 56147
rect 14361 56095 14433 56147
rect 14485 56095 14557 56147
rect 14609 56095 14717 56147
rect 12817 56023 14717 56095
rect 12817 55971 14185 56023
rect 14237 55971 14309 56023
rect 14361 55971 14433 56023
rect 14485 55971 14557 56023
rect 14609 55971 14717 56023
rect 12817 55899 14717 55971
rect 12817 55847 14185 55899
rect 14237 55847 14309 55899
rect 14361 55847 14433 55899
rect 14485 55847 14557 55899
rect 14609 55847 14717 55899
rect 12817 55775 14717 55847
rect 12817 55723 14185 55775
rect 14237 55723 14309 55775
rect 14361 55723 14433 55775
rect 14485 55723 14557 55775
rect 14609 55723 14717 55775
rect 12817 55651 14717 55723
rect 12817 55599 14185 55651
rect 14237 55599 14309 55651
rect 14361 55599 14433 55651
rect 14485 55599 14557 55651
rect 14609 55599 14717 55651
rect 12817 55527 14717 55599
rect 12817 55475 14185 55527
rect 14237 55475 14309 55527
rect 14361 55475 14433 55527
rect 14485 55475 14557 55527
rect 14609 55475 14717 55527
rect 12817 55403 14717 55475
rect 12817 55351 14185 55403
rect 14237 55351 14309 55403
rect 14361 55351 14433 55403
rect 14485 55351 14557 55403
rect 14609 55351 14717 55403
rect 12817 55279 14717 55351
rect 12817 55227 14185 55279
rect 14237 55227 14309 55279
rect 14361 55227 14433 55279
rect 14485 55227 14557 55279
rect 14609 55227 14717 55279
rect 12817 55155 14717 55227
rect 12817 55103 14185 55155
rect 14237 55103 14309 55155
rect 14361 55103 14433 55155
rect 14485 55103 14557 55155
rect 14609 55103 14717 55155
rect 12817 55031 14717 55103
rect 12817 54979 14185 55031
rect 14237 54979 14309 55031
rect 14361 54979 14433 55031
rect 14485 54979 14557 55031
rect 14609 54979 14717 55031
rect 12817 54907 14717 54979
rect 12817 54855 14185 54907
rect 14237 54855 14309 54907
rect 14361 54855 14433 54907
rect 14485 54855 14557 54907
rect 14609 54855 14717 54907
rect 12817 54783 14717 54855
rect 12817 54731 14185 54783
rect 14237 54731 14309 54783
rect 14361 54731 14433 54783
rect 14485 54731 14557 54783
rect 14609 54731 14717 54783
rect 12817 54659 14717 54731
rect 12817 54607 14185 54659
rect 14237 54607 14309 54659
rect 14361 54607 14433 54659
rect 14485 54607 14557 54659
rect 14609 54607 14717 54659
rect 12817 54535 14717 54607
rect 12817 54483 14185 54535
rect 14237 54483 14309 54535
rect 14361 54483 14433 54535
rect 14485 54483 14557 54535
rect 14609 54483 14717 54535
rect 12817 54411 14717 54483
rect 12817 54359 14185 54411
rect 14237 54359 14309 54411
rect 14361 54359 14433 54411
rect 14485 54359 14557 54411
rect 14609 54359 14717 54411
rect 12817 54287 14717 54359
rect 12817 54235 14185 54287
rect 14237 54235 14309 54287
rect 14361 54235 14433 54287
rect 14485 54235 14557 54287
rect 14609 54235 14717 54287
rect 12817 54163 14717 54235
rect 12817 54111 14185 54163
rect 14237 54111 14309 54163
rect 14361 54111 14433 54163
rect 14485 54111 14557 54163
rect 14609 54111 14717 54163
rect 12817 54039 14717 54111
rect 12817 53987 14185 54039
rect 14237 53987 14309 54039
rect 14361 53987 14433 54039
rect 14485 53987 14557 54039
rect 14609 53987 14717 54039
rect 12817 53915 14717 53987
rect 12817 53863 14185 53915
rect 14237 53863 14309 53915
rect 14361 53863 14433 53915
rect 14485 53863 14557 53915
rect 14609 53863 14717 53915
rect 12817 53791 14717 53863
rect 12817 53739 14185 53791
rect 14237 53739 14309 53791
rect 14361 53739 14433 53791
rect 14485 53739 14557 53791
rect 14609 53739 14717 53791
rect 12817 53667 14717 53739
rect 12817 53615 14185 53667
rect 14237 53615 14309 53667
rect 14361 53615 14433 53667
rect 14485 53615 14557 53667
rect 14609 53615 14717 53667
rect 12817 53543 14717 53615
rect 12817 53491 14185 53543
rect 14237 53491 14309 53543
rect 14361 53491 14433 53543
rect 14485 53491 14557 53543
rect 14609 53491 14717 53543
rect 12817 53483 14717 53491
rect 12817 53431 12869 53483
rect 12921 53431 12977 53483
rect 13029 53431 13085 53483
rect 13137 53431 13193 53483
rect 13245 53431 13301 53483
rect 13353 53431 13409 53483
rect 13461 53431 13517 53483
rect 13569 53431 13625 53483
rect 13677 53431 13733 53483
rect 13785 53431 13841 53483
rect 13893 53431 13949 53483
rect 14001 53431 14057 53483
rect 14109 53431 14717 53483
rect 12817 53419 14717 53431
rect 12817 53375 14185 53419
rect 12817 53323 12869 53375
rect 12921 53323 12977 53375
rect 13029 53323 13085 53375
rect 13137 53323 13193 53375
rect 13245 53323 13301 53375
rect 13353 53323 13409 53375
rect 13461 53323 13517 53375
rect 13569 53323 13625 53375
rect 13677 53323 13733 53375
rect 13785 53323 13841 53375
rect 13893 53323 13949 53375
rect 14001 53323 14057 53375
rect 14109 53367 14185 53375
rect 14237 53367 14309 53419
rect 14361 53367 14433 53419
rect 14485 53367 14557 53419
rect 14609 53367 14717 53419
rect 14109 53323 14717 53367
rect 12817 53295 14717 53323
rect 12817 53267 14185 53295
rect 12817 53215 12869 53267
rect 12921 53215 12977 53267
rect 13029 53215 13085 53267
rect 13137 53215 13193 53267
rect 13245 53215 13301 53267
rect 13353 53215 13409 53267
rect 13461 53215 13517 53267
rect 13569 53215 13625 53267
rect 13677 53215 13733 53267
rect 13785 53215 13841 53267
rect 13893 53215 13949 53267
rect 14001 53215 14057 53267
rect 14109 53243 14185 53267
rect 14237 53243 14309 53295
rect 14361 53243 14433 53295
rect 14485 53243 14557 53295
rect 14609 53243 14717 53295
rect 14109 53215 14717 53243
rect 12817 52548 14717 53215
rect 12817 52492 12871 52548
rect 12927 52492 12995 52548
rect 13051 52492 13119 52548
rect 13175 52492 13243 52548
rect 13299 52492 13367 52548
rect 13423 52492 13491 52548
rect 13547 52492 13615 52548
rect 13671 52492 13739 52548
rect 13795 52492 13863 52548
rect 13919 52492 13987 52548
rect 14043 52492 14111 52548
rect 14167 52492 14235 52548
rect 14291 52492 14359 52548
rect 14415 52492 14483 52548
rect 14539 52492 14607 52548
rect 14663 52492 14717 52548
rect 12817 52424 14717 52492
rect 12817 52368 12871 52424
rect 12927 52368 12995 52424
rect 13051 52368 13119 52424
rect 13175 52368 13243 52424
rect 13299 52368 13367 52424
rect 13423 52368 13491 52424
rect 13547 52368 13615 52424
rect 13671 52368 13739 52424
rect 13795 52368 13863 52424
rect 13919 52368 13987 52424
rect 14043 52368 14111 52424
rect 14167 52368 14235 52424
rect 14291 52368 14359 52424
rect 14415 52368 14483 52424
rect 14539 52368 14607 52424
rect 14663 52368 14717 52424
rect 12817 52300 14717 52368
rect 12817 52244 12871 52300
rect 12927 52244 12995 52300
rect 13051 52244 13119 52300
rect 13175 52244 13243 52300
rect 13299 52244 13367 52300
rect 13423 52244 13491 52300
rect 13547 52244 13615 52300
rect 13671 52244 13739 52300
rect 13795 52244 13863 52300
rect 13919 52244 13987 52300
rect 14043 52244 14111 52300
rect 14167 52244 14235 52300
rect 14291 52244 14359 52300
rect 14415 52244 14483 52300
rect 14539 52244 14607 52300
rect 14663 52244 14717 52300
rect 12817 52176 14717 52244
rect 12817 52120 12871 52176
rect 12927 52120 12995 52176
rect 13051 52120 13119 52176
rect 13175 52120 13243 52176
rect 13299 52120 13367 52176
rect 13423 52120 13491 52176
rect 13547 52120 13615 52176
rect 13671 52120 13739 52176
rect 13795 52120 13863 52176
rect 13919 52120 13987 52176
rect 14043 52120 14111 52176
rect 14167 52120 14235 52176
rect 14291 52120 14359 52176
rect 14415 52120 14483 52176
rect 14539 52120 14607 52176
rect 14663 52120 14717 52176
rect 12817 52052 14717 52120
rect 12817 51996 12871 52052
rect 12927 51996 12995 52052
rect 13051 51996 13119 52052
rect 13175 51996 13243 52052
rect 13299 51996 13367 52052
rect 13423 51996 13491 52052
rect 13547 51996 13615 52052
rect 13671 51996 13739 52052
rect 13795 51996 13863 52052
rect 13919 51996 13987 52052
rect 14043 51996 14111 52052
rect 14167 51996 14235 52052
rect 14291 51996 14359 52052
rect 14415 51996 14483 52052
rect 14539 51996 14607 52052
rect 14663 51996 14717 52052
rect 12817 51928 14717 51996
rect 12817 51872 12871 51928
rect 12927 51872 12995 51928
rect 13051 51872 13119 51928
rect 13175 51872 13243 51928
rect 13299 51872 13367 51928
rect 13423 51872 13491 51928
rect 13547 51872 13615 51928
rect 13671 51872 13739 51928
rect 13795 51872 13863 51928
rect 13919 51872 13987 51928
rect 14043 51872 14111 51928
rect 14167 51872 14235 51928
rect 14291 51872 14359 51928
rect 14415 51872 14483 51928
rect 14539 51872 14607 51928
rect 14663 51872 14717 51928
rect 12817 51804 14717 51872
rect 12817 51748 12871 51804
rect 12927 51748 12995 51804
rect 13051 51748 13119 51804
rect 13175 51748 13243 51804
rect 13299 51748 13367 51804
rect 13423 51748 13491 51804
rect 13547 51748 13615 51804
rect 13671 51748 13739 51804
rect 13795 51748 13863 51804
rect 13919 51748 13987 51804
rect 14043 51748 14111 51804
rect 14167 51748 14235 51804
rect 14291 51748 14359 51804
rect 14415 51748 14483 51804
rect 14539 51748 14607 51804
rect 14663 51748 14717 51804
rect 12817 51680 14717 51748
rect 12817 51624 12871 51680
rect 12927 51624 12995 51680
rect 13051 51624 13119 51680
rect 13175 51624 13243 51680
rect 13299 51624 13367 51680
rect 13423 51624 13491 51680
rect 13547 51624 13615 51680
rect 13671 51624 13739 51680
rect 13795 51624 13863 51680
rect 13919 51624 13987 51680
rect 14043 51624 14111 51680
rect 14167 51624 14235 51680
rect 14291 51624 14359 51680
rect 14415 51624 14483 51680
rect 14539 51624 14607 51680
rect 14663 51624 14717 51680
rect 12817 51556 14717 51624
rect 12817 51500 12871 51556
rect 12927 51500 12995 51556
rect 13051 51500 13119 51556
rect 13175 51500 13243 51556
rect 13299 51500 13367 51556
rect 13423 51500 13491 51556
rect 13547 51500 13615 51556
rect 13671 51500 13739 51556
rect 13795 51500 13863 51556
rect 13919 51500 13987 51556
rect 14043 51500 14111 51556
rect 14167 51500 14235 51556
rect 14291 51500 14359 51556
rect 14415 51500 14483 51556
rect 14539 51500 14607 51556
rect 14663 51500 14717 51556
rect 12817 51432 14717 51500
rect 12817 51376 12871 51432
rect 12927 51376 12995 51432
rect 13051 51376 13119 51432
rect 13175 51376 13243 51432
rect 13299 51376 13367 51432
rect 13423 51376 13491 51432
rect 13547 51376 13615 51432
rect 13671 51376 13739 51432
rect 13795 51376 13863 51432
rect 13919 51376 13987 51432
rect 14043 51376 14111 51432
rect 14167 51376 14235 51432
rect 14291 51376 14359 51432
rect 14415 51376 14483 51432
rect 14539 51376 14607 51432
rect 14663 51376 14717 51432
rect 12817 51308 14717 51376
rect 12817 51252 12871 51308
rect 12927 51252 12995 51308
rect 13051 51252 13119 51308
rect 13175 51252 13243 51308
rect 13299 51252 13367 51308
rect 13423 51252 13491 51308
rect 13547 51252 13615 51308
rect 13671 51252 13739 51308
rect 13795 51252 13863 51308
rect 13919 51252 13987 51308
rect 14043 51252 14111 51308
rect 14167 51252 14235 51308
rect 14291 51252 14359 51308
rect 14415 51252 14483 51308
rect 14539 51252 14607 51308
rect 14663 51252 14717 51308
rect 12817 47163 14717 51252
rect 14892 57259 14989 57271
rect 14892 57207 14904 57259
rect 14956 57207 14989 57259
rect 14892 57151 14989 57207
rect 14892 57099 14904 57151
rect 14956 57099 14989 57151
rect 14892 57043 14989 57099
rect 14892 56991 14904 57043
rect 14956 56991 14989 57043
rect 14892 56935 14989 56991
rect 14892 56883 14904 56935
rect 14956 56883 14989 56935
rect 14892 56827 14989 56883
rect 14892 56775 14904 56827
rect 14956 56775 14989 56827
rect 14892 56719 14989 56775
rect 14892 56667 14904 56719
rect 14956 56667 14989 56719
rect 14892 56611 14989 56667
rect 14892 56559 14904 56611
rect 14956 56559 14989 56611
rect 14892 56503 14989 56559
rect 14892 56451 14904 56503
rect 14956 56451 14989 56503
rect 14892 56395 14989 56451
rect 14892 56343 14904 56395
rect 14956 56343 14989 56395
rect 14892 56287 14989 56343
rect 14892 56235 14904 56287
rect 14956 56235 14989 56287
rect 14892 56179 14989 56235
rect 14892 56127 14904 56179
rect 14956 56127 14989 56179
rect 14892 56071 14989 56127
rect 14892 56019 14904 56071
rect 14956 56019 14989 56071
rect 14892 54174 14989 56019
rect 14892 54122 14904 54174
rect 14956 54122 14989 54174
rect 14892 54066 14989 54122
rect 14892 54014 14904 54066
rect 14956 54014 14989 54066
rect 14892 53958 14989 54014
rect 14892 53906 14904 53958
rect 14956 53906 14989 53958
rect 14892 53850 14989 53906
rect 14892 53798 14904 53850
rect 14956 53798 14989 53850
rect 14892 53742 14989 53798
rect 14892 53690 14904 53742
rect 14956 53690 14989 53742
rect 14892 53634 14989 53690
rect 14892 53582 14904 53634
rect 14956 53582 14989 53634
rect 14892 53526 14989 53582
rect 14892 53474 14904 53526
rect 14956 53474 14989 53526
rect 14892 53418 14989 53474
rect 14892 53366 14904 53418
rect 14956 53366 14989 53418
rect 14892 53310 14989 53366
rect 14892 53258 14904 53310
rect 14956 53258 14989 53310
rect 14892 53202 14989 53258
rect 14892 53150 14904 53202
rect 14956 53150 14989 53202
rect 14892 53094 14989 53150
rect 14892 53042 14904 53094
rect 14956 53042 14989 53094
rect 14892 52986 14989 53042
rect 14892 52934 14904 52986
rect 14956 52934 14989 52986
rect 14892 52878 14989 52934
rect 14892 52826 14904 52878
rect 14956 52826 14989 52878
rect 14892 52576 14989 52826
rect 14892 51224 14902 52576
rect 14958 51224 14989 52576
rect 14892 49374 14989 51224
rect 14892 49322 14904 49374
rect 14956 49322 14989 49374
rect 14892 49266 14989 49322
rect 14892 49214 14904 49266
rect 14956 49214 14989 49266
rect 14892 49158 14989 49214
rect 14892 49106 14904 49158
rect 14956 49106 14989 49158
rect 14892 49050 14989 49106
rect 14892 48998 14904 49050
rect 14956 48998 14989 49050
rect 14892 48942 14989 48998
rect 14892 48890 14904 48942
rect 14956 48890 14989 48942
rect 14892 48834 14989 48890
rect 14892 48782 14904 48834
rect 14956 48782 14989 48834
rect 14892 48726 14989 48782
rect 14892 48674 14904 48726
rect 14956 48674 14989 48726
rect 14892 48618 14989 48674
rect 14892 48566 14904 48618
rect 14956 48566 14989 48618
rect 14892 48510 14989 48566
rect 14892 48458 14904 48510
rect 14956 48458 14989 48510
rect 14892 48402 14989 48458
rect 14892 48350 14904 48402
rect 14956 48350 14989 48402
rect 14892 48294 14989 48350
rect 14892 48242 14904 48294
rect 14956 48242 14989 48294
rect 14892 48186 14989 48242
rect 14892 48134 14904 48186
rect 14956 48134 14989 48186
rect 14892 48078 14989 48134
rect 14892 48026 14904 48078
rect 14956 48026 14989 48078
rect 14892 46174 14989 48026
rect 2798 44842 4734 46158
rect 5168 44842 7104 46158
rect 7874 44842 9810 46158
rect 10244 44842 12180 46158
rect 12861 44842 14673 46158
rect 14892 46122 14904 46174
rect 14956 46122 14989 46174
rect 14892 46066 14989 46122
rect 14892 46014 14904 46066
rect 14956 46014 14989 46066
rect 14892 45958 14989 46014
rect 14892 45906 14904 45958
rect 14956 45906 14989 45958
rect 14892 45850 14989 45906
rect 14892 45798 14904 45850
rect 14956 45798 14989 45850
rect 14892 45742 14989 45798
rect 14892 45690 14904 45742
rect 14956 45690 14989 45742
rect 14892 45634 14989 45690
rect 14892 45582 14904 45634
rect 14956 45582 14989 45634
rect 14892 45526 14989 45582
rect 14892 45474 14904 45526
rect 14956 45474 14989 45526
rect 14892 45418 14989 45474
rect 14892 45366 14904 45418
rect 14956 45366 14989 45418
rect 14892 45310 14989 45366
rect 14892 45258 14904 45310
rect 14956 45258 14989 45310
rect 14892 45202 14989 45258
rect 14892 45150 14904 45202
rect 14956 45150 14989 45202
rect 14892 45094 14989 45150
rect 14892 45042 14904 45094
rect 14956 45042 14989 45094
rect 14892 44986 14989 45042
rect 14892 44934 14904 44986
rect 14956 44934 14989 44986
rect 14892 44878 14989 44934
rect 14892 44826 14904 44878
rect 14956 44826 14989 44878
rect 2481 43242 2681 44558
rect 4851 43242 5051 44558
rect 7265 43242 7713 44558
rect 9927 43242 10127 44558
rect 12297 43242 12497 44558
rect 2481 41642 2681 42958
rect 4851 41642 5051 42958
rect 7265 41642 7713 42958
rect 9927 41642 10127 42958
rect 12297 41642 12497 42958
rect 2481 40042 2681 41358
rect 4851 40042 5051 41358
rect 7265 40042 7713 41358
rect 9927 40042 10127 41358
rect 12297 40042 12497 41358
rect 2292 39671 2302 39727
rect 2358 39671 2368 39727
rect 2292 39595 2368 39671
rect 2292 39539 2302 39595
rect 2358 39539 2368 39595
rect 2292 39463 2368 39539
rect 2292 39407 2302 39463
rect 2358 39407 2368 39463
rect 2292 39331 2368 39407
rect 2292 39275 2302 39331
rect 2358 39275 2368 39331
rect 2292 39199 2368 39275
rect 2292 39143 2302 39199
rect 2358 39143 2368 39199
rect 2292 39067 2368 39143
rect 2292 39011 2302 39067
rect 2358 39011 2368 39067
rect 2292 38935 2368 39011
rect 2292 38879 2302 38935
rect 2358 38879 2368 38935
rect 2292 38803 2368 38879
rect 2292 38747 2302 38803
rect 2358 38747 2368 38803
rect 2292 38671 2368 38747
rect 2292 38615 2302 38671
rect 2358 38615 2368 38671
rect 2292 38539 2368 38615
rect 2292 38483 2302 38539
rect 2358 38483 2368 38539
rect 2292 38400 2368 38483
rect -11 36824 20 38176
rect 76 36824 86 38176
rect 14892 38176 14989 44826
rect 2491 38098 2547 38154
rect 2615 38098 2671 38154
rect 4861 38098 4917 38154
rect 4985 38098 5041 38154
rect 7275 38098 7331 38154
rect 7399 38098 7455 38154
rect 7523 38098 7579 38154
rect 7647 38098 7703 38154
rect 9937 38098 9993 38154
rect 10061 38098 10117 38154
rect 12307 38098 12363 38154
rect 12431 38098 12487 38154
rect 2491 37974 2547 38030
rect 2615 37974 2671 38030
rect 4861 37974 4917 38030
rect 4985 37974 5041 38030
rect 7275 37974 7331 38030
rect 7399 37974 7455 38030
rect 7523 37974 7579 38030
rect 7647 37974 7703 38030
rect 9937 37974 9993 38030
rect 10061 37974 10117 38030
rect 12307 37974 12363 38030
rect 12431 37974 12487 38030
rect 2491 37850 2547 37906
rect 2615 37850 2671 37906
rect 4861 37850 4917 37906
rect 4985 37850 5041 37906
rect 7275 37850 7331 37906
rect 7399 37850 7455 37906
rect 7523 37850 7579 37906
rect 7647 37850 7703 37906
rect 9937 37850 9993 37906
rect 10061 37850 10117 37906
rect 12307 37850 12363 37906
rect 12431 37850 12487 37906
rect 2491 37726 2547 37782
rect 2615 37726 2671 37782
rect 4861 37726 4917 37782
rect 4985 37726 5041 37782
rect 7275 37726 7331 37782
rect 7399 37726 7455 37782
rect 7523 37726 7579 37782
rect 7647 37726 7703 37782
rect 9937 37726 9993 37782
rect 10061 37726 10117 37782
rect 12307 37726 12363 37782
rect 12431 37726 12487 37782
rect 2491 37602 2547 37658
rect 2615 37602 2671 37658
rect 4861 37602 4917 37658
rect 4985 37602 5041 37658
rect 7275 37602 7331 37658
rect 7399 37602 7455 37658
rect 7523 37602 7579 37658
rect 7647 37602 7703 37658
rect 9937 37602 9993 37658
rect 10061 37602 10117 37658
rect 12307 37602 12363 37658
rect 12431 37602 12487 37658
rect 2491 37478 2547 37534
rect 2615 37478 2671 37534
rect 4861 37478 4917 37534
rect 4985 37478 5041 37534
rect 7275 37478 7331 37534
rect 7399 37478 7455 37534
rect 7523 37478 7579 37534
rect 7647 37478 7703 37534
rect 9937 37478 9993 37534
rect 10061 37478 10117 37534
rect 12307 37478 12363 37534
rect 12431 37478 12487 37534
rect 2491 37354 2547 37410
rect 2615 37354 2671 37410
rect 4861 37354 4917 37410
rect 4985 37354 5041 37410
rect 7275 37354 7331 37410
rect 7399 37354 7455 37410
rect 7523 37354 7579 37410
rect 7647 37354 7703 37410
rect 9937 37354 9993 37410
rect 10061 37354 10117 37410
rect 12307 37354 12363 37410
rect 12431 37354 12487 37410
rect 2491 37230 2547 37286
rect 2615 37230 2671 37286
rect 4861 37230 4917 37286
rect 4985 37230 5041 37286
rect 7275 37230 7331 37286
rect 7399 37230 7455 37286
rect 7523 37230 7579 37286
rect 7647 37230 7703 37286
rect 9937 37230 9993 37286
rect 10061 37230 10117 37286
rect 12307 37230 12363 37286
rect 12431 37230 12487 37286
rect 2491 37106 2547 37162
rect 2615 37106 2671 37162
rect 4861 37106 4917 37162
rect 4985 37106 5041 37162
rect 7275 37106 7331 37162
rect 7399 37106 7455 37162
rect 7523 37106 7579 37162
rect 7647 37106 7703 37162
rect 9937 37106 9993 37162
rect 10061 37106 10117 37162
rect 12307 37106 12363 37162
rect 12431 37106 12487 37162
rect 2491 36982 2547 37038
rect 2615 36982 2671 37038
rect 4861 36982 4917 37038
rect 4985 36982 5041 37038
rect 7275 36982 7331 37038
rect 7399 36982 7455 37038
rect 7523 36982 7579 37038
rect 7647 36982 7703 37038
rect 9937 36982 9993 37038
rect 10061 36982 10117 37038
rect 12307 36982 12363 37038
rect 12431 36982 12487 37038
rect 2491 36858 2547 36914
rect 2615 36858 2671 36914
rect 4861 36858 4917 36914
rect 4985 36858 5041 36914
rect 7275 36858 7331 36914
rect 7399 36858 7455 36914
rect 7523 36858 7579 36914
rect 7647 36858 7703 36914
rect 9937 36858 9993 36914
rect 10061 36858 10117 36914
rect 12307 36858 12363 36914
rect 12431 36858 12487 36914
rect -11 36584 86 36824
rect -11 36532 22 36584
rect 74 36532 86 36584
rect 14892 36824 14902 38176
rect 14958 36824 14989 38176
rect 14892 36584 14989 36824
rect -11 36476 86 36532
rect -11 36424 22 36476
rect 74 36424 86 36476
rect -11 36368 86 36424
rect -11 36316 22 36368
rect 74 36316 86 36368
rect -11 36260 86 36316
rect -11 36208 22 36260
rect 74 36208 86 36260
rect -11 36152 86 36208
rect -11 36100 22 36152
rect 74 36100 86 36152
rect -11 36044 86 36100
rect -11 35992 22 36044
rect 74 35992 86 36044
rect -11 35936 86 35992
rect -11 35884 22 35936
rect 74 35884 86 35936
rect -11 35828 86 35884
rect -11 35776 22 35828
rect 74 35776 86 35828
rect -11 35720 86 35776
rect -11 35668 22 35720
rect 74 35668 86 35720
rect -11 35612 86 35668
rect -11 35560 22 35612
rect 74 35560 86 35612
rect -11 35504 86 35560
rect -11 35452 22 35504
rect 74 35452 86 35504
rect -11 35396 86 35452
rect -11 35344 22 35396
rect 74 35344 86 35396
rect -11 35288 86 35344
rect -11 35236 22 35288
rect 74 35236 86 35288
rect -11 35180 86 35236
rect -11 35128 22 35180
rect 74 35128 86 35180
rect -11 35072 86 35128
rect -11 35020 22 35072
rect 74 35020 86 35072
rect -11 34964 86 35020
rect -11 34912 22 34964
rect 74 34912 86 34964
rect -11 34856 86 34912
rect -11 34804 22 34856
rect 74 34804 86 34856
rect -11 34748 86 34804
rect -11 34696 22 34748
rect 74 34696 86 34748
rect -11 34640 86 34696
rect -11 34588 22 34640
rect 74 34588 86 34640
rect -11 34532 86 34588
rect -11 34480 22 34532
rect 74 34480 86 34532
rect -11 34424 86 34480
rect -11 34372 22 34424
rect 74 34372 86 34424
rect -11 34316 86 34372
rect -11 34264 22 34316
rect 74 34264 86 34316
rect -11 34208 86 34264
rect -11 34156 22 34208
rect 74 34156 86 34208
rect -11 34100 86 34156
rect -11 34048 22 34100
rect 74 34048 86 34100
rect -11 33992 86 34048
rect -11 33940 22 33992
rect 74 33940 86 33992
rect -11 33884 86 33940
rect -11 33832 22 33884
rect 74 33832 86 33884
rect -11 33776 86 33832
rect -11 33724 22 33776
rect 74 33724 86 33776
rect -11 33668 86 33724
rect -11 33616 22 33668
rect 74 33616 86 33668
rect 305 33636 2117 36564
rect 2798 33636 4734 36564
rect 5168 33636 7104 36564
rect 7874 33636 9810 36564
rect 10244 33636 12180 36564
rect 12861 33636 14673 36564
rect 14892 36532 14904 36584
rect 14956 36532 14989 36584
rect 14892 36476 14989 36532
rect 14892 36424 14904 36476
rect 14956 36424 14989 36476
rect 14892 36368 14989 36424
rect 14892 36316 14904 36368
rect 14956 36316 14989 36368
rect 14892 36260 14989 36316
rect 14892 36208 14904 36260
rect 14956 36208 14989 36260
rect 14892 36152 14989 36208
rect 14892 36100 14904 36152
rect 14956 36100 14989 36152
rect 14892 36044 14989 36100
rect 14892 35992 14904 36044
rect 14956 35992 14989 36044
rect 14892 35936 14989 35992
rect 14892 35884 14904 35936
rect 14956 35884 14989 35936
rect 14892 35828 14989 35884
rect 14892 35776 14904 35828
rect 14956 35776 14989 35828
rect 14892 35720 14989 35776
rect 14892 35668 14904 35720
rect 14956 35668 14989 35720
rect 14892 35612 14989 35668
rect 14892 35560 14904 35612
rect 14956 35560 14989 35612
rect 14892 35504 14989 35560
rect 14892 35452 14904 35504
rect 14956 35452 14989 35504
rect 14892 35396 14989 35452
rect 14892 35344 14904 35396
rect 14956 35344 14989 35396
rect 14892 35288 14989 35344
rect 14892 35236 14904 35288
rect 14956 35236 14989 35288
rect 14892 35180 14989 35236
rect 14892 35128 14904 35180
rect 14956 35128 14989 35180
rect 14892 35072 14989 35128
rect 14892 35020 14904 35072
rect 14956 35020 14989 35072
rect 14892 34964 14989 35020
rect 14892 34912 14904 34964
rect 14956 34912 14989 34964
rect 14892 34856 14989 34912
rect 14892 34804 14904 34856
rect 14956 34804 14989 34856
rect 14892 34748 14989 34804
rect 14892 34696 14904 34748
rect 14956 34696 14989 34748
rect 14892 34640 14989 34696
rect 14892 34588 14904 34640
rect 14956 34588 14989 34640
rect 14892 34532 14989 34588
rect 14892 34480 14904 34532
rect 14956 34480 14989 34532
rect 14892 34424 14989 34480
rect 14892 34372 14904 34424
rect 14956 34372 14989 34424
rect 14892 34316 14989 34372
rect 14892 34264 14904 34316
rect 14956 34264 14989 34316
rect 14892 34208 14989 34264
rect 14892 34156 14904 34208
rect 14956 34156 14989 34208
rect 14892 34100 14989 34156
rect 14892 34048 14904 34100
rect 14956 34048 14989 34100
rect 14892 33992 14989 34048
rect 14892 33940 14904 33992
rect 14956 33940 14989 33992
rect 14892 33884 14989 33940
rect 14892 33832 14904 33884
rect 14956 33832 14989 33884
rect 14892 33776 14989 33832
rect 14892 33724 14904 33776
rect 14956 33724 14989 33776
rect 14892 33668 14989 33724
rect -11 28574 86 33616
rect 14892 33616 14904 33668
rect 14956 33616 14989 33668
rect 2481 30436 2681 33364
rect 4851 30436 5051 33364
rect 7265 30436 7713 33364
rect 9927 30436 10127 33364
rect 12297 30436 12497 33364
rect 2481 28842 2681 30158
rect 4851 28842 5051 30158
rect 7265 28842 7713 30158
rect 9927 28842 10127 30158
rect 12297 28842 12497 30158
rect -11 28522 22 28574
rect 74 28522 86 28574
rect 14892 28574 14989 33616
rect -11 28466 86 28522
rect -11 28414 22 28466
rect 74 28414 86 28466
rect -11 28358 86 28414
rect -11 28306 22 28358
rect 74 28306 86 28358
rect -11 28250 86 28306
rect -11 28198 22 28250
rect 74 28198 86 28250
rect -11 28142 86 28198
rect -11 28090 22 28142
rect 74 28090 86 28142
rect -11 28034 86 28090
rect -11 27982 22 28034
rect 74 27982 86 28034
rect -11 27926 86 27982
rect -11 27874 22 27926
rect 74 27874 86 27926
rect -11 27818 86 27874
rect -11 27766 22 27818
rect 74 27766 86 27818
rect -11 27710 86 27766
rect -11 27658 22 27710
rect 74 27658 86 27710
rect -11 27602 86 27658
rect -11 27550 22 27602
rect 74 27550 86 27602
rect -11 27494 86 27550
rect -11 27442 22 27494
rect 74 27442 86 27494
rect -11 27386 86 27442
rect -11 27334 22 27386
rect 74 27334 86 27386
rect -11 27278 86 27334
rect -11 27226 22 27278
rect 74 27226 86 27278
rect 305 27242 2117 28558
rect 2798 27242 4734 28558
rect 5168 27242 7104 28558
rect 7874 27242 9810 28558
rect 10244 27242 12180 28558
rect 12861 27242 14673 28558
rect 14892 28522 14904 28574
rect 14956 28522 14989 28574
rect 14892 28466 14989 28522
rect 14892 28414 14904 28466
rect 14956 28414 14989 28466
rect 14892 28358 14989 28414
rect 14892 28306 14904 28358
rect 14956 28306 14989 28358
rect 14892 28250 14989 28306
rect 14892 28198 14904 28250
rect 14956 28198 14989 28250
rect 14892 28142 14989 28198
rect 14892 28090 14904 28142
rect 14956 28090 14989 28142
rect 14892 28034 14989 28090
rect 14892 27982 14904 28034
rect 14956 27982 14989 28034
rect 14892 27926 14989 27982
rect 14892 27874 14904 27926
rect 14956 27874 14989 27926
rect 14892 27818 14989 27874
rect 14892 27766 14904 27818
rect 14956 27766 14989 27818
rect 14892 27710 14989 27766
rect 14892 27658 14904 27710
rect 14956 27658 14989 27710
rect 14892 27602 14989 27658
rect 14892 27550 14904 27602
rect 14956 27550 14989 27602
rect 14892 27494 14989 27550
rect 14892 27442 14904 27494
rect 14956 27442 14989 27494
rect 14892 27386 14989 27442
rect 14892 27334 14904 27386
rect 14956 27334 14989 27386
rect 14892 27278 14989 27334
rect -11 14174 86 27226
rect 14892 27226 14904 27278
rect 14956 27226 14989 27278
rect 2481 24036 2681 26964
rect 4851 24036 5051 26964
rect 7265 24036 7713 26964
rect 9927 24036 10127 26964
rect 12297 24036 12497 26964
rect 2481 20836 2681 23764
rect 4851 20836 5051 23764
rect 7265 20836 7713 23764
rect 9927 20836 10127 23764
rect 12297 20836 12497 23764
rect 2481 17636 2681 20564
rect 4851 17636 5051 20564
rect 7265 17636 7713 20564
rect 9927 17636 10127 20564
rect 12297 17636 12497 20564
rect 2481 14436 2681 17364
rect 4851 14436 5051 17364
rect 7265 14436 7713 17364
rect 9927 14436 10127 17364
rect 12297 14436 12497 17364
rect -11 14122 22 14174
rect 74 14122 86 14174
rect 14892 14174 14989 27226
rect -11 14066 86 14122
rect -11 14014 22 14066
rect 74 14014 86 14066
rect -11 13958 86 14014
rect -11 13906 22 13958
rect 74 13906 86 13958
rect -11 13850 86 13906
rect -11 13798 22 13850
rect 74 13798 86 13850
rect -11 13742 86 13798
rect -11 13690 22 13742
rect 74 13690 86 13742
rect -11 13634 86 13690
rect -11 13582 22 13634
rect 74 13582 86 13634
rect -11 13526 86 13582
rect -11 13474 22 13526
rect 74 13474 86 13526
rect -11 13418 86 13474
rect -11 13366 22 13418
rect 74 13366 86 13418
rect -11 13310 86 13366
rect -11 13258 22 13310
rect 74 13258 86 13310
rect -11 13202 86 13258
rect -11 13150 22 13202
rect 74 13150 86 13202
rect -11 13094 86 13150
rect -11 13042 22 13094
rect 74 13042 86 13094
rect -11 12986 86 13042
rect -11 12934 22 12986
rect 74 12934 86 12986
rect -11 12878 86 12934
rect -11 12826 22 12878
rect 74 12826 86 12878
rect 305 12842 2117 14158
rect 2798 12842 4734 14158
rect 5168 12842 7104 14158
rect 7874 12842 9810 14158
rect 10244 12842 12180 14158
rect 12861 12842 14673 14158
rect 14892 14122 14904 14174
rect 14956 14122 14989 14174
rect 14892 14066 14989 14122
rect 14892 14014 14904 14066
rect 14956 14014 14989 14066
rect 14892 13958 14989 14014
rect 14892 13906 14904 13958
rect 14956 13906 14989 13958
rect 14892 13850 14989 13906
rect 14892 13798 14904 13850
rect 14956 13798 14989 13850
rect 14892 13742 14989 13798
rect 14892 13690 14904 13742
rect 14956 13690 14989 13742
rect 14892 13634 14989 13690
rect 14892 13582 14904 13634
rect 14956 13582 14989 13634
rect 14892 13526 14989 13582
rect 14892 13474 14904 13526
rect 14956 13474 14989 13526
rect 14892 13418 14989 13474
rect 14892 13366 14904 13418
rect 14956 13366 14989 13418
rect 14892 13310 14989 13366
rect 14892 13258 14904 13310
rect 14956 13258 14989 13310
rect 14892 13202 14989 13258
rect 14892 13150 14904 13202
rect 14956 13150 14989 13202
rect 14892 13094 14989 13150
rect 14892 13042 14904 13094
rect 14956 13042 14989 13094
rect 14892 12986 14989 13042
rect 14892 12934 14904 12986
rect 14956 12934 14989 12986
rect 14892 12878 14989 12934
rect -11 10984 86 12826
rect 14892 12826 14904 12878
rect 14956 12826 14989 12878
rect 2481 11242 2681 12558
rect 4851 11242 5051 12558
rect 7265 11242 7713 12558
rect 9927 11242 10127 12558
rect 12297 11242 12497 12558
rect -11 10932 22 10984
rect 74 10932 86 10984
rect 14892 10984 14989 12826
rect -11 10876 86 10932
rect -11 10824 22 10876
rect 74 10824 86 10876
rect -11 10768 86 10824
rect -11 10716 22 10768
rect 74 10716 86 10768
rect -11 10660 86 10716
rect -11 10608 22 10660
rect 74 10608 86 10660
rect -11 10552 86 10608
rect -11 10500 22 10552
rect 74 10500 86 10552
rect -11 10444 86 10500
rect -11 10392 22 10444
rect 74 10392 86 10444
rect -11 10336 86 10392
rect -11 10284 22 10336
rect 74 10284 86 10336
rect -11 10228 86 10284
rect -11 10176 22 10228
rect 74 10176 86 10228
rect -11 10120 86 10176
rect -11 10068 22 10120
rect 74 10068 86 10120
rect -11 10012 86 10068
rect -11 9960 22 10012
rect 74 9960 86 10012
rect -11 9904 86 9960
rect -11 9852 22 9904
rect 74 9852 86 9904
rect -11 9796 86 9852
rect -11 9744 22 9796
rect 74 9744 86 9796
rect -11 9688 86 9744
rect -11 9636 22 9688
rect 74 9636 86 9688
rect -11 9580 86 9636
rect -11 9528 22 9580
rect 74 9528 86 9580
rect -11 9472 86 9528
rect -11 9420 22 9472
rect 74 9420 86 9472
rect -11 9364 86 9420
rect -11 9312 22 9364
rect 74 9312 86 9364
rect -11 9256 86 9312
rect -11 9204 22 9256
rect 74 9204 86 9256
rect -11 9148 86 9204
rect -11 9096 22 9148
rect 74 9096 86 9148
rect -11 9040 86 9096
rect -11 8988 22 9040
rect 74 8988 86 9040
rect -11 8932 86 8988
rect -11 8880 22 8932
rect 74 8880 86 8932
rect -11 8824 86 8880
rect -11 8772 22 8824
rect 74 8772 86 8824
rect -11 8716 86 8772
rect -11 8664 22 8716
rect 74 8664 86 8716
rect -11 8608 86 8664
rect -11 8556 22 8608
rect 74 8556 86 8608
rect -11 8500 86 8556
rect -11 8448 22 8500
rect 74 8448 86 8500
rect -11 8392 86 8448
rect -11 8340 22 8392
rect 74 8340 86 8392
rect -11 8284 86 8340
rect -11 8232 22 8284
rect 74 8232 86 8284
rect -11 8176 86 8232
rect -11 8124 22 8176
rect 74 8124 86 8176
rect -11 8068 86 8124
rect -11 8016 22 8068
rect 74 8016 86 8068
rect 305 8036 2117 10964
rect 2798 8036 4734 10964
rect 5168 8036 7104 10964
rect 7874 8036 9810 10964
rect 10244 8036 12180 10964
rect 12861 8036 14673 10964
rect 14892 10932 14904 10984
rect 14956 10932 14989 10984
rect 14892 10876 14989 10932
rect 14892 10824 14904 10876
rect 14956 10824 14989 10876
rect 14892 10768 14989 10824
rect 14892 10716 14904 10768
rect 14956 10716 14989 10768
rect 14892 10660 14989 10716
rect 14892 10608 14904 10660
rect 14956 10608 14989 10660
rect 14892 10552 14989 10608
rect 14892 10500 14904 10552
rect 14956 10500 14989 10552
rect 14892 10444 14989 10500
rect 14892 10392 14904 10444
rect 14956 10392 14989 10444
rect 14892 10336 14989 10392
rect 14892 10284 14904 10336
rect 14956 10284 14989 10336
rect 14892 10228 14989 10284
rect 14892 10176 14904 10228
rect 14956 10176 14989 10228
rect 14892 10120 14989 10176
rect 14892 10068 14904 10120
rect 14956 10068 14989 10120
rect 14892 10012 14989 10068
rect 14892 9960 14904 10012
rect 14956 9960 14989 10012
rect 14892 9904 14989 9960
rect 14892 9852 14904 9904
rect 14956 9852 14989 9904
rect 14892 9796 14989 9852
rect 14892 9744 14904 9796
rect 14956 9744 14989 9796
rect 14892 9688 14989 9744
rect 14892 9636 14904 9688
rect 14956 9636 14989 9688
rect 14892 9580 14989 9636
rect 14892 9528 14904 9580
rect 14956 9528 14989 9580
rect 14892 9472 14989 9528
rect 14892 9420 14904 9472
rect 14956 9420 14989 9472
rect 14892 9364 14989 9420
rect 14892 9312 14904 9364
rect 14956 9312 14989 9364
rect 14892 9256 14989 9312
rect 14892 9204 14904 9256
rect 14956 9204 14989 9256
rect 14892 9148 14989 9204
rect 14892 9096 14904 9148
rect 14956 9096 14989 9148
rect 14892 9040 14989 9096
rect 14892 8988 14904 9040
rect 14956 8988 14989 9040
rect 14892 8932 14989 8988
rect 14892 8880 14904 8932
rect 14956 8880 14989 8932
rect 14892 8824 14989 8880
rect 14892 8772 14904 8824
rect 14956 8772 14989 8824
rect 14892 8716 14989 8772
rect 14892 8664 14904 8716
rect 14956 8664 14989 8716
rect 14892 8608 14989 8664
rect 14892 8556 14904 8608
rect 14956 8556 14989 8608
rect 14892 8500 14989 8556
rect 14892 8448 14904 8500
rect 14956 8448 14989 8500
rect 14892 8392 14989 8448
rect 14892 8340 14904 8392
rect 14956 8340 14989 8392
rect 14892 8284 14989 8340
rect 14892 8232 14904 8284
rect 14956 8232 14989 8284
rect 14892 8176 14989 8232
rect 14892 8124 14904 8176
rect 14956 8124 14989 8176
rect 14892 8068 14989 8124
rect -11 7784 86 8016
rect -11 7732 22 7784
rect 74 7732 86 7784
rect 14892 8016 14904 8068
rect 14956 8016 14989 8068
rect 14892 7784 14989 8016
rect -11 7676 86 7732
rect -11 7624 22 7676
rect 74 7624 86 7676
rect -11 7568 86 7624
rect -11 7516 22 7568
rect 74 7516 86 7568
rect -11 7460 86 7516
rect -11 7408 22 7460
rect 74 7408 86 7460
rect -11 7352 86 7408
rect -11 7300 22 7352
rect 74 7300 86 7352
rect -11 7244 86 7300
rect -11 7192 22 7244
rect 74 7192 86 7244
rect -11 7136 86 7192
rect -11 7084 22 7136
rect 74 7084 86 7136
rect -11 7028 86 7084
rect -11 6976 22 7028
rect 74 6976 86 7028
rect -11 6920 86 6976
rect -11 6868 22 6920
rect 74 6868 86 6920
rect -11 6812 86 6868
rect -11 6760 22 6812
rect 74 6760 86 6812
rect -11 6704 86 6760
rect -11 6652 22 6704
rect 74 6652 86 6704
rect -11 6596 86 6652
rect -11 6544 22 6596
rect 74 6544 86 6596
rect -11 6488 86 6544
rect -11 6436 22 6488
rect 74 6436 86 6488
rect -11 6380 86 6436
rect -11 6328 22 6380
rect 74 6328 86 6380
rect -11 6272 86 6328
rect -11 6220 22 6272
rect 74 6220 86 6272
rect -11 6164 86 6220
rect -11 6112 22 6164
rect 74 6112 86 6164
rect -11 6056 86 6112
rect -11 6004 22 6056
rect 74 6004 86 6056
rect -11 5948 86 6004
rect -11 5896 22 5948
rect 74 5896 86 5948
rect -11 5840 86 5896
rect -11 5788 22 5840
rect 74 5788 86 5840
rect -11 5732 86 5788
rect -11 5680 22 5732
rect 74 5680 86 5732
rect -11 5624 86 5680
rect -11 5572 22 5624
rect 74 5572 86 5624
rect -11 5516 86 5572
rect -11 5464 22 5516
rect 74 5464 86 5516
rect -11 5408 86 5464
rect -11 5356 22 5408
rect 74 5356 86 5408
rect -11 5300 86 5356
rect -11 5248 22 5300
rect 74 5248 86 5300
rect -11 5192 86 5248
rect -11 5140 22 5192
rect 74 5140 86 5192
rect -11 5084 86 5140
rect -11 5032 22 5084
rect 74 5032 86 5084
rect -11 4976 86 5032
rect -11 4924 22 4976
rect 74 4924 86 4976
rect -11 4868 86 4924
rect -11 4816 22 4868
rect 74 4816 86 4868
rect 305 4836 2117 7764
rect 2798 4836 4734 7764
rect 5168 4836 7104 7764
rect 7874 4836 9810 7764
rect 10244 4836 12180 7764
rect 12861 4836 14673 7764
rect 14892 7732 14904 7784
rect 14956 7732 14989 7784
rect 14892 7676 14989 7732
rect 14892 7624 14904 7676
rect 14956 7624 14989 7676
rect 14892 7568 14989 7624
rect 14892 7516 14904 7568
rect 14956 7516 14989 7568
rect 14892 7460 14989 7516
rect 14892 7408 14904 7460
rect 14956 7408 14989 7460
rect 14892 7352 14989 7408
rect 14892 7300 14904 7352
rect 14956 7300 14989 7352
rect 14892 7244 14989 7300
rect 14892 7192 14904 7244
rect 14956 7192 14989 7244
rect 14892 7136 14989 7192
rect 14892 7084 14904 7136
rect 14956 7084 14989 7136
rect 14892 7028 14989 7084
rect 14892 6976 14904 7028
rect 14956 6976 14989 7028
rect 14892 6920 14989 6976
rect 14892 6868 14904 6920
rect 14956 6868 14989 6920
rect 14892 6812 14989 6868
rect 14892 6760 14904 6812
rect 14956 6760 14989 6812
rect 14892 6704 14989 6760
rect 14892 6652 14904 6704
rect 14956 6652 14989 6704
rect 14892 6596 14989 6652
rect 14892 6544 14904 6596
rect 14956 6544 14989 6596
rect 14892 6488 14989 6544
rect 14892 6436 14904 6488
rect 14956 6436 14989 6488
rect 14892 6380 14989 6436
rect 14892 6328 14904 6380
rect 14956 6328 14989 6380
rect 14892 6272 14989 6328
rect 14892 6220 14904 6272
rect 14956 6220 14989 6272
rect 14892 6164 14989 6220
rect 14892 6112 14904 6164
rect 14956 6112 14989 6164
rect 14892 6056 14989 6112
rect 14892 6004 14904 6056
rect 14956 6004 14989 6056
rect 14892 5948 14989 6004
rect 14892 5896 14904 5948
rect 14956 5896 14989 5948
rect 14892 5840 14989 5896
rect 14892 5788 14904 5840
rect 14956 5788 14989 5840
rect 14892 5732 14989 5788
rect 14892 5680 14904 5732
rect 14956 5680 14989 5732
rect 14892 5624 14989 5680
rect 14892 5572 14904 5624
rect 14956 5572 14989 5624
rect 14892 5516 14989 5572
rect 14892 5464 14904 5516
rect 14956 5464 14989 5516
rect 14892 5408 14989 5464
rect 14892 5356 14904 5408
rect 14956 5356 14989 5408
rect 14892 5300 14989 5356
rect 14892 5248 14904 5300
rect 14956 5248 14989 5300
rect 14892 5192 14989 5248
rect 14892 5140 14904 5192
rect 14956 5140 14989 5192
rect 14892 5084 14989 5140
rect 14892 5032 14904 5084
rect 14956 5032 14989 5084
rect 14892 4976 14989 5032
rect 14892 4924 14904 4976
rect 14956 4924 14989 4976
rect 14892 4868 14989 4924
rect -11 4584 86 4816
rect -11 4532 22 4584
rect 74 4532 86 4584
rect 14892 4816 14904 4868
rect 14956 4816 14989 4868
rect 14892 4584 14989 4816
rect -11 4476 86 4532
rect -11 4424 22 4476
rect 74 4424 86 4476
rect -11 4368 86 4424
rect -11 4316 22 4368
rect 74 4316 86 4368
rect -11 4260 86 4316
rect -11 4208 22 4260
rect 74 4208 86 4260
rect -11 4152 86 4208
rect -11 4100 22 4152
rect 74 4100 86 4152
rect -11 4044 86 4100
rect -11 3992 22 4044
rect 74 3992 86 4044
rect -11 3936 86 3992
rect -11 3884 22 3936
rect 74 3884 86 3936
rect -11 3828 86 3884
rect -11 3776 22 3828
rect 74 3776 86 3828
rect -11 3720 86 3776
rect -11 3668 22 3720
rect 74 3668 86 3720
rect -11 3612 86 3668
rect -11 3560 22 3612
rect 74 3560 86 3612
rect -11 3504 86 3560
rect -11 3452 22 3504
rect 74 3452 86 3504
rect -11 3396 86 3452
rect -11 3344 22 3396
rect 74 3344 86 3396
rect -11 3288 86 3344
rect -11 3236 22 3288
rect 74 3236 86 3288
rect -11 3180 86 3236
rect -11 3128 22 3180
rect 74 3128 86 3180
rect -11 3072 86 3128
rect -11 3020 22 3072
rect 74 3020 86 3072
rect -11 2964 86 3020
rect -11 2912 22 2964
rect 74 2912 86 2964
rect -11 2856 86 2912
rect -11 2804 22 2856
rect 74 2804 86 2856
rect -11 2748 86 2804
rect -11 2696 22 2748
rect 74 2696 86 2748
rect -11 2640 86 2696
rect -11 2588 22 2640
rect 74 2588 86 2640
rect -11 2532 86 2588
rect -11 2480 22 2532
rect 74 2480 86 2532
rect -11 2424 86 2480
rect -11 2372 22 2424
rect 74 2372 86 2424
rect -11 2316 86 2372
rect -11 2264 22 2316
rect 74 2264 86 2316
rect -11 2208 86 2264
rect -11 2156 22 2208
rect 74 2156 86 2208
rect -11 2100 86 2156
rect -11 2048 22 2100
rect 74 2048 86 2100
rect -11 1992 86 2048
rect -11 1940 22 1992
rect 74 1940 86 1992
rect -11 1884 86 1940
rect -11 1832 22 1884
rect 74 1832 86 1884
rect -11 1776 86 1832
rect -11 1724 22 1776
rect 74 1724 86 1776
rect -11 1668 86 1724
rect -11 1616 22 1668
rect 74 1616 86 1668
rect 305 1636 2117 4564
rect 2798 1636 4734 4564
rect 5168 1636 7104 4564
rect 7874 1636 9810 4564
rect 10244 1636 12180 4564
rect 12861 1636 14673 4564
rect 14892 4532 14904 4584
rect 14956 4532 14989 4584
rect 14892 4476 14989 4532
rect 14892 4424 14904 4476
rect 14956 4424 14989 4476
rect 14892 4368 14989 4424
rect 14892 4316 14904 4368
rect 14956 4316 14989 4368
rect 14892 4260 14989 4316
rect 14892 4208 14904 4260
rect 14956 4208 14989 4260
rect 14892 4152 14989 4208
rect 14892 4100 14904 4152
rect 14956 4100 14989 4152
rect 14892 4044 14989 4100
rect 14892 3992 14904 4044
rect 14956 3992 14989 4044
rect 14892 3936 14989 3992
rect 14892 3884 14904 3936
rect 14956 3884 14989 3936
rect 14892 3828 14989 3884
rect 14892 3776 14904 3828
rect 14956 3776 14989 3828
rect 14892 3720 14989 3776
rect 14892 3668 14904 3720
rect 14956 3668 14989 3720
rect 14892 3612 14989 3668
rect 14892 3560 14904 3612
rect 14956 3560 14989 3612
rect 14892 3504 14989 3560
rect 14892 3452 14904 3504
rect 14956 3452 14989 3504
rect 14892 3396 14989 3452
rect 14892 3344 14904 3396
rect 14956 3344 14989 3396
rect 14892 3288 14989 3344
rect 14892 3236 14904 3288
rect 14956 3236 14989 3288
rect 14892 3180 14989 3236
rect 14892 3128 14904 3180
rect 14956 3128 14989 3180
rect 14892 3072 14989 3128
rect 14892 3020 14904 3072
rect 14956 3020 14989 3072
rect 14892 2964 14989 3020
rect 14892 2912 14904 2964
rect 14956 2912 14989 2964
rect 14892 2856 14989 2912
rect 14892 2804 14904 2856
rect 14956 2804 14989 2856
rect 14892 2748 14989 2804
rect 14892 2696 14904 2748
rect 14956 2696 14989 2748
rect 14892 2640 14989 2696
rect 14892 2588 14904 2640
rect 14956 2588 14989 2640
rect 14892 2532 14989 2588
rect 14892 2480 14904 2532
rect 14956 2480 14989 2532
rect 14892 2424 14989 2480
rect 14892 2372 14904 2424
rect 14956 2372 14989 2424
rect 14892 2316 14989 2372
rect 14892 2264 14904 2316
rect 14956 2264 14989 2316
rect 14892 2208 14989 2264
rect 14892 2156 14904 2208
rect 14956 2156 14989 2208
rect 14892 2100 14989 2156
rect 14892 2048 14904 2100
rect 14956 2048 14989 2100
rect 14892 1992 14989 2048
rect 14892 1940 14904 1992
rect 14956 1940 14989 1992
rect 14892 1884 14989 1940
rect 14892 1832 14904 1884
rect 14956 1832 14989 1884
rect 14892 1776 14989 1832
rect 14892 1724 14904 1776
rect 14956 1724 14989 1776
rect 14892 1668 14989 1724
rect -11 1604 86 1616
rect 14892 1616 14904 1668
rect 14956 1616 14989 1668
rect 14892 1604 14989 1616
rect 261 0 2161 1190
rect 2741 0 4791 1190
rect 5111 0 7161 1190
rect 7817 0 9867 1190
rect 10187 0 12237 1190
rect 12817 0 14717 1190
<< via2 >>
rect 20 52574 76 52576
rect 20 52522 22 52574
rect 22 52522 74 52574
rect 74 52522 76 52574
rect 20 52466 76 52522
rect 20 52414 22 52466
rect 22 52414 74 52466
rect 74 52414 76 52466
rect 20 52358 76 52414
rect 20 52306 22 52358
rect 22 52306 74 52358
rect 74 52306 76 52358
rect 20 52250 76 52306
rect 20 52198 22 52250
rect 22 52198 74 52250
rect 74 52198 76 52250
rect 20 52142 76 52198
rect 20 52090 22 52142
rect 22 52090 74 52142
rect 74 52090 76 52142
rect 20 52034 76 52090
rect 20 51982 22 52034
rect 22 51982 74 52034
rect 74 51982 76 52034
rect 20 51926 76 51982
rect 20 51874 22 51926
rect 22 51874 74 51926
rect 74 51874 76 51926
rect 20 51818 76 51874
rect 20 51766 22 51818
rect 22 51766 74 51818
rect 74 51766 76 51818
rect 20 51710 76 51766
rect 20 51658 22 51710
rect 22 51658 74 51710
rect 74 51658 76 51710
rect 20 51602 76 51658
rect 20 51550 22 51602
rect 22 51550 74 51602
rect 74 51550 76 51602
rect 20 51494 76 51550
rect 20 51442 22 51494
rect 22 51442 74 51494
rect 74 51442 76 51494
rect 20 51386 76 51442
rect 20 51334 22 51386
rect 22 51334 74 51386
rect 74 51334 76 51386
rect 20 51278 76 51334
rect 20 51226 22 51278
rect 22 51226 74 51278
rect 74 51226 76 51278
rect 20 51224 76 51226
rect 315 52492 371 52548
rect 439 52492 495 52548
rect 563 52492 619 52548
rect 687 52492 743 52548
rect 811 52492 867 52548
rect 935 52492 991 52548
rect 1059 52492 1115 52548
rect 1183 52492 1239 52548
rect 1307 52492 1363 52548
rect 1431 52492 1487 52548
rect 1555 52492 1611 52548
rect 1679 52492 1735 52548
rect 1803 52492 1859 52548
rect 1927 52492 1983 52548
rect 2051 52492 2107 52548
rect 315 52368 371 52424
rect 439 52368 495 52424
rect 563 52368 619 52424
rect 687 52368 743 52424
rect 811 52368 867 52424
rect 935 52368 991 52424
rect 1059 52368 1115 52424
rect 1183 52368 1239 52424
rect 1307 52368 1363 52424
rect 1431 52368 1487 52424
rect 1555 52368 1611 52424
rect 1679 52368 1735 52424
rect 1803 52368 1859 52424
rect 1927 52368 1983 52424
rect 2051 52368 2107 52424
rect 315 52244 371 52300
rect 439 52244 495 52300
rect 563 52244 619 52300
rect 687 52244 743 52300
rect 811 52244 867 52300
rect 935 52244 991 52300
rect 1059 52244 1115 52300
rect 1183 52244 1239 52300
rect 1307 52244 1363 52300
rect 1431 52244 1487 52300
rect 1555 52244 1611 52300
rect 1679 52244 1735 52300
rect 1803 52244 1859 52300
rect 1927 52244 1983 52300
rect 2051 52244 2107 52300
rect 315 52120 371 52176
rect 439 52120 495 52176
rect 563 52120 619 52176
rect 687 52120 743 52176
rect 811 52120 867 52176
rect 935 52120 991 52176
rect 1059 52120 1115 52176
rect 1183 52120 1239 52176
rect 1307 52120 1363 52176
rect 1431 52120 1487 52176
rect 1555 52120 1611 52176
rect 1679 52120 1735 52176
rect 1803 52120 1859 52176
rect 1927 52120 1983 52176
rect 2051 52120 2107 52176
rect 315 51996 371 52052
rect 439 51996 495 52052
rect 563 51996 619 52052
rect 687 51996 743 52052
rect 811 51996 867 52052
rect 935 51996 991 52052
rect 1059 51996 1115 52052
rect 1183 51996 1239 52052
rect 1307 51996 1363 52052
rect 1431 51996 1487 52052
rect 1555 51996 1611 52052
rect 1679 51996 1735 52052
rect 1803 51996 1859 52052
rect 1927 51996 1983 52052
rect 2051 51996 2107 52052
rect 315 51872 371 51928
rect 439 51872 495 51928
rect 563 51872 619 51928
rect 687 51872 743 51928
rect 811 51872 867 51928
rect 935 51872 991 51928
rect 1059 51872 1115 51928
rect 1183 51872 1239 51928
rect 1307 51872 1363 51928
rect 1431 51872 1487 51928
rect 1555 51872 1611 51928
rect 1679 51872 1735 51928
rect 1803 51872 1859 51928
rect 1927 51872 1983 51928
rect 2051 51872 2107 51928
rect 315 51748 371 51804
rect 439 51748 495 51804
rect 563 51748 619 51804
rect 687 51748 743 51804
rect 811 51748 867 51804
rect 935 51748 991 51804
rect 1059 51748 1115 51804
rect 1183 51748 1239 51804
rect 1307 51748 1363 51804
rect 1431 51748 1487 51804
rect 1555 51748 1611 51804
rect 1679 51748 1735 51804
rect 1803 51748 1859 51804
rect 1927 51748 1983 51804
rect 2051 51748 2107 51804
rect 315 51624 371 51680
rect 439 51624 495 51680
rect 563 51624 619 51680
rect 687 51624 743 51680
rect 811 51624 867 51680
rect 935 51624 991 51680
rect 1059 51624 1115 51680
rect 1183 51624 1239 51680
rect 1307 51624 1363 51680
rect 1431 51624 1487 51680
rect 1555 51624 1611 51680
rect 1679 51624 1735 51680
rect 1803 51624 1859 51680
rect 1927 51624 1983 51680
rect 2051 51624 2107 51680
rect 315 51500 371 51556
rect 439 51500 495 51556
rect 563 51500 619 51556
rect 687 51500 743 51556
rect 811 51500 867 51556
rect 935 51500 991 51556
rect 1059 51500 1115 51556
rect 1183 51500 1239 51556
rect 1307 51500 1363 51556
rect 1431 51500 1487 51556
rect 1555 51500 1611 51556
rect 1679 51500 1735 51556
rect 1803 51500 1859 51556
rect 1927 51500 1983 51556
rect 2051 51500 2107 51556
rect 315 51376 371 51432
rect 439 51376 495 51432
rect 563 51376 619 51432
rect 687 51376 743 51432
rect 811 51376 867 51432
rect 935 51376 991 51432
rect 1059 51376 1115 51432
rect 1183 51376 1239 51432
rect 1307 51376 1363 51432
rect 1431 51376 1487 51432
rect 1555 51376 1611 51432
rect 1679 51376 1735 51432
rect 1803 51376 1859 51432
rect 1927 51376 1983 51432
rect 2051 51376 2107 51432
rect 315 51252 371 51308
rect 439 51252 495 51308
rect 563 51252 619 51308
rect 687 51252 743 51308
rect 811 51252 867 51308
rect 935 51252 991 51308
rect 1059 51252 1115 51308
rect 1183 51252 1239 51308
rect 1307 51252 1363 51308
rect 1431 51252 1487 51308
rect 1555 51252 1611 51308
rect 1679 51252 1735 51308
rect 1803 51252 1859 51308
rect 1927 51252 1983 51308
rect 2051 51252 2107 51308
rect 2302 50870 2358 50926
rect 2302 50738 2358 50794
rect 2302 50606 2358 50662
rect 2302 50474 2358 50530
rect 2302 50342 2358 50398
rect 2302 50210 2358 50266
rect 2302 50078 2358 50134
rect 2302 49946 2358 50002
rect 2302 49814 2358 49870
rect 2302 49682 2358 49738
rect 2491 50892 2547 50948
rect 2615 50922 2642 50948
rect 2642 50922 2671 50948
rect 2615 50892 2671 50922
rect 2491 50768 2547 50824
rect 2615 50814 2642 50824
rect 2642 50814 2671 50824
rect 2615 50768 2671 50814
rect 2491 50644 2547 50700
rect 2615 50650 2671 50700
rect 2615 50644 2642 50650
rect 2642 50644 2671 50650
rect 2491 50520 2547 50576
rect 2615 50542 2671 50576
rect 2615 50520 2642 50542
rect 2642 50520 2671 50542
rect 2491 50396 2547 50452
rect 2615 50434 2671 50452
rect 2615 50396 2642 50434
rect 2642 50396 2671 50434
rect 2491 50272 2547 50328
rect 2615 50326 2671 50328
rect 2615 50274 2642 50326
rect 2642 50274 2671 50326
rect 2615 50272 2671 50274
rect 2491 50148 2547 50204
rect 2615 50166 2642 50204
rect 2642 50166 2671 50204
rect 2615 50148 2671 50166
rect 2491 50024 2547 50080
rect 2615 50058 2642 50080
rect 2642 50058 2671 50080
rect 2615 50024 2671 50058
rect 2491 49900 2547 49956
rect 2615 49950 2642 49956
rect 2642 49950 2671 49956
rect 2615 49900 2671 49950
rect 2491 49776 2547 49832
rect 2615 49786 2671 49832
rect 2615 49776 2642 49786
rect 2642 49776 2671 49786
rect 2491 49652 2547 49708
rect 2615 49678 2671 49708
rect 2615 49652 2642 49678
rect 2642 49652 2671 49678
rect 2808 52492 2864 52548
rect 2932 52492 2988 52548
rect 3056 52492 3112 52548
rect 3180 52492 3236 52548
rect 3304 52492 3360 52548
rect 3428 52492 3484 52548
rect 3552 52492 3608 52548
rect 3676 52492 3732 52548
rect 3800 52492 3856 52548
rect 3924 52492 3980 52548
rect 4048 52492 4104 52548
rect 4172 52492 4228 52548
rect 4296 52492 4352 52548
rect 4420 52492 4476 52548
rect 4544 52492 4600 52548
rect 4668 52492 4724 52548
rect 2808 52368 2864 52424
rect 2932 52368 2988 52424
rect 3056 52368 3112 52424
rect 3180 52368 3236 52424
rect 3304 52368 3360 52424
rect 3428 52368 3484 52424
rect 3552 52368 3608 52424
rect 3676 52368 3732 52424
rect 3800 52368 3856 52424
rect 3924 52368 3980 52424
rect 4048 52368 4104 52424
rect 4172 52368 4228 52424
rect 4296 52368 4352 52424
rect 4420 52368 4476 52424
rect 4544 52368 4600 52424
rect 4668 52368 4724 52424
rect 2808 52244 2864 52300
rect 2932 52244 2988 52300
rect 3056 52244 3112 52300
rect 3180 52244 3236 52300
rect 3304 52244 3360 52300
rect 3428 52244 3484 52300
rect 3552 52244 3608 52300
rect 3676 52244 3732 52300
rect 3800 52244 3856 52300
rect 3924 52244 3980 52300
rect 4048 52244 4104 52300
rect 4172 52244 4228 52300
rect 4296 52244 4352 52300
rect 4420 52244 4476 52300
rect 4544 52244 4600 52300
rect 4668 52244 4724 52300
rect 2808 52120 2864 52176
rect 2932 52120 2988 52176
rect 3056 52120 3112 52176
rect 3180 52120 3236 52176
rect 3304 52120 3360 52176
rect 3428 52120 3484 52176
rect 3552 52120 3608 52176
rect 3676 52120 3732 52176
rect 3800 52120 3856 52176
rect 3924 52120 3980 52176
rect 4048 52120 4104 52176
rect 4172 52120 4228 52176
rect 4296 52120 4352 52176
rect 4420 52120 4476 52176
rect 4544 52120 4600 52176
rect 4668 52120 4724 52176
rect 2808 51996 2864 52052
rect 2932 51996 2988 52052
rect 3056 51996 3112 52052
rect 3180 52009 3236 52052
rect 3304 52009 3360 52052
rect 3428 52009 3484 52052
rect 3552 52009 3608 52052
rect 3676 52009 3732 52052
rect 3800 52009 3856 52052
rect 3924 52009 3980 52052
rect 4048 52009 4104 52052
rect 4172 52009 4228 52052
rect 4296 52009 4352 52052
rect 4420 52009 4476 52052
rect 4544 52009 4600 52052
rect 4668 52009 4724 52052
rect 3180 51996 3213 52009
rect 3213 51996 3236 52009
rect 3304 51996 3321 52009
rect 3321 51996 3360 52009
rect 3428 51996 3429 52009
rect 3429 51996 3484 52009
rect 3552 51996 3593 52009
rect 3593 51996 3608 52009
rect 3676 51996 3701 52009
rect 3701 51996 3732 52009
rect 3800 51996 3809 52009
rect 3809 51996 3856 52009
rect 3924 51996 3969 52009
rect 3969 51996 3980 52009
rect 4048 51996 4077 52009
rect 4077 51996 4104 52009
rect 4172 51996 4185 52009
rect 4185 51996 4228 52009
rect 4296 51996 4349 52009
rect 4349 51996 4352 52009
rect 4420 51996 4457 52009
rect 4457 51996 4476 52009
rect 4544 51996 4565 52009
rect 4565 51996 4600 52009
rect 4668 51996 4673 52009
rect 4673 51996 4724 52009
rect 2808 51872 2864 51928
rect 2932 51872 2988 51928
rect 3056 51872 3112 51928
rect 3180 51901 3236 51928
rect 3304 51901 3360 51928
rect 3428 51901 3484 51928
rect 3552 51901 3608 51928
rect 3676 51901 3732 51928
rect 3800 51901 3856 51928
rect 3924 51901 3980 51928
rect 4048 51901 4104 51928
rect 4172 51901 4228 51928
rect 4296 51901 4352 51928
rect 4420 51901 4476 51928
rect 4544 51901 4600 51928
rect 4668 51901 4724 51928
rect 3180 51872 3213 51901
rect 3213 51872 3236 51901
rect 3304 51872 3321 51901
rect 3321 51872 3360 51901
rect 3428 51872 3429 51901
rect 3429 51872 3484 51901
rect 3552 51872 3593 51901
rect 3593 51872 3608 51901
rect 3676 51872 3701 51901
rect 3701 51872 3732 51901
rect 3800 51872 3809 51901
rect 3809 51872 3856 51901
rect 3924 51872 3969 51901
rect 3969 51872 3980 51901
rect 4048 51872 4077 51901
rect 4077 51872 4104 51901
rect 4172 51872 4185 51901
rect 4185 51872 4228 51901
rect 4296 51872 4349 51901
rect 4349 51872 4352 51901
rect 4420 51872 4457 51901
rect 4457 51872 4476 51901
rect 4544 51872 4565 51901
rect 4565 51872 4600 51901
rect 4668 51872 4673 51901
rect 4673 51872 4724 51901
rect 2808 51748 2864 51804
rect 2932 51748 2988 51804
rect 3056 51748 3112 51804
rect 3180 51748 3236 51804
rect 3304 51748 3360 51804
rect 3428 51748 3484 51804
rect 3552 51748 3608 51804
rect 3676 51748 3732 51804
rect 3800 51748 3856 51804
rect 3924 51748 3980 51804
rect 4048 51748 4104 51804
rect 4172 51748 4228 51804
rect 4296 51748 4352 51804
rect 4420 51748 4476 51804
rect 4544 51748 4600 51804
rect 4668 51748 4724 51804
rect 2808 51624 2864 51680
rect 2932 51624 2988 51680
rect 3056 51624 3112 51680
rect 3180 51624 3236 51680
rect 3304 51624 3360 51680
rect 3428 51624 3484 51680
rect 3552 51624 3608 51680
rect 3676 51624 3732 51680
rect 3800 51624 3856 51680
rect 3924 51624 3980 51680
rect 4048 51624 4104 51680
rect 4172 51624 4228 51680
rect 4296 51624 4352 51680
rect 4420 51624 4476 51680
rect 4544 51624 4600 51680
rect 4668 51624 4724 51680
rect 2808 51500 2864 51556
rect 2932 51500 2988 51556
rect 3056 51500 3112 51556
rect 3180 51500 3236 51556
rect 3304 51500 3360 51556
rect 3428 51500 3484 51556
rect 3552 51500 3608 51556
rect 3676 51500 3732 51556
rect 3800 51500 3856 51556
rect 3924 51500 3980 51556
rect 4048 51500 4104 51556
rect 4172 51500 4228 51556
rect 4296 51500 4352 51556
rect 4420 51500 4476 51556
rect 4544 51500 4600 51556
rect 4668 51500 4724 51556
rect 2808 51376 2864 51432
rect 2932 51376 2988 51432
rect 3056 51376 3112 51432
rect 3180 51376 3236 51432
rect 3304 51376 3360 51432
rect 3428 51376 3484 51432
rect 3552 51376 3608 51432
rect 3676 51376 3732 51432
rect 3800 51376 3856 51432
rect 3924 51376 3980 51432
rect 4048 51376 4104 51432
rect 4172 51376 4228 51432
rect 4296 51376 4352 51432
rect 4420 51376 4476 51432
rect 4544 51376 4600 51432
rect 4668 51376 4724 51432
rect 2808 51252 2864 51308
rect 2932 51252 2988 51308
rect 3056 51252 3112 51308
rect 3180 51252 3236 51308
rect 3304 51252 3360 51308
rect 3428 51252 3484 51308
rect 3552 51252 3608 51308
rect 3676 51252 3732 51308
rect 3800 51252 3856 51308
rect 3924 51252 3980 51308
rect 4048 51252 4104 51308
rect 4172 51252 4228 51308
rect 4296 51252 4352 51308
rect 4420 51252 4476 51308
rect 4544 51252 4600 51308
rect 4668 51252 4724 51308
rect 4861 50892 4917 50948
rect 4985 50892 5041 50948
rect 4861 50768 4917 50824
rect 4985 50768 5041 50824
rect 4861 50685 4917 50700
rect 4985 50685 5041 50700
rect 4861 50644 4871 50685
rect 4871 50644 4917 50685
rect 4985 50644 5031 50685
rect 5031 50644 5041 50685
rect 4861 50525 4871 50576
rect 4871 50525 4917 50576
rect 4985 50525 5031 50576
rect 5031 50525 5041 50576
rect 4861 50520 4917 50525
rect 4985 50520 5041 50525
rect 4861 50396 4917 50452
rect 4985 50396 5041 50452
rect 4861 50272 4917 50328
rect 4985 50272 5041 50328
rect 4861 50148 4917 50204
rect 4985 50148 5041 50204
rect 4861 50024 4917 50080
rect 4985 50024 5041 50080
rect 4861 49900 4917 49956
rect 4985 49900 5041 49956
rect 4861 49776 4917 49832
rect 4985 49776 5041 49832
rect 4861 49699 4871 49708
rect 4871 49699 4917 49708
rect 4985 49699 5031 49708
rect 5031 49699 5041 49708
rect 4861 49652 4917 49699
rect 4985 49652 5041 49699
rect 5178 52492 5234 52548
rect 5302 52492 5358 52548
rect 5426 52492 5482 52548
rect 5550 52492 5606 52548
rect 5674 52492 5730 52548
rect 5798 52492 5854 52548
rect 5922 52492 5978 52548
rect 6046 52492 6102 52548
rect 6170 52492 6226 52548
rect 6294 52492 6350 52548
rect 6418 52492 6474 52548
rect 6542 52492 6598 52548
rect 6666 52492 6722 52548
rect 6790 52492 6846 52548
rect 6914 52492 6970 52548
rect 7038 52492 7094 52548
rect 5178 52368 5234 52424
rect 5302 52368 5358 52424
rect 5426 52368 5482 52424
rect 5550 52368 5606 52424
rect 5674 52368 5730 52424
rect 5798 52368 5854 52424
rect 5922 52368 5978 52424
rect 6046 52368 6102 52424
rect 6170 52368 6226 52424
rect 6294 52368 6350 52424
rect 6418 52368 6474 52424
rect 6542 52368 6598 52424
rect 6666 52368 6722 52424
rect 6790 52368 6846 52424
rect 6914 52368 6970 52424
rect 7038 52368 7094 52424
rect 5178 52244 5234 52300
rect 5302 52244 5358 52300
rect 5426 52244 5482 52300
rect 5550 52244 5606 52300
rect 5674 52244 5730 52300
rect 5798 52244 5854 52300
rect 5922 52244 5978 52300
rect 6046 52244 6102 52300
rect 6170 52244 6226 52300
rect 6294 52244 6350 52300
rect 6418 52244 6474 52300
rect 6542 52244 6598 52300
rect 6666 52244 6722 52300
rect 6790 52244 6846 52300
rect 6914 52244 6970 52300
rect 7038 52244 7094 52300
rect 5178 52120 5234 52176
rect 5302 52120 5358 52176
rect 5426 52120 5482 52176
rect 5550 52120 5606 52176
rect 5674 52120 5730 52176
rect 5798 52120 5854 52176
rect 5922 52120 5978 52176
rect 6046 52120 6102 52176
rect 6170 52120 6226 52176
rect 6294 52120 6350 52176
rect 6418 52120 6474 52176
rect 6542 52120 6598 52176
rect 6666 52120 6722 52176
rect 6790 52120 6846 52176
rect 6914 52120 6970 52176
rect 7038 52120 7094 52176
rect 5178 52009 5234 52052
rect 5302 52009 5358 52052
rect 5426 52009 5482 52052
rect 5550 52009 5606 52052
rect 5674 52009 5730 52052
rect 5798 52009 5854 52052
rect 5922 52009 5978 52052
rect 6046 52009 6102 52052
rect 6170 52009 6226 52052
rect 6294 52009 6350 52052
rect 6418 52009 6474 52052
rect 6542 52009 6598 52052
rect 6666 52009 6722 52052
rect 6790 52009 6846 52052
rect 6914 52009 6970 52052
rect 7038 52009 7094 52052
rect 5178 51996 5190 52009
rect 5190 51996 5234 52009
rect 5302 51996 5354 52009
rect 5354 51996 5358 52009
rect 5426 51996 5462 52009
rect 5462 51996 5482 52009
rect 5550 51996 5570 52009
rect 5570 51996 5606 52009
rect 5674 51996 5678 52009
rect 5678 51996 5730 52009
rect 5798 51996 5838 52009
rect 5838 51996 5854 52009
rect 5922 51996 5946 52009
rect 5946 51996 5978 52009
rect 6046 51996 6054 52009
rect 6054 51996 6102 52009
rect 6170 51996 6218 52009
rect 6218 51996 6226 52009
rect 6294 51996 6326 52009
rect 6326 51996 6350 52009
rect 6418 51996 6434 52009
rect 6434 51996 6474 52009
rect 6542 51996 6594 52009
rect 6594 51996 6598 52009
rect 6666 51996 6702 52009
rect 6702 51996 6722 52009
rect 6790 51996 6810 52009
rect 6810 51996 6846 52009
rect 6914 51996 6918 52009
rect 6918 51996 6970 52009
rect 7038 51996 7082 52009
rect 7082 51996 7094 52009
rect 5178 51901 5234 51928
rect 5302 51901 5358 51928
rect 5426 51901 5482 51928
rect 5550 51901 5606 51928
rect 5674 51901 5730 51928
rect 5798 51901 5854 51928
rect 5922 51901 5978 51928
rect 6046 51901 6102 51928
rect 6170 51901 6226 51928
rect 6294 51901 6350 51928
rect 6418 51901 6474 51928
rect 6542 51901 6598 51928
rect 6666 51901 6722 51928
rect 6790 51901 6846 51928
rect 6914 51901 6970 51928
rect 7038 51901 7094 51928
rect 5178 51872 5190 51901
rect 5190 51872 5234 51901
rect 5302 51872 5354 51901
rect 5354 51872 5358 51901
rect 5426 51872 5462 51901
rect 5462 51872 5482 51901
rect 5550 51872 5570 51901
rect 5570 51872 5606 51901
rect 5674 51872 5678 51901
rect 5678 51872 5730 51901
rect 5798 51872 5838 51901
rect 5838 51872 5854 51901
rect 5922 51872 5946 51901
rect 5946 51872 5978 51901
rect 6046 51872 6054 51901
rect 6054 51872 6102 51901
rect 6170 51872 6218 51901
rect 6218 51872 6226 51901
rect 6294 51872 6326 51901
rect 6326 51872 6350 51901
rect 6418 51872 6434 51901
rect 6434 51872 6474 51901
rect 6542 51872 6594 51901
rect 6594 51872 6598 51901
rect 6666 51872 6702 51901
rect 6702 51872 6722 51901
rect 6790 51872 6810 51901
rect 6810 51872 6846 51901
rect 6914 51872 6918 51901
rect 6918 51872 6970 51901
rect 7038 51872 7082 51901
rect 7082 51872 7094 51901
rect 5178 51748 5234 51804
rect 5302 51748 5358 51804
rect 5426 51748 5482 51804
rect 5550 51748 5606 51804
rect 5674 51748 5730 51804
rect 5798 51748 5854 51804
rect 5922 51748 5978 51804
rect 6046 51748 6102 51804
rect 6170 51748 6226 51804
rect 6294 51748 6350 51804
rect 6418 51748 6474 51804
rect 6542 51748 6598 51804
rect 6666 51748 6722 51804
rect 6790 51748 6846 51804
rect 6914 51748 6970 51804
rect 7038 51748 7094 51804
rect 5178 51624 5234 51680
rect 5302 51624 5358 51680
rect 5426 51624 5482 51680
rect 5550 51624 5606 51680
rect 5674 51624 5730 51680
rect 5798 51624 5854 51680
rect 5922 51624 5978 51680
rect 6046 51624 6102 51680
rect 6170 51624 6226 51680
rect 6294 51624 6350 51680
rect 6418 51624 6474 51680
rect 6542 51624 6598 51680
rect 6666 51624 6722 51680
rect 6790 51624 6846 51680
rect 6914 51624 6970 51680
rect 7038 51624 7094 51680
rect 5178 51500 5234 51556
rect 5302 51500 5358 51556
rect 5426 51500 5482 51556
rect 5550 51500 5606 51556
rect 5674 51500 5730 51556
rect 5798 51500 5854 51556
rect 5922 51500 5978 51556
rect 6046 51500 6102 51556
rect 6170 51500 6226 51556
rect 6294 51500 6350 51556
rect 6418 51500 6474 51556
rect 6542 51500 6598 51556
rect 6666 51500 6722 51556
rect 6790 51500 6846 51556
rect 6914 51500 6970 51556
rect 7038 51500 7094 51556
rect 5178 51376 5234 51432
rect 5302 51376 5358 51432
rect 5426 51376 5482 51432
rect 5550 51376 5606 51432
rect 5674 51376 5730 51432
rect 5798 51376 5854 51432
rect 5922 51376 5978 51432
rect 6046 51376 6102 51432
rect 6170 51376 6226 51432
rect 6294 51376 6350 51432
rect 6418 51376 6474 51432
rect 6542 51376 6598 51432
rect 6666 51376 6722 51432
rect 6790 51376 6846 51432
rect 6914 51376 6970 51432
rect 7038 51376 7094 51432
rect 5178 51252 5234 51308
rect 5302 51252 5358 51308
rect 5426 51252 5482 51308
rect 5550 51252 5606 51308
rect 5674 51252 5730 51308
rect 5798 51252 5854 51308
rect 5922 51252 5978 51308
rect 6046 51252 6102 51308
rect 6170 51252 6226 51308
rect 6294 51252 6350 51308
rect 6418 51252 6474 51308
rect 6542 51252 6598 51308
rect 6666 51252 6722 51308
rect 6790 51252 6846 51308
rect 6914 51252 6970 51308
rect 7038 51252 7094 51308
rect 7275 50892 7331 50948
rect 7399 50892 7455 50948
rect 7523 50892 7579 50948
rect 7647 50892 7703 50948
rect 7275 50768 7331 50824
rect 7399 50768 7455 50824
rect 7523 50768 7579 50824
rect 7647 50768 7703 50824
rect 7275 50685 7331 50700
rect 7399 50685 7455 50700
rect 7523 50685 7579 50700
rect 7647 50685 7703 50700
rect 7275 50644 7299 50685
rect 7299 50644 7331 50685
rect 7399 50644 7407 50685
rect 7407 50644 7455 50685
rect 7523 50644 7571 50685
rect 7571 50644 7579 50685
rect 7647 50644 7679 50685
rect 7679 50644 7703 50685
rect 7275 50525 7299 50576
rect 7299 50525 7331 50576
rect 7399 50525 7407 50576
rect 7407 50525 7455 50576
rect 7523 50525 7571 50576
rect 7571 50525 7579 50576
rect 7647 50525 7679 50576
rect 7679 50525 7703 50576
rect 7275 50520 7331 50525
rect 7399 50520 7455 50525
rect 7523 50520 7579 50525
rect 7647 50520 7703 50525
rect 7275 50396 7331 50452
rect 7399 50396 7455 50452
rect 7523 50396 7579 50452
rect 7647 50396 7703 50452
rect 7275 50272 7331 50328
rect 7399 50272 7455 50328
rect 7523 50272 7579 50328
rect 7647 50272 7703 50328
rect 7275 50148 7331 50204
rect 7399 50148 7455 50204
rect 7523 50148 7579 50204
rect 7647 50148 7703 50204
rect 7275 50024 7331 50080
rect 7399 50024 7455 50080
rect 7523 50024 7579 50080
rect 7647 50024 7703 50080
rect 7275 49900 7331 49956
rect 7399 49900 7455 49956
rect 7523 49900 7579 49956
rect 7647 49900 7703 49956
rect 7275 49776 7331 49832
rect 7399 49776 7455 49832
rect 7523 49776 7579 49832
rect 7647 49776 7703 49832
rect 7275 49699 7299 49708
rect 7299 49699 7331 49708
rect 7399 49699 7407 49708
rect 7407 49699 7455 49708
rect 7523 49699 7571 49708
rect 7571 49699 7579 49708
rect 7647 49699 7679 49708
rect 7679 49699 7703 49708
rect 7275 49652 7331 49699
rect 7399 49652 7455 49699
rect 7523 49652 7579 49699
rect 7647 49652 7703 49699
rect 7884 52492 7940 52548
rect 8008 52492 8064 52548
rect 8132 52492 8188 52548
rect 8256 52492 8312 52548
rect 8380 52492 8436 52548
rect 8504 52492 8560 52548
rect 8628 52492 8684 52548
rect 8752 52492 8808 52548
rect 8876 52492 8932 52548
rect 9000 52492 9056 52548
rect 9124 52492 9180 52548
rect 9248 52492 9304 52548
rect 9372 52492 9428 52548
rect 9496 52492 9552 52548
rect 9620 52492 9676 52548
rect 9744 52492 9800 52548
rect 7884 52368 7940 52424
rect 8008 52368 8064 52424
rect 8132 52368 8188 52424
rect 8256 52368 8312 52424
rect 8380 52368 8436 52424
rect 8504 52368 8560 52424
rect 8628 52368 8684 52424
rect 8752 52368 8808 52424
rect 8876 52368 8932 52424
rect 9000 52368 9056 52424
rect 9124 52368 9180 52424
rect 9248 52368 9304 52424
rect 9372 52368 9428 52424
rect 9496 52368 9552 52424
rect 9620 52368 9676 52424
rect 9744 52368 9800 52424
rect 7884 52244 7940 52300
rect 8008 52244 8064 52300
rect 8132 52244 8188 52300
rect 8256 52244 8312 52300
rect 8380 52244 8436 52300
rect 8504 52244 8560 52300
rect 8628 52244 8684 52300
rect 8752 52244 8808 52300
rect 8876 52244 8932 52300
rect 9000 52244 9056 52300
rect 9124 52244 9180 52300
rect 9248 52244 9304 52300
rect 9372 52244 9428 52300
rect 9496 52244 9552 52300
rect 9620 52244 9676 52300
rect 9744 52244 9800 52300
rect 7884 52120 7940 52176
rect 8008 52120 8064 52176
rect 8132 52120 8188 52176
rect 8256 52120 8312 52176
rect 8380 52120 8436 52176
rect 8504 52120 8560 52176
rect 8628 52120 8684 52176
rect 8752 52120 8808 52176
rect 8876 52120 8932 52176
rect 9000 52120 9056 52176
rect 9124 52120 9180 52176
rect 9248 52120 9304 52176
rect 9372 52120 9428 52176
rect 9496 52120 9552 52176
rect 9620 52120 9676 52176
rect 9744 52120 9800 52176
rect 7884 52009 7940 52052
rect 8008 52009 8064 52052
rect 8132 52009 8188 52052
rect 8256 52009 8312 52052
rect 8380 52009 8436 52052
rect 8504 52009 8560 52052
rect 8628 52009 8684 52052
rect 8752 52009 8808 52052
rect 8876 52009 8932 52052
rect 9000 52009 9056 52052
rect 9124 52009 9180 52052
rect 9248 52009 9304 52052
rect 9372 52009 9428 52052
rect 9496 52009 9552 52052
rect 9620 52009 9676 52052
rect 9744 52009 9800 52052
rect 7884 51996 7896 52009
rect 7896 51996 7940 52009
rect 8008 51996 8060 52009
rect 8060 51996 8064 52009
rect 8132 51996 8168 52009
rect 8168 51996 8188 52009
rect 8256 51996 8276 52009
rect 8276 51996 8312 52009
rect 8380 51996 8384 52009
rect 8384 51996 8436 52009
rect 8504 51996 8544 52009
rect 8544 51996 8560 52009
rect 8628 51996 8652 52009
rect 8652 51996 8684 52009
rect 8752 51996 8760 52009
rect 8760 51996 8808 52009
rect 8876 51996 8924 52009
rect 8924 51996 8932 52009
rect 9000 51996 9032 52009
rect 9032 51996 9056 52009
rect 9124 51996 9140 52009
rect 9140 51996 9180 52009
rect 9248 51996 9300 52009
rect 9300 51996 9304 52009
rect 9372 51996 9408 52009
rect 9408 51996 9428 52009
rect 9496 51996 9516 52009
rect 9516 51996 9552 52009
rect 9620 51996 9624 52009
rect 9624 51996 9676 52009
rect 9744 51996 9788 52009
rect 9788 51996 9800 52009
rect 7884 51901 7940 51928
rect 8008 51901 8064 51928
rect 8132 51901 8188 51928
rect 8256 51901 8312 51928
rect 8380 51901 8436 51928
rect 8504 51901 8560 51928
rect 8628 51901 8684 51928
rect 8752 51901 8808 51928
rect 8876 51901 8932 51928
rect 9000 51901 9056 51928
rect 9124 51901 9180 51928
rect 9248 51901 9304 51928
rect 9372 51901 9428 51928
rect 9496 51901 9552 51928
rect 9620 51901 9676 51928
rect 9744 51901 9800 51928
rect 7884 51872 7896 51901
rect 7896 51872 7940 51901
rect 8008 51872 8060 51901
rect 8060 51872 8064 51901
rect 8132 51872 8168 51901
rect 8168 51872 8188 51901
rect 8256 51872 8276 51901
rect 8276 51872 8312 51901
rect 8380 51872 8384 51901
rect 8384 51872 8436 51901
rect 8504 51872 8544 51901
rect 8544 51872 8560 51901
rect 8628 51872 8652 51901
rect 8652 51872 8684 51901
rect 8752 51872 8760 51901
rect 8760 51872 8808 51901
rect 8876 51872 8924 51901
rect 8924 51872 8932 51901
rect 9000 51872 9032 51901
rect 9032 51872 9056 51901
rect 9124 51872 9140 51901
rect 9140 51872 9180 51901
rect 9248 51872 9300 51901
rect 9300 51872 9304 51901
rect 9372 51872 9408 51901
rect 9408 51872 9428 51901
rect 9496 51872 9516 51901
rect 9516 51872 9552 51901
rect 9620 51872 9624 51901
rect 9624 51872 9676 51901
rect 9744 51872 9788 51901
rect 9788 51872 9800 51901
rect 7884 51748 7940 51804
rect 8008 51748 8064 51804
rect 8132 51748 8188 51804
rect 8256 51748 8312 51804
rect 8380 51748 8436 51804
rect 8504 51748 8560 51804
rect 8628 51748 8684 51804
rect 8752 51748 8808 51804
rect 8876 51748 8932 51804
rect 9000 51748 9056 51804
rect 9124 51748 9180 51804
rect 9248 51748 9304 51804
rect 9372 51748 9428 51804
rect 9496 51748 9552 51804
rect 9620 51748 9676 51804
rect 9744 51748 9800 51804
rect 7884 51624 7940 51680
rect 8008 51624 8064 51680
rect 8132 51624 8188 51680
rect 8256 51624 8312 51680
rect 8380 51624 8436 51680
rect 8504 51624 8560 51680
rect 8628 51624 8684 51680
rect 8752 51624 8808 51680
rect 8876 51624 8932 51680
rect 9000 51624 9056 51680
rect 9124 51624 9180 51680
rect 9248 51624 9304 51680
rect 9372 51624 9428 51680
rect 9496 51624 9552 51680
rect 9620 51624 9676 51680
rect 9744 51624 9800 51680
rect 7884 51500 7940 51556
rect 8008 51500 8064 51556
rect 8132 51500 8188 51556
rect 8256 51500 8312 51556
rect 8380 51500 8436 51556
rect 8504 51500 8560 51556
rect 8628 51500 8684 51556
rect 8752 51500 8808 51556
rect 8876 51500 8932 51556
rect 9000 51500 9056 51556
rect 9124 51500 9180 51556
rect 9248 51500 9304 51556
rect 9372 51500 9428 51556
rect 9496 51500 9552 51556
rect 9620 51500 9676 51556
rect 9744 51500 9800 51556
rect 7884 51376 7940 51432
rect 8008 51376 8064 51432
rect 8132 51376 8188 51432
rect 8256 51376 8312 51432
rect 8380 51376 8436 51432
rect 8504 51376 8560 51432
rect 8628 51376 8684 51432
rect 8752 51376 8808 51432
rect 8876 51376 8932 51432
rect 9000 51376 9056 51432
rect 9124 51376 9180 51432
rect 9248 51376 9304 51432
rect 9372 51376 9428 51432
rect 9496 51376 9552 51432
rect 9620 51376 9676 51432
rect 9744 51376 9800 51432
rect 7884 51252 7940 51308
rect 8008 51252 8064 51308
rect 8132 51252 8188 51308
rect 8256 51252 8312 51308
rect 8380 51252 8436 51308
rect 8504 51252 8560 51308
rect 8628 51252 8684 51308
rect 8752 51252 8808 51308
rect 8876 51252 8932 51308
rect 9000 51252 9056 51308
rect 9124 51252 9180 51308
rect 9248 51252 9304 51308
rect 9372 51252 9428 51308
rect 9496 51252 9552 51308
rect 9620 51252 9676 51308
rect 9744 51252 9800 51308
rect 9937 50892 9993 50948
rect 10061 50892 10117 50948
rect 9937 50768 9993 50824
rect 10061 50768 10117 50824
rect 9937 50685 9993 50700
rect 10061 50685 10117 50700
rect 9937 50644 9947 50685
rect 9947 50644 9993 50685
rect 10061 50644 10107 50685
rect 10107 50644 10117 50685
rect 9937 50525 9947 50576
rect 9947 50525 9993 50576
rect 10061 50525 10107 50576
rect 10107 50525 10117 50576
rect 9937 50520 9993 50525
rect 10061 50520 10117 50525
rect 9937 50396 9993 50452
rect 10061 50396 10117 50452
rect 9937 50272 9993 50328
rect 10061 50272 10117 50328
rect 9937 50148 9993 50204
rect 10061 50148 10117 50204
rect 9937 50024 9993 50080
rect 10061 50024 10117 50080
rect 9937 49900 9993 49956
rect 10061 49900 10117 49956
rect 9937 49776 9993 49832
rect 10061 49776 10117 49832
rect 9937 49699 9947 49708
rect 9947 49699 9993 49708
rect 10061 49699 10107 49708
rect 10107 49699 10117 49708
rect 9937 49652 9993 49699
rect 10061 49652 10117 49699
rect 10254 52492 10310 52548
rect 10378 52492 10434 52548
rect 10502 52492 10558 52548
rect 10626 52492 10682 52548
rect 10750 52492 10806 52548
rect 10874 52492 10930 52548
rect 10998 52492 11054 52548
rect 11122 52492 11178 52548
rect 11246 52492 11302 52548
rect 11370 52492 11426 52548
rect 11494 52492 11550 52548
rect 11618 52492 11674 52548
rect 11742 52492 11798 52548
rect 11866 52492 11922 52548
rect 11990 52492 12046 52548
rect 12114 52492 12170 52548
rect 10254 52368 10310 52424
rect 10378 52368 10434 52424
rect 10502 52368 10558 52424
rect 10626 52368 10682 52424
rect 10750 52368 10806 52424
rect 10874 52368 10930 52424
rect 10998 52368 11054 52424
rect 11122 52368 11178 52424
rect 11246 52368 11302 52424
rect 11370 52368 11426 52424
rect 11494 52368 11550 52424
rect 11618 52368 11674 52424
rect 11742 52368 11798 52424
rect 11866 52368 11922 52424
rect 11990 52368 12046 52424
rect 12114 52368 12170 52424
rect 10254 52244 10310 52300
rect 10378 52244 10434 52300
rect 10502 52244 10558 52300
rect 10626 52244 10682 52300
rect 10750 52244 10806 52300
rect 10874 52244 10930 52300
rect 10998 52244 11054 52300
rect 11122 52244 11178 52300
rect 11246 52244 11302 52300
rect 11370 52244 11426 52300
rect 11494 52244 11550 52300
rect 11618 52244 11674 52300
rect 11742 52244 11798 52300
rect 11866 52244 11922 52300
rect 11990 52244 12046 52300
rect 12114 52244 12170 52300
rect 10254 52120 10310 52176
rect 10378 52120 10434 52176
rect 10502 52120 10558 52176
rect 10626 52120 10682 52176
rect 10750 52120 10806 52176
rect 10874 52120 10930 52176
rect 10998 52120 11054 52176
rect 11122 52120 11178 52176
rect 11246 52120 11302 52176
rect 11370 52120 11426 52176
rect 11494 52120 11550 52176
rect 11618 52120 11674 52176
rect 11742 52120 11798 52176
rect 11866 52120 11922 52176
rect 11990 52120 12046 52176
rect 12114 52120 12170 52176
rect 10254 52009 10310 52052
rect 10378 52009 10434 52052
rect 10502 52009 10558 52052
rect 10626 52009 10682 52052
rect 10750 52009 10806 52052
rect 10874 52009 10930 52052
rect 10998 52009 11054 52052
rect 11122 52009 11178 52052
rect 11246 52009 11302 52052
rect 11370 52009 11426 52052
rect 11494 52009 11550 52052
rect 11618 52009 11674 52052
rect 11742 52009 11798 52052
rect 10254 51996 10305 52009
rect 10305 51996 10310 52009
rect 10378 51996 10413 52009
rect 10413 51996 10434 52009
rect 10502 51996 10521 52009
rect 10521 51996 10558 52009
rect 10626 51996 10629 52009
rect 10629 51996 10682 52009
rect 10750 51996 10793 52009
rect 10793 51996 10806 52009
rect 10874 51996 10901 52009
rect 10901 51996 10930 52009
rect 10998 51996 11009 52009
rect 11009 51996 11054 52009
rect 11122 51996 11169 52009
rect 11169 51996 11178 52009
rect 11246 51996 11277 52009
rect 11277 51996 11302 52009
rect 11370 51996 11385 52009
rect 11385 51996 11426 52009
rect 11494 51996 11549 52009
rect 11549 51996 11550 52009
rect 11618 51996 11657 52009
rect 11657 51996 11674 52009
rect 11742 51996 11765 52009
rect 11765 51996 11798 52009
rect 11866 51996 11922 52052
rect 11990 51996 12046 52052
rect 12114 51996 12170 52052
rect 10254 51901 10310 51928
rect 10378 51901 10434 51928
rect 10502 51901 10558 51928
rect 10626 51901 10682 51928
rect 10750 51901 10806 51928
rect 10874 51901 10930 51928
rect 10998 51901 11054 51928
rect 11122 51901 11178 51928
rect 11246 51901 11302 51928
rect 11370 51901 11426 51928
rect 11494 51901 11550 51928
rect 11618 51901 11674 51928
rect 11742 51901 11798 51928
rect 10254 51872 10305 51901
rect 10305 51872 10310 51901
rect 10378 51872 10413 51901
rect 10413 51872 10434 51901
rect 10502 51872 10521 51901
rect 10521 51872 10558 51901
rect 10626 51872 10629 51901
rect 10629 51872 10682 51901
rect 10750 51872 10793 51901
rect 10793 51872 10806 51901
rect 10874 51872 10901 51901
rect 10901 51872 10930 51901
rect 10998 51872 11009 51901
rect 11009 51872 11054 51901
rect 11122 51872 11169 51901
rect 11169 51872 11178 51901
rect 11246 51872 11277 51901
rect 11277 51872 11302 51901
rect 11370 51872 11385 51901
rect 11385 51872 11426 51901
rect 11494 51872 11549 51901
rect 11549 51872 11550 51901
rect 11618 51872 11657 51901
rect 11657 51872 11674 51901
rect 11742 51872 11765 51901
rect 11765 51872 11798 51901
rect 11866 51872 11922 51928
rect 11990 51872 12046 51928
rect 12114 51872 12170 51928
rect 10254 51748 10310 51804
rect 10378 51748 10434 51804
rect 10502 51748 10558 51804
rect 10626 51748 10682 51804
rect 10750 51748 10806 51804
rect 10874 51748 10930 51804
rect 10998 51748 11054 51804
rect 11122 51748 11178 51804
rect 11246 51748 11302 51804
rect 11370 51748 11426 51804
rect 11494 51748 11550 51804
rect 11618 51748 11674 51804
rect 11742 51748 11798 51804
rect 11866 51748 11922 51804
rect 11990 51748 12046 51804
rect 12114 51748 12170 51804
rect 10254 51624 10310 51680
rect 10378 51624 10434 51680
rect 10502 51624 10558 51680
rect 10626 51624 10682 51680
rect 10750 51624 10806 51680
rect 10874 51624 10930 51680
rect 10998 51624 11054 51680
rect 11122 51624 11178 51680
rect 11246 51624 11302 51680
rect 11370 51624 11426 51680
rect 11494 51624 11550 51680
rect 11618 51624 11674 51680
rect 11742 51624 11798 51680
rect 11866 51624 11922 51680
rect 11990 51624 12046 51680
rect 12114 51624 12170 51680
rect 10254 51500 10310 51556
rect 10378 51500 10434 51556
rect 10502 51500 10558 51556
rect 10626 51500 10682 51556
rect 10750 51500 10806 51556
rect 10874 51500 10930 51556
rect 10998 51500 11054 51556
rect 11122 51500 11178 51556
rect 11246 51500 11302 51556
rect 11370 51500 11426 51556
rect 11494 51500 11550 51556
rect 11618 51500 11674 51556
rect 11742 51500 11798 51556
rect 11866 51500 11922 51556
rect 11990 51500 12046 51556
rect 12114 51500 12170 51556
rect 10254 51376 10310 51432
rect 10378 51376 10434 51432
rect 10502 51376 10558 51432
rect 10626 51376 10682 51432
rect 10750 51376 10806 51432
rect 10874 51376 10930 51432
rect 10998 51376 11054 51432
rect 11122 51376 11178 51432
rect 11246 51376 11302 51432
rect 11370 51376 11426 51432
rect 11494 51376 11550 51432
rect 11618 51376 11674 51432
rect 11742 51376 11798 51432
rect 11866 51376 11922 51432
rect 11990 51376 12046 51432
rect 12114 51376 12170 51432
rect 10254 51252 10310 51308
rect 10378 51252 10434 51308
rect 10502 51252 10558 51308
rect 10626 51252 10682 51308
rect 10750 51252 10806 51308
rect 10874 51252 10930 51308
rect 10998 51252 11054 51308
rect 11122 51252 11178 51308
rect 11246 51252 11302 51308
rect 11370 51252 11426 51308
rect 11494 51252 11550 51308
rect 11618 51252 11674 51308
rect 11742 51252 11798 51308
rect 11866 51252 11922 51308
rect 11990 51252 12046 51308
rect 12114 51252 12170 51308
rect 12307 50922 12336 50948
rect 12336 50922 12363 50948
rect 12307 50892 12363 50922
rect 12431 50892 12487 50948
rect 12307 50814 12336 50824
rect 12336 50814 12363 50824
rect 12307 50768 12363 50814
rect 12431 50768 12487 50824
rect 12307 50650 12363 50700
rect 12307 50644 12336 50650
rect 12336 50644 12363 50650
rect 12431 50644 12487 50700
rect 12307 50542 12363 50576
rect 12307 50520 12336 50542
rect 12336 50520 12363 50542
rect 12431 50520 12487 50576
rect 12307 50434 12363 50452
rect 12307 50396 12336 50434
rect 12336 50396 12363 50434
rect 12431 50396 12487 50452
rect 12307 50326 12363 50328
rect 12307 50274 12336 50326
rect 12336 50274 12363 50326
rect 12307 50272 12363 50274
rect 12431 50272 12487 50328
rect 12307 50166 12336 50204
rect 12336 50166 12363 50204
rect 12307 50148 12363 50166
rect 12431 50148 12487 50204
rect 12307 50058 12336 50080
rect 12336 50058 12363 50080
rect 12307 50024 12363 50058
rect 12431 50024 12487 50080
rect 12307 49950 12336 49956
rect 12336 49950 12363 49956
rect 12307 49900 12363 49950
rect 12431 49900 12487 49956
rect 12307 49786 12363 49832
rect 12307 49776 12336 49786
rect 12336 49776 12363 49786
rect 12431 49776 12487 49832
rect 12307 49678 12363 49708
rect 12307 49652 12336 49678
rect 12336 49652 12363 49678
rect 12431 49652 12487 49708
rect 12871 52492 12927 52548
rect 12995 52492 13051 52548
rect 13119 52492 13175 52548
rect 13243 52492 13299 52548
rect 13367 52492 13423 52548
rect 13491 52492 13547 52548
rect 13615 52492 13671 52548
rect 13739 52492 13795 52548
rect 13863 52492 13919 52548
rect 13987 52492 14043 52548
rect 14111 52492 14167 52548
rect 14235 52492 14291 52548
rect 14359 52492 14415 52548
rect 14483 52492 14539 52548
rect 14607 52492 14663 52548
rect 12871 52368 12927 52424
rect 12995 52368 13051 52424
rect 13119 52368 13175 52424
rect 13243 52368 13299 52424
rect 13367 52368 13423 52424
rect 13491 52368 13547 52424
rect 13615 52368 13671 52424
rect 13739 52368 13795 52424
rect 13863 52368 13919 52424
rect 13987 52368 14043 52424
rect 14111 52368 14167 52424
rect 14235 52368 14291 52424
rect 14359 52368 14415 52424
rect 14483 52368 14539 52424
rect 14607 52368 14663 52424
rect 12871 52244 12927 52300
rect 12995 52244 13051 52300
rect 13119 52244 13175 52300
rect 13243 52244 13299 52300
rect 13367 52244 13423 52300
rect 13491 52244 13547 52300
rect 13615 52244 13671 52300
rect 13739 52244 13795 52300
rect 13863 52244 13919 52300
rect 13987 52244 14043 52300
rect 14111 52244 14167 52300
rect 14235 52244 14291 52300
rect 14359 52244 14415 52300
rect 14483 52244 14539 52300
rect 14607 52244 14663 52300
rect 12871 52120 12927 52176
rect 12995 52120 13051 52176
rect 13119 52120 13175 52176
rect 13243 52120 13299 52176
rect 13367 52120 13423 52176
rect 13491 52120 13547 52176
rect 13615 52120 13671 52176
rect 13739 52120 13795 52176
rect 13863 52120 13919 52176
rect 13987 52120 14043 52176
rect 14111 52120 14167 52176
rect 14235 52120 14291 52176
rect 14359 52120 14415 52176
rect 14483 52120 14539 52176
rect 14607 52120 14663 52176
rect 12871 51996 12927 52052
rect 12995 51996 13051 52052
rect 13119 51996 13175 52052
rect 13243 51996 13299 52052
rect 13367 51996 13423 52052
rect 13491 51996 13547 52052
rect 13615 51996 13671 52052
rect 13739 51996 13795 52052
rect 13863 51996 13919 52052
rect 13987 51996 14043 52052
rect 14111 51996 14167 52052
rect 14235 51996 14291 52052
rect 14359 51996 14415 52052
rect 14483 51996 14539 52052
rect 14607 51996 14663 52052
rect 12871 51872 12927 51928
rect 12995 51872 13051 51928
rect 13119 51872 13175 51928
rect 13243 51872 13299 51928
rect 13367 51872 13423 51928
rect 13491 51872 13547 51928
rect 13615 51872 13671 51928
rect 13739 51872 13795 51928
rect 13863 51872 13919 51928
rect 13987 51872 14043 51928
rect 14111 51872 14167 51928
rect 14235 51872 14291 51928
rect 14359 51872 14415 51928
rect 14483 51872 14539 51928
rect 14607 51872 14663 51928
rect 12871 51748 12927 51804
rect 12995 51748 13051 51804
rect 13119 51748 13175 51804
rect 13243 51748 13299 51804
rect 13367 51748 13423 51804
rect 13491 51748 13547 51804
rect 13615 51748 13671 51804
rect 13739 51748 13795 51804
rect 13863 51748 13919 51804
rect 13987 51748 14043 51804
rect 14111 51748 14167 51804
rect 14235 51748 14291 51804
rect 14359 51748 14415 51804
rect 14483 51748 14539 51804
rect 14607 51748 14663 51804
rect 12871 51624 12927 51680
rect 12995 51624 13051 51680
rect 13119 51624 13175 51680
rect 13243 51624 13299 51680
rect 13367 51624 13423 51680
rect 13491 51624 13547 51680
rect 13615 51624 13671 51680
rect 13739 51624 13795 51680
rect 13863 51624 13919 51680
rect 13987 51624 14043 51680
rect 14111 51624 14167 51680
rect 14235 51624 14291 51680
rect 14359 51624 14415 51680
rect 14483 51624 14539 51680
rect 14607 51624 14663 51680
rect 12871 51500 12927 51556
rect 12995 51500 13051 51556
rect 13119 51500 13175 51556
rect 13243 51500 13299 51556
rect 13367 51500 13423 51556
rect 13491 51500 13547 51556
rect 13615 51500 13671 51556
rect 13739 51500 13795 51556
rect 13863 51500 13919 51556
rect 13987 51500 14043 51556
rect 14111 51500 14167 51556
rect 14235 51500 14291 51556
rect 14359 51500 14415 51556
rect 14483 51500 14539 51556
rect 14607 51500 14663 51556
rect 12871 51376 12927 51432
rect 12995 51376 13051 51432
rect 13119 51376 13175 51432
rect 13243 51376 13299 51432
rect 13367 51376 13423 51432
rect 13491 51376 13547 51432
rect 13615 51376 13671 51432
rect 13739 51376 13795 51432
rect 13863 51376 13919 51432
rect 13987 51376 14043 51432
rect 14111 51376 14167 51432
rect 14235 51376 14291 51432
rect 14359 51376 14415 51432
rect 14483 51376 14539 51432
rect 14607 51376 14663 51432
rect 12871 51252 12927 51308
rect 12995 51252 13051 51308
rect 13119 51252 13175 51308
rect 13243 51252 13299 51308
rect 13367 51252 13423 51308
rect 13491 51252 13547 51308
rect 13615 51252 13671 51308
rect 13739 51252 13795 51308
rect 13863 51252 13919 51308
rect 13987 51252 14043 51308
rect 14111 51252 14167 51308
rect 14235 51252 14291 51308
rect 14359 51252 14415 51308
rect 14483 51252 14539 51308
rect 14607 51252 14663 51308
rect 14902 52574 14958 52576
rect 14902 52522 14904 52574
rect 14904 52522 14956 52574
rect 14956 52522 14958 52574
rect 14902 52466 14958 52522
rect 14902 52414 14904 52466
rect 14904 52414 14956 52466
rect 14956 52414 14958 52466
rect 14902 52358 14958 52414
rect 14902 52306 14904 52358
rect 14904 52306 14956 52358
rect 14956 52306 14958 52358
rect 14902 52250 14958 52306
rect 14902 52198 14904 52250
rect 14904 52198 14956 52250
rect 14956 52198 14958 52250
rect 14902 52142 14958 52198
rect 14902 52090 14904 52142
rect 14904 52090 14956 52142
rect 14956 52090 14958 52142
rect 14902 52034 14958 52090
rect 14902 51982 14904 52034
rect 14904 51982 14956 52034
rect 14956 51982 14958 52034
rect 14902 51926 14958 51982
rect 14902 51874 14904 51926
rect 14904 51874 14956 51926
rect 14956 51874 14958 51926
rect 14902 51818 14958 51874
rect 14902 51766 14904 51818
rect 14904 51766 14956 51818
rect 14956 51766 14958 51818
rect 14902 51710 14958 51766
rect 14902 51658 14904 51710
rect 14904 51658 14956 51710
rect 14956 51658 14958 51710
rect 14902 51602 14958 51658
rect 14902 51550 14904 51602
rect 14904 51550 14956 51602
rect 14956 51550 14958 51602
rect 14902 51494 14958 51550
rect 14902 51442 14904 51494
rect 14904 51442 14956 51494
rect 14956 51442 14958 51494
rect 14902 51386 14958 51442
rect 14902 51334 14904 51386
rect 14904 51334 14956 51386
rect 14956 51334 14958 51386
rect 14902 51278 14958 51334
rect 14902 51226 14904 51278
rect 14904 51226 14956 51278
rect 14956 51226 14958 51278
rect 14902 51224 14958 51226
rect 2302 39671 2358 39727
rect 2491 39692 2547 39748
rect 2615 39692 2671 39748
rect 4861 39692 4917 39748
rect 4985 39692 5041 39748
rect 7275 39692 7331 39748
rect 7399 39692 7455 39748
rect 7523 39692 7579 39748
rect 7647 39692 7703 39748
rect 9937 39692 9993 39748
rect 10061 39692 10117 39748
rect 12307 39692 12363 39748
rect 12431 39692 12487 39748
rect 2302 39539 2358 39595
rect 2491 39568 2547 39624
rect 2615 39568 2671 39624
rect 4861 39568 4917 39624
rect 4985 39568 5041 39624
rect 7275 39568 7331 39624
rect 7399 39568 7455 39624
rect 7523 39568 7579 39624
rect 7647 39568 7703 39624
rect 9937 39568 9993 39624
rect 10061 39568 10117 39624
rect 12307 39568 12363 39624
rect 12431 39568 12487 39624
rect 2302 39407 2358 39463
rect 2491 39444 2547 39500
rect 2615 39444 2671 39500
rect 4861 39444 4917 39500
rect 4985 39444 5041 39500
rect 7275 39444 7331 39500
rect 7399 39444 7455 39500
rect 7523 39444 7579 39500
rect 7647 39444 7703 39500
rect 9937 39444 9993 39500
rect 10061 39444 10117 39500
rect 12307 39444 12363 39500
rect 12431 39444 12487 39500
rect 2302 39275 2358 39331
rect 2491 39320 2547 39376
rect 2615 39320 2671 39376
rect 4861 39320 4917 39376
rect 4985 39320 5041 39376
rect 7275 39320 7331 39376
rect 7399 39320 7455 39376
rect 7523 39320 7579 39376
rect 7647 39320 7703 39376
rect 9937 39320 9993 39376
rect 10061 39320 10117 39376
rect 12307 39320 12363 39376
rect 12431 39320 12487 39376
rect 2302 39143 2358 39199
rect 2491 39196 2547 39252
rect 2615 39196 2671 39252
rect 4861 39196 4917 39252
rect 4985 39196 5041 39252
rect 7275 39196 7331 39252
rect 7399 39196 7455 39252
rect 7523 39196 7579 39252
rect 7647 39196 7703 39252
rect 9937 39196 9993 39252
rect 10061 39196 10117 39252
rect 12307 39196 12363 39252
rect 12431 39196 12487 39252
rect 2491 39072 2547 39128
rect 2615 39072 2671 39128
rect 4861 39072 4917 39128
rect 4985 39072 5041 39128
rect 7275 39072 7331 39128
rect 7399 39072 7455 39128
rect 7523 39072 7579 39128
rect 7647 39072 7703 39128
rect 9937 39072 9993 39128
rect 10061 39072 10117 39128
rect 12307 39072 12363 39128
rect 12431 39072 12487 39128
rect 2302 39011 2358 39067
rect 2491 38948 2547 39004
rect 2615 38948 2671 39004
rect 4861 38948 4917 39004
rect 4985 38948 5041 39004
rect 7275 38948 7331 39004
rect 7399 38948 7455 39004
rect 7523 38948 7579 39004
rect 7647 38948 7703 39004
rect 9937 38948 9993 39004
rect 10061 38948 10117 39004
rect 12307 38948 12363 39004
rect 12431 38948 12487 39004
rect 2302 38879 2358 38935
rect 2491 38824 2547 38880
rect 2615 38824 2671 38880
rect 4861 38824 4917 38880
rect 4985 38824 5041 38880
rect 7275 38824 7331 38880
rect 7399 38824 7455 38880
rect 7523 38824 7579 38880
rect 7647 38824 7703 38880
rect 9937 38824 9993 38880
rect 10061 38824 10117 38880
rect 12307 38824 12363 38880
rect 12431 38824 12487 38880
rect 2302 38747 2358 38803
rect 2491 38700 2547 38756
rect 2615 38700 2671 38756
rect 4861 38700 4917 38756
rect 4985 38700 5041 38756
rect 7275 38700 7331 38756
rect 7399 38700 7455 38756
rect 7523 38700 7579 38756
rect 7647 38700 7703 38756
rect 9937 38700 9993 38756
rect 10061 38700 10117 38756
rect 12307 38700 12363 38756
rect 12431 38700 12487 38756
rect 2302 38615 2358 38671
rect 2491 38576 2547 38632
rect 2615 38576 2671 38632
rect 4861 38576 4917 38632
rect 4985 38576 5041 38632
rect 7275 38576 7331 38632
rect 7399 38576 7455 38632
rect 7523 38576 7579 38632
rect 7647 38576 7703 38632
rect 9937 38576 9993 38632
rect 10061 38576 10117 38632
rect 12307 38576 12363 38632
rect 12431 38576 12487 38632
rect 2302 38483 2358 38539
rect 2491 38452 2547 38508
rect 2615 38452 2671 38508
rect 4861 38452 4917 38508
rect 4985 38452 5041 38508
rect 7275 38452 7331 38508
rect 7399 38452 7455 38508
rect 7523 38452 7579 38508
rect 7647 38452 7703 38508
rect 9937 38452 9993 38508
rect 10061 38452 10117 38508
rect 12307 38452 12363 38508
rect 12431 38452 12487 38508
rect 20 38174 76 38176
rect 20 38122 22 38174
rect 22 38122 74 38174
rect 74 38122 76 38174
rect 20 38066 76 38122
rect 20 38014 22 38066
rect 22 38014 74 38066
rect 74 38014 76 38066
rect 20 37958 76 38014
rect 20 37906 22 37958
rect 22 37906 74 37958
rect 74 37906 76 37958
rect 20 37850 76 37906
rect 20 37798 22 37850
rect 22 37798 74 37850
rect 74 37798 76 37850
rect 20 37742 76 37798
rect 20 37690 22 37742
rect 22 37690 74 37742
rect 74 37690 76 37742
rect 20 37634 76 37690
rect 20 37582 22 37634
rect 22 37582 74 37634
rect 74 37582 76 37634
rect 20 37526 76 37582
rect 20 37474 22 37526
rect 22 37474 74 37526
rect 74 37474 76 37526
rect 20 37418 76 37474
rect 20 37366 22 37418
rect 22 37366 74 37418
rect 74 37366 76 37418
rect 20 37310 76 37366
rect 20 37258 22 37310
rect 22 37258 74 37310
rect 74 37258 76 37310
rect 20 37202 76 37258
rect 20 37150 22 37202
rect 22 37150 74 37202
rect 74 37150 76 37202
rect 20 37094 76 37150
rect 20 37042 22 37094
rect 22 37042 74 37094
rect 74 37042 76 37094
rect 20 36986 76 37042
rect 20 36934 22 36986
rect 22 36934 74 36986
rect 74 36934 76 36986
rect 20 36878 76 36934
rect 20 36826 22 36878
rect 22 36826 74 36878
rect 74 36826 76 36878
rect 20 36824 76 36826
rect 315 38092 371 38148
rect 439 38092 495 38148
rect 563 38092 619 38148
rect 687 38092 743 38148
rect 811 38092 867 38148
rect 935 38092 991 38148
rect 1059 38092 1115 38148
rect 1183 38092 1239 38148
rect 1307 38092 1363 38148
rect 1431 38092 1487 38148
rect 1555 38092 1611 38148
rect 1679 38092 1735 38148
rect 1803 38092 1859 38148
rect 1927 38092 1983 38148
rect 2051 38092 2107 38148
rect 2808 38092 2864 38148
rect 2932 38092 2988 38148
rect 3056 38092 3112 38148
rect 3180 38092 3236 38148
rect 3304 38092 3360 38148
rect 3428 38092 3484 38148
rect 3552 38092 3608 38148
rect 3676 38092 3732 38148
rect 3800 38092 3856 38148
rect 3924 38092 3980 38148
rect 4048 38092 4104 38148
rect 4172 38092 4228 38148
rect 4296 38092 4352 38148
rect 4420 38092 4476 38148
rect 4544 38092 4600 38148
rect 4668 38092 4724 38148
rect 5178 38092 5234 38148
rect 5302 38092 5358 38148
rect 5426 38092 5482 38148
rect 5550 38092 5606 38148
rect 5674 38092 5730 38148
rect 5798 38092 5854 38148
rect 5922 38092 5978 38148
rect 6046 38092 6102 38148
rect 6170 38092 6226 38148
rect 6294 38092 6350 38148
rect 6418 38092 6474 38148
rect 6542 38092 6598 38148
rect 6666 38092 6722 38148
rect 6790 38092 6846 38148
rect 6914 38092 6970 38148
rect 7038 38092 7094 38148
rect 7884 38092 7940 38148
rect 8008 38092 8064 38148
rect 8132 38092 8188 38148
rect 8256 38092 8312 38148
rect 8380 38092 8436 38148
rect 8504 38092 8560 38148
rect 8628 38092 8684 38148
rect 8752 38092 8808 38148
rect 8876 38092 8932 38148
rect 9000 38092 9056 38148
rect 9124 38092 9180 38148
rect 9248 38092 9304 38148
rect 9372 38092 9428 38148
rect 9496 38092 9552 38148
rect 9620 38092 9676 38148
rect 9744 38092 9800 38148
rect 10254 38092 10310 38148
rect 10378 38092 10434 38148
rect 10502 38092 10558 38148
rect 10626 38092 10682 38148
rect 10750 38092 10806 38148
rect 10874 38092 10930 38148
rect 10998 38092 11054 38148
rect 11122 38092 11178 38148
rect 11246 38092 11302 38148
rect 11370 38092 11426 38148
rect 11494 38092 11550 38148
rect 11618 38092 11674 38148
rect 11742 38092 11798 38148
rect 11866 38092 11922 38148
rect 11990 38092 12046 38148
rect 12114 38092 12170 38148
rect 12871 38092 12927 38148
rect 12995 38092 13051 38148
rect 13119 38092 13175 38148
rect 13243 38092 13299 38148
rect 13367 38092 13423 38148
rect 13491 38092 13547 38148
rect 13615 38092 13671 38148
rect 13739 38092 13795 38148
rect 13863 38092 13919 38148
rect 13987 38092 14043 38148
rect 14111 38092 14167 38148
rect 14235 38092 14291 38148
rect 14359 38092 14415 38148
rect 14483 38092 14539 38148
rect 14607 38092 14663 38148
rect 315 37968 371 38024
rect 439 37968 495 38024
rect 563 37968 619 38024
rect 687 37968 743 38024
rect 811 37968 867 38024
rect 935 37968 991 38024
rect 1059 37968 1115 38024
rect 1183 37968 1239 38024
rect 1307 37968 1363 38024
rect 1431 37968 1487 38024
rect 1555 37968 1611 38024
rect 1679 37968 1735 38024
rect 1803 37968 1859 38024
rect 1927 37968 1983 38024
rect 2051 37968 2107 38024
rect 2808 37968 2864 38024
rect 2932 37968 2988 38024
rect 3056 37968 3112 38024
rect 3180 37968 3236 38024
rect 3304 37968 3360 38024
rect 3428 37968 3484 38024
rect 3552 37968 3608 38024
rect 3676 37968 3732 38024
rect 3800 37968 3856 38024
rect 3924 37968 3980 38024
rect 4048 37968 4104 38024
rect 4172 37968 4228 38024
rect 4296 37968 4352 38024
rect 4420 37968 4476 38024
rect 4544 37968 4600 38024
rect 4668 37968 4724 38024
rect 5178 37968 5234 38024
rect 5302 37968 5358 38024
rect 5426 37968 5482 38024
rect 5550 37968 5606 38024
rect 5674 37968 5730 38024
rect 5798 37968 5854 38024
rect 5922 37968 5978 38024
rect 6046 37968 6102 38024
rect 6170 37968 6226 38024
rect 6294 37968 6350 38024
rect 6418 37968 6474 38024
rect 6542 37968 6598 38024
rect 6666 37968 6722 38024
rect 6790 37968 6846 38024
rect 6914 37968 6970 38024
rect 7038 37968 7094 38024
rect 7884 37968 7940 38024
rect 8008 37968 8064 38024
rect 8132 37968 8188 38024
rect 8256 37968 8312 38024
rect 8380 37968 8436 38024
rect 8504 37968 8560 38024
rect 8628 37968 8684 38024
rect 8752 37968 8808 38024
rect 8876 37968 8932 38024
rect 9000 37968 9056 38024
rect 9124 37968 9180 38024
rect 9248 37968 9304 38024
rect 9372 37968 9428 38024
rect 9496 37968 9552 38024
rect 9620 37968 9676 38024
rect 9744 37968 9800 38024
rect 10254 37968 10310 38024
rect 10378 37968 10434 38024
rect 10502 37968 10558 38024
rect 10626 37968 10682 38024
rect 10750 37968 10806 38024
rect 10874 37968 10930 38024
rect 10998 37968 11054 38024
rect 11122 37968 11178 38024
rect 11246 37968 11302 38024
rect 11370 37968 11426 38024
rect 11494 37968 11550 38024
rect 11618 37968 11674 38024
rect 11742 37968 11798 38024
rect 11866 37968 11922 38024
rect 11990 37968 12046 38024
rect 12114 37968 12170 38024
rect 12871 37968 12927 38024
rect 12995 37968 13051 38024
rect 13119 37968 13175 38024
rect 13243 37968 13299 38024
rect 13367 37968 13423 38024
rect 13491 37968 13547 38024
rect 13615 37968 13671 38024
rect 13739 37968 13795 38024
rect 13863 37968 13919 38024
rect 13987 37968 14043 38024
rect 14111 37968 14167 38024
rect 14235 37968 14291 38024
rect 14359 37968 14415 38024
rect 14483 37968 14539 38024
rect 14607 37968 14663 38024
rect 315 37844 371 37900
rect 439 37844 495 37900
rect 563 37844 619 37900
rect 687 37844 743 37900
rect 811 37844 867 37900
rect 935 37844 991 37900
rect 1059 37844 1115 37900
rect 1183 37844 1239 37900
rect 1307 37844 1363 37900
rect 1431 37844 1487 37900
rect 1555 37844 1611 37900
rect 1679 37844 1735 37900
rect 1803 37844 1859 37900
rect 1927 37844 1983 37900
rect 2051 37844 2107 37900
rect 2808 37844 2864 37900
rect 2932 37844 2988 37900
rect 3056 37844 3112 37900
rect 3180 37844 3236 37900
rect 3304 37844 3360 37900
rect 3428 37844 3484 37900
rect 3552 37844 3608 37900
rect 3676 37844 3732 37900
rect 3800 37844 3856 37900
rect 3924 37844 3980 37900
rect 4048 37844 4104 37900
rect 4172 37844 4228 37900
rect 4296 37844 4352 37900
rect 4420 37844 4476 37900
rect 4544 37844 4600 37900
rect 4668 37844 4724 37900
rect 5178 37844 5234 37900
rect 5302 37844 5358 37900
rect 5426 37844 5482 37900
rect 5550 37844 5606 37900
rect 5674 37844 5730 37900
rect 5798 37844 5854 37900
rect 5922 37844 5978 37900
rect 6046 37844 6102 37900
rect 6170 37844 6226 37900
rect 6294 37844 6350 37900
rect 6418 37844 6474 37900
rect 6542 37844 6598 37900
rect 6666 37844 6722 37900
rect 6790 37844 6846 37900
rect 6914 37844 6970 37900
rect 7038 37844 7094 37900
rect 7884 37844 7940 37900
rect 8008 37844 8064 37900
rect 8132 37844 8188 37900
rect 8256 37844 8312 37900
rect 8380 37844 8436 37900
rect 8504 37844 8560 37900
rect 8628 37844 8684 37900
rect 8752 37844 8808 37900
rect 8876 37844 8932 37900
rect 9000 37844 9056 37900
rect 9124 37844 9180 37900
rect 9248 37844 9304 37900
rect 9372 37844 9428 37900
rect 9496 37844 9552 37900
rect 9620 37844 9676 37900
rect 9744 37844 9800 37900
rect 10254 37844 10310 37900
rect 10378 37844 10434 37900
rect 10502 37844 10558 37900
rect 10626 37844 10682 37900
rect 10750 37844 10806 37900
rect 10874 37844 10930 37900
rect 10998 37844 11054 37900
rect 11122 37844 11178 37900
rect 11246 37844 11302 37900
rect 11370 37844 11426 37900
rect 11494 37844 11550 37900
rect 11618 37844 11674 37900
rect 11742 37844 11798 37900
rect 11866 37844 11922 37900
rect 11990 37844 12046 37900
rect 12114 37844 12170 37900
rect 12871 37844 12927 37900
rect 12995 37844 13051 37900
rect 13119 37844 13175 37900
rect 13243 37844 13299 37900
rect 13367 37844 13423 37900
rect 13491 37844 13547 37900
rect 13615 37844 13671 37900
rect 13739 37844 13795 37900
rect 13863 37844 13919 37900
rect 13987 37844 14043 37900
rect 14111 37844 14167 37900
rect 14235 37844 14291 37900
rect 14359 37844 14415 37900
rect 14483 37844 14539 37900
rect 14607 37844 14663 37900
rect 315 37720 371 37776
rect 439 37720 495 37776
rect 563 37720 619 37776
rect 687 37720 743 37776
rect 811 37720 867 37776
rect 935 37720 991 37776
rect 1059 37720 1115 37776
rect 1183 37720 1239 37776
rect 1307 37720 1363 37776
rect 1431 37720 1487 37776
rect 1555 37720 1611 37776
rect 1679 37720 1735 37776
rect 1803 37720 1859 37776
rect 1927 37720 1983 37776
rect 2051 37720 2107 37776
rect 2808 37720 2864 37776
rect 2932 37720 2988 37776
rect 3056 37720 3112 37776
rect 3180 37720 3236 37776
rect 3304 37720 3360 37776
rect 3428 37720 3484 37776
rect 3552 37720 3608 37776
rect 3676 37720 3732 37776
rect 3800 37720 3856 37776
rect 3924 37720 3980 37776
rect 4048 37720 4104 37776
rect 4172 37720 4228 37776
rect 4296 37720 4352 37776
rect 4420 37720 4476 37776
rect 4544 37720 4600 37776
rect 4668 37720 4724 37776
rect 5178 37720 5234 37776
rect 5302 37720 5358 37776
rect 5426 37720 5482 37776
rect 5550 37720 5606 37776
rect 5674 37720 5730 37776
rect 5798 37720 5854 37776
rect 5922 37720 5978 37776
rect 6046 37720 6102 37776
rect 6170 37720 6226 37776
rect 6294 37720 6350 37776
rect 6418 37720 6474 37776
rect 6542 37720 6598 37776
rect 6666 37720 6722 37776
rect 6790 37720 6846 37776
rect 6914 37720 6970 37776
rect 7038 37720 7094 37776
rect 7884 37720 7940 37776
rect 8008 37720 8064 37776
rect 8132 37720 8188 37776
rect 8256 37720 8312 37776
rect 8380 37720 8436 37776
rect 8504 37720 8560 37776
rect 8628 37720 8684 37776
rect 8752 37720 8808 37776
rect 8876 37720 8932 37776
rect 9000 37720 9056 37776
rect 9124 37720 9180 37776
rect 9248 37720 9304 37776
rect 9372 37720 9428 37776
rect 9496 37720 9552 37776
rect 9620 37720 9676 37776
rect 9744 37720 9800 37776
rect 10254 37720 10310 37776
rect 10378 37720 10434 37776
rect 10502 37720 10558 37776
rect 10626 37720 10682 37776
rect 10750 37720 10806 37776
rect 10874 37720 10930 37776
rect 10998 37720 11054 37776
rect 11122 37720 11178 37776
rect 11246 37720 11302 37776
rect 11370 37720 11426 37776
rect 11494 37720 11550 37776
rect 11618 37720 11674 37776
rect 11742 37720 11798 37776
rect 11866 37720 11922 37776
rect 11990 37720 12046 37776
rect 12114 37720 12170 37776
rect 12871 37720 12927 37776
rect 12995 37720 13051 37776
rect 13119 37720 13175 37776
rect 13243 37720 13299 37776
rect 13367 37720 13423 37776
rect 13491 37720 13547 37776
rect 13615 37720 13671 37776
rect 13739 37720 13795 37776
rect 13863 37720 13919 37776
rect 13987 37720 14043 37776
rect 14111 37720 14167 37776
rect 14235 37720 14291 37776
rect 14359 37720 14415 37776
rect 14483 37720 14539 37776
rect 14607 37720 14663 37776
rect 315 37596 371 37652
rect 439 37596 495 37652
rect 563 37596 619 37652
rect 687 37596 743 37652
rect 811 37596 867 37652
rect 935 37596 991 37652
rect 1059 37596 1115 37652
rect 1183 37596 1239 37652
rect 1307 37596 1363 37652
rect 1431 37596 1487 37652
rect 1555 37596 1611 37652
rect 1679 37596 1735 37652
rect 1803 37596 1859 37652
rect 1927 37596 1983 37652
rect 2051 37596 2107 37652
rect 2808 37596 2864 37652
rect 2932 37596 2988 37652
rect 3056 37596 3112 37652
rect 3180 37596 3236 37652
rect 3304 37596 3360 37652
rect 3428 37596 3484 37652
rect 3552 37596 3608 37652
rect 3676 37596 3732 37652
rect 3800 37596 3856 37652
rect 3924 37596 3980 37652
rect 4048 37596 4104 37652
rect 4172 37596 4228 37652
rect 4296 37596 4352 37652
rect 4420 37596 4476 37652
rect 4544 37596 4600 37652
rect 4668 37596 4724 37652
rect 5178 37596 5234 37652
rect 5302 37596 5358 37652
rect 5426 37596 5482 37652
rect 5550 37596 5606 37652
rect 5674 37596 5730 37652
rect 5798 37596 5854 37652
rect 5922 37596 5978 37652
rect 6046 37596 6102 37652
rect 6170 37596 6226 37652
rect 6294 37596 6350 37652
rect 6418 37596 6474 37652
rect 6542 37596 6598 37652
rect 6666 37596 6722 37652
rect 6790 37596 6846 37652
rect 6914 37596 6970 37652
rect 7038 37596 7094 37652
rect 7884 37596 7940 37652
rect 8008 37596 8064 37652
rect 8132 37596 8188 37652
rect 8256 37596 8312 37652
rect 8380 37596 8436 37652
rect 8504 37596 8560 37652
rect 8628 37596 8684 37652
rect 8752 37596 8808 37652
rect 8876 37596 8932 37652
rect 9000 37596 9056 37652
rect 9124 37596 9180 37652
rect 9248 37596 9304 37652
rect 9372 37596 9428 37652
rect 9496 37596 9552 37652
rect 9620 37596 9676 37652
rect 9744 37596 9800 37652
rect 10254 37596 10310 37652
rect 10378 37596 10434 37652
rect 10502 37596 10558 37652
rect 10626 37596 10682 37652
rect 10750 37596 10806 37652
rect 10874 37596 10930 37652
rect 10998 37596 11054 37652
rect 11122 37596 11178 37652
rect 11246 37596 11302 37652
rect 11370 37596 11426 37652
rect 11494 37596 11550 37652
rect 11618 37596 11674 37652
rect 11742 37596 11798 37652
rect 11866 37596 11922 37652
rect 11990 37596 12046 37652
rect 12114 37596 12170 37652
rect 12871 37596 12927 37652
rect 12995 37596 13051 37652
rect 13119 37596 13175 37652
rect 13243 37596 13299 37652
rect 13367 37596 13423 37652
rect 13491 37596 13547 37652
rect 13615 37596 13671 37652
rect 13739 37596 13795 37652
rect 13863 37596 13919 37652
rect 13987 37596 14043 37652
rect 14111 37596 14167 37652
rect 14235 37596 14291 37652
rect 14359 37596 14415 37652
rect 14483 37596 14539 37652
rect 14607 37596 14663 37652
rect 315 37472 371 37528
rect 439 37472 495 37528
rect 563 37472 619 37528
rect 687 37472 743 37528
rect 811 37472 867 37528
rect 935 37472 991 37528
rect 1059 37472 1115 37528
rect 1183 37472 1239 37528
rect 1307 37472 1363 37528
rect 1431 37472 1487 37528
rect 1555 37472 1611 37528
rect 1679 37472 1735 37528
rect 1803 37472 1859 37528
rect 1927 37472 1983 37528
rect 2051 37472 2107 37528
rect 2808 37472 2864 37528
rect 2932 37472 2988 37528
rect 3056 37472 3112 37528
rect 3180 37472 3236 37528
rect 3304 37472 3360 37528
rect 3428 37472 3484 37528
rect 3552 37472 3608 37528
rect 3676 37472 3732 37528
rect 3800 37472 3856 37528
rect 3924 37472 3980 37528
rect 4048 37472 4104 37528
rect 4172 37472 4228 37528
rect 4296 37472 4352 37528
rect 4420 37472 4476 37528
rect 4544 37472 4600 37528
rect 4668 37472 4724 37528
rect 5178 37472 5234 37528
rect 5302 37472 5358 37528
rect 5426 37472 5482 37528
rect 5550 37472 5606 37528
rect 5674 37472 5730 37528
rect 5798 37472 5854 37528
rect 5922 37472 5978 37528
rect 6046 37472 6102 37528
rect 6170 37472 6226 37528
rect 6294 37472 6350 37528
rect 6418 37472 6474 37528
rect 6542 37472 6598 37528
rect 6666 37472 6722 37528
rect 6790 37472 6846 37528
rect 6914 37472 6970 37528
rect 7038 37472 7094 37528
rect 7884 37472 7940 37528
rect 8008 37472 8064 37528
rect 8132 37472 8188 37528
rect 8256 37472 8312 37528
rect 8380 37472 8436 37528
rect 8504 37472 8560 37528
rect 8628 37472 8684 37528
rect 8752 37472 8808 37528
rect 8876 37472 8932 37528
rect 9000 37472 9056 37528
rect 9124 37472 9180 37528
rect 9248 37472 9304 37528
rect 9372 37472 9428 37528
rect 9496 37472 9552 37528
rect 9620 37472 9676 37528
rect 9744 37472 9800 37528
rect 10254 37472 10310 37528
rect 10378 37472 10434 37528
rect 10502 37472 10558 37528
rect 10626 37472 10682 37528
rect 10750 37472 10806 37528
rect 10874 37472 10930 37528
rect 10998 37472 11054 37528
rect 11122 37472 11178 37528
rect 11246 37472 11302 37528
rect 11370 37472 11426 37528
rect 11494 37472 11550 37528
rect 11618 37472 11674 37528
rect 11742 37472 11798 37528
rect 11866 37472 11922 37528
rect 11990 37472 12046 37528
rect 12114 37472 12170 37528
rect 12871 37472 12927 37528
rect 12995 37472 13051 37528
rect 13119 37472 13175 37528
rect 13243 37472 13299 37528
rect 13367 37472 13423 37528
rect 13491 37472 13547 37528
rect 13615 37472 13671 37528
rect 13739 37472 13795 37528
rect 13863 37472 13919 37528
rect 13987 37472 14043 37528
rect 14111 37472 14167 37528
rect 14235 37472 14291 37528
rect 14359 37472 14415 37528
rect 14483 37472 14539 37528
rect 14607 37472 14663 37528
rect 315 37348 371 37404
rect 439 37348 495 37404
rect 563 37348 619 37404
rect 687 37348 743 37404
rect 811 37348 867 37404
rect 935 37348 991 37404
rect 1059 37348 1115 37404
rect 1183 37348 1239 37404
rect 1307 37348 1363 37404
rect 1431 37348 1487 37404
rect 1555 37348 1611 37404
rect 1679 37348 1735 37404
rect 1803 37348 1859 37404
rect 1927 37348 1983 37404
rect 2051 37348 2107 37404
rect 2808 37348 2864 37404
rect 2932 37348 2988 37404
rect 3056 37348 3112 37404
rect 3180 37348 3236 37404
rect 3304 37348 3360 37404
rect 3428 37348 3484 37404
rect 3552 37348 3608 37404
rect 3676 37348 3732 37404
rect 3800 37348 3856 37404
rect 3924 37348 3980 37404
rect 4048 37348 4104 37404
rect 4172 37348 4228 37404
rect 4296 37348 4352 37404
rect 4420 37348 4476 37404
rect 4544 37348 4600 37404
rect 4668 37348 4724 37404
rect 5178 37348 5234 37404
rect 5302 37348 5358 37404
rect 5426 37348 5482 37404
rect 5550 37348 5606 37404
rect 5674 37348 5730 37404
rect 5798 37348 5854 37404
rect 5922 37348 5978 37404
rect 6046 37348 6102 37404
rect 6170 37348 6226 37404
rect 6294 37348 6350 37404
rect 6418 37348 6474 37404
rect 6542 37348 6598 37404
rect 6666 37348 6722 37404
rect 6790 37348 6846 37404
rect 6914 37348 6970 37404
rect 7038 37348 7094 37404
rect 7884 37348 7940 37404
rect 8008 37348 8064 37404
rect 8132 37348 8188 37404
rect 8256 37348 8312 37404
rect 8380 37348 8436 37404
rect 8504 37348 8560 37404
rect 8628 37348 8684 37404
rect 8752 37348 8808 37404
rect 8876 37348 8932 37404
rect 9000 37348 9056 37404
rect 9124 37348 9180 37404
rect 9248 37348 9304 37404
rect 9372 37348 9428 37404
rect 9496 37348 9552 37404
rect 9620 37348 9676 37404
rect 9744 37348 9800 37404
rect 10254 37348 10310 37404
rect 10378 37348 10434 37404
rect 10502 37348 10558 37404
rect 10626 37348 10682 37404
rect 10750 37348 10806 37404
rect 10874 37348 10930 37404
rect 10998 37348 11054 37404
rect 11122 37348 11178 37404
rect 11246 37348 11302 37404
rect 11370 37348 11426 37404
rect 11494 37348 11550 37404
rect 11618 37348 11674 37404
rect 11742 37348 11798 37404
rect 11866 37348 11922 37404
rect 11990 37348 12046 37404
rect 12114 37348 12170 37404
rect 12871 37348 12927 37404
rect 12995 37348 13051 37404
rect 13119 37348 13175 37404
rect 13243 37348 13299 37404
rect 13367 37348 13423 37404
rect 13491 37348 13547 37404
rect 13615 37348 13671 37404
rect 13739 37348 13795 37404
rect 13863 37348 13919 37404
rect 13987 37348 14043 37404
rect 14111 37348 14167 37404
rect 14235 37348 14291 37404
rect 14359 37348 14415 37404
rect 14483 37348 14539 37404
rect 14607 37348 14663 37404
rect 315 37224 371 37280
rect 439 37224 495 37280
rect 563 37224 619 37280
rect 687 37224 743 37280
rect 811 37224 867 37280
rect 935 37224 991 37280
rect 1059 37224 1115 37280
rect 1183 37224 1239 37280
rect 1307 37224 1363 37280
rect 1431 37224 1487 37280
rect 1555 37224 1611 37280
rect 1679 37224 1735 37280
rect 1803 37224 1859 37280
rect 1927 37224 1983 37280
rect 2051 37224 2107 37280
rect 2808 37224 2864 37280
rect 2932 37224 2988 37280
rect 3056 37224 3112 37280
rect 3180 37224 3236 37280
rect 3304 37224 3360 37280
rect 3428 37224 3484 37280
rect 3552 37224 3608 37280
rect 3676 37224 3732 37280
rect 3800 37224 3856 37280
rect 3924 37224 3980 37280
rect 4048 37224 4104 37280
rect 4172 37224 4228 37280
rect 4296 37224 4352 37280
rect 4420 37224 4476 37280
rect 4544 37224 4600 37280
rect 4668 37224 4724 37280
rect 5178 37224 5234 37280
rect 5302 37224 5358 37280
rect 5426 37224 5482 37280
rect 5550 37224 5606 37280
rect 5674 37224 5730 37280
rect 5798 37224 5854 37280
rect 5922 37224 5978 37280
rect 6046 37224 6102 37280
rect 6170 37224 6226 37280
rect 6294 37224 6350 37280
rect 6418 37224 6474 37280
rect 6542 37224 6598 37280
rect 6666 37224 6722 37280
rect 6790 37224 6846 37280
rect 6914 37224 6970 37280
rect 7038 37224 7094 37280
rect 7884 37224 7940 37280
rect 8008 37224 8064 37280
rect 8132 37224 8188 37280
rect 8256 37224 8312 37280
rect 8380 37224 8436 37280
rect 8504 37224 8560 37280
rect 8628 37224 8684 37280
rect 8752 37224 8808 37280
rect 8876 37224 8932 37280
rect 9000 37224 9056 37280
rect 9124 37224 9180 37280
rect 9248 37224 9304 37280
rect 9372 37224 9428 37280
rect 9496 37224 9552 37280
rect 9620 37224 9676 37280
rect 9744 37224 9800 37280
rect 10254 37224 10310 37280
rect 10378 37224 10434 37280
rect 10502 37224 10558 37280
rect 10626 37224 10682 37280
rect 10750 37224 10806 37280
rect 10874 37224 10930 37280
rect 10998 37224 11054 37280
rect 11122 37224 11178 37280
rect 11246 37224 11302 37280
rect 11370 37224 11426 37280
rect 11494 37224 11550 37280
rect 11618 37224 11674 37280
rect 11742 37224 11798 37280
rect 11866 37224 11922 37280
rect 11990 37224 12046 37280
rect 12114 37224 12170 37280
rect 12871 37224 12927 37280
rect 12995 37224 13051 37280
rect 13119 37224 13175 37280
rect 13243 37224 13299 37280
rect 13367 37224 13423 37280
rect 13491 37224 13547 37280
rect 13615 37224 13671 37280
rect 13739 37224 13795 37280
rect 13863 37224 13919 37280
rect 13987 37224 14043 37280
rect 14111 37224 14167 37280
rect 14235 37224 14291 37280
rect 14359 37224 14415 37280
rect 14483 37224 14539 37280
rect 14607 37224 14663 37280
rect 315 37100 371 37156
rect 439 37100 495 37156
rect 563 37100 619 37156
rect 687 37100 743 37156
rect 811 37100 867 37156
rect 935 37100 991 37156
rect 1059 37100 1115 37156
rect 1183 37100 1239 37156
rect 1307 37100 1363 37156
rect 1431 37100 1487 37156
rect 1555 37100 1611 37156
rect 1679 37100 1735 37156
rect 1803 37100 1859 37156
rect 1927 37100 1983 37156
rect 2051 37100 2107 37156
rect 2808 37100 2864 37156
rect 2932 37100 2988 37156
rect 3056 37100 3112 37156
rect 3180 37100 3236 37156
rect 3304 37100 3360 37156
rect 3428 37100 3484 37156
rect 3552 37100 3608 37156
rect 3676 37100 3732 37156
rect 3800 37100 3856 37156
rect 3924 37100 3980 37156
rect 4048 37100 4104 37156
rect 4172 37100 4228 37156
rect 4296 37100 4352 37156
rect 4420 37100 4476 37156
rect 4544 37100 4600 37156
rect 4668 37100 4724 37156
rect 5178 37100 5234 37156
rect 5302 37100 5358 37156
rect 5426 37100 5482 37156
rect 5550 37100 5606 37156
rect 5674 37100 5730 37156
rect 5798 37100 5854 37156
rect 5922 37100 5978 37156
rect 6046 37100 6102 37156
rect 6170 37100 6226 37156
rect 6294 37100 6350 37156
rect 6418 37100 6474 37156
rect 6542 37100 6598 37156
rect 6666 37100 6722 37156
rect 6790 37100 6846 37156
rect 6914 37100 6970 37156
rect 7038 37100 7094 37156
rect 7884 37100 7940 37156
rect 8008 37100 8064 37156
rect 8132 37100 8188 37156
rect 8256 37100 8312 37156
rect 8380 37100 8436 37156
rect 8504 37100 8560 37156
rect 8628 37100 8684 37156
rect 8752 37100 8808 37156
rect 8876 37100 8932 37156
rect 9000 37100 9056 37156
rect 9124 37100 9180 37156
rect 9248 37100 9304 37156
rect 9372 37100 9428 37156
rect 9496 37100 9552 37156
rect 9620 37100 9676 37156
rect 9744 37100 9800 37156
rect 10254 37100 10310 37156
rect 10378 37100 10434 37156
rect 10502 37100 10558 37156
rect 10626 37100 10682 37156
rect 10750 37100 10806 37156
rect 10874 37100 10930 37156
rect 10998 37100 11054 37156
rect 11122 37100 11178 37156
rect 11246 37100 11302 37156
rect 11370 37100 11426 37156
rect 11494 37100 11550 37156
rect 11618 37100 11674 37156
rect 11742 37100 11798 37156
rect 11866 37100 11922 37156
rect 11990 37100 12046 37156
rect 12114 37100 12170 37156
rect 12871 37100 12927 37156
rect 12995 37100 13051 37156
rect 13119 37100 13175 37156
rect 13243 37100 13299 37156
rect 13367 37100 13423 37156
rect 13491 37100 13547 37156
rect 13615 37100 13671 37156
rect 13739 37100 13795 37156
rect 13863 37100 13919 37156
rect 13987 37100 14043 37156
rect 14111 37100 14167 37156
rect 14235 37100 14291 37156
rect 14359 37100 14415 37156
rect 14483 37100 14539 37156
rect 14607 37100 14663 37156
rect 315 36976 371 37032
rect 439 36976 495 37032
rect 563 36976 619 37032
rect 687 36976 743 37032
rect 811 36976 867 37032
rect 935 36976 991 37032
rect 1059 36976 1115 37032
rect 1183 36976 1239 37032
rect 1307 36976 1363 37032
rect 1431 36976 1487 37032
rect 1555 36976 1611 37032
rect 1679 36976 1735 37032
rect 1803 36976 1859 37032
rect 1927 36976 1983 37032
rect 2051 36976 2107 37032
rect 2808 36976 2864 37032
rect 2932 36976 2988 37032
rect 3056 36976 3112 37032
rect 3180 36976 3236 37032
rect 3304 36976 3360 37032
rect 3428 36976 3484 37032
rect 3552 36976 3608 37032
rect 3676 36976 3732 37032
rect 3800 36976 3856 37032
rect 3924 36976 3980 37032
rect 4048 36976 4104 37032
rect 4172 36976 4228 37032
rect 4296 36976 4352 37032
rect 4420 36976 4476 37032
rect 4544 36976 4600 37032
rect 4668 36976 4724 37032
rect 5178 36976 5234 37032
rect 5302 36976 5358 37032
rect 5426 36976 5482 37032
rect 5550 36976 5606 37032
rect 5674 36976 5730 37032
rect 5798 36976 5854 37032
rect 5922 36976 5978 37032
rect 6046 36976 6102 37032
rect 6170 36976 6226 37032
rect 6294 36976 6350 37032
rect 6418 36976 6474 37032
rect 6542 36976 6598 37032
rect 6666 36976 6722 37032
rect 6790 36976 6846 37032
rect 6914 36976 6970 37032
rect 7038 36976 7094 37032
rect 7884 36976 7940 37032
rect 8008 36976 8064 37032
rect 8132 36976 8188 37032
rect 8256 36976 8312 37032
rect 8380 36976 8436 37032
rect 8504 36976 8560 37032
rect 8628 36976 8684 37032
rect 8752 36976 8808 37032
rect 8876 36976 8932 37032
rect 9000 36976 9056 37032
rect 9124 36976 9180 37032
rect 9248 36976 9304 37032
rect 9372 36976 9428 37032
rect 9496 36976 9552 37032
rect 9620 36976 9676 37032
rect 9744 36976 9800 37032
rect 10254 36976 10310 37032
rect 10378 36976 10434 37032
rect 10502 36976 10558 37032
rect 10626 36976 10682 37032
rect 10750 36976 10806 37032
rect 10874 36976 10930 37032
rect 10998 36976 11054 37032
rect 11122 36976 11178 37032
rect 11246 36976 11302 37032
rect 11370 36976 11426 37032
rect 11494 36976 11550 37032
rect 11618 36976 11674 37032
rect 11742 36976 11798 37032
rect 11866 36976 11922 37032
rect 11990 36976 12046 37032
rect 12114 36976 12170 37032
rect 12871 36976 12927 37032
rect 12995 36976 13051 37032
rect 13119 36976 13175 37032
rect 13243 36976 13299 37032
rect 13367 36976 13423 37032
rect 13491 36976 13547 37032
rect 13615 36976 13671 37032
rect 13739 36976 13795 37032
rect 13863 36976 13919 37032
rect 13987 36976 14043 37032
rect 14111 36976 14167 37032
rect 14235 36976 14291 37032
rect 14359 36976 14415 37032
rect 14483 36976 14539 37032
rect 14607 36976 14663 37032
rect 315 36852 371 36908
rect 439 36852 495 36908
rect 563 36852 619 36908
rect 687 36852 743 36908
rect 811 36852 867 36908
rect 935 36852 991 36908
rect 1059 36852 1115 36908
rect 1183 36852 1239 36908
rect 1307 36852 1363 36908
rect 1431 36852 1487 36908
rect 1555 36852 1611 36908
rect 1679 36852 1735 36908
rect 1803 36852 1859 36908
rect 1927 36852 1983 36908
rect 2051 36852 2107 36908
rect 2808 36852 2864 36908
rect 2932 36852 2988 36908
rect 3056 36852 3112 36908
rect 3180 36852 3236 36908
rect 3304 36852 3360 36908
rect 3428 36852 3484 36908
rect 3552 36852 3608 36908
rect 3676 36852 3732 36908
rect 3800 36852 3856 36908
rect 3924 36852 3980 36908
rect 4048 36852 4104 36908
rect 4172 36852 4228 36908
rect 4296 36852 4352 36908
rect 4420 36852 4476 36908
rect 4544 36852 4600 36908
rect 4668 36852 4724 36908
rect 5178 36852 5234 36908
rect 5302 36852 5358 36908
rect 5426 36852 5482 36908
rect 5550 36852 5606 36908
rect 5674 36852 5730 36908
rect 5798 36852 5854 36908
rect 5922 36852 5978 36908
rect 6046 36852 6102 36908
rect 6170 36852 6226 36908
rect 6294 36852 6350 36908
rect 6418 36852 6474 36908
rect 6542 36852 6598 36908
rect 6666 36852 6722 36908
rect 6790 36852 6846 36908
rect 6914 36852 6970 36908
rect 7038 36852 7094 36908
rect 7884 36852 7940 36908
rect 8008 36852 8064 36908
rect 8132 36852 8188 36908
rect 8256 36852 8312 36908
rect 8380 36852 8436 36908
rect 8504 36852 8560 36908
rect 8628 36852 8684 36908
rect 8752 36852 8808 36908
rect 8876 36852 8932 36908
rect 9000 36852 9056 36908
rect 9124 36852 9180 36908
rect 9248 36852 9304 36908
rect 9372 36852 9428 36908
rect 9496 36852 9552 36908
rect 9620 36852 9676 36908
rect 9744 36852 9800 36908
rect 10254 36852 10310 36908
rect 10378 36852 10434 36908
rect 10502 36852 10558 36908
rect 10626 36852 10682 36908
rect 10750 36852 10806 36908
rect 10874 36852 10930 36908
rect 10998 36852 11054 36908
rect 11122 36852 11178 36908
rect 11246 36852 11302 36908
rect 11370 36852 11426 36908
rect 11494 36852 11550 36908
rect 11618 36852 11674 36908
rect 11742 36852 11798 36908
rect 11866 36852 11922 36908
rect 11990 36852 12046 36908
rect 12114 36852 12170 36908
rect 12871 36852 12927 36908
rect 12995 36852 13051 36908
rect 13119 36852 13175 36908
rect 13243 36852 13299 36908
rect 13367 36852 13423 36908
rect 13491 36852 13547 36908
rect 13615 36852 13671 36908
rect 13739 36852 13795 36908
rect 13863 36852 13919 36908
rect 13987 36852 14043 36908
rect 14111 36852 14167 36908
rect 14235 36852 14291 36908
rect 14359 36852 14415 36908
rect 14483 36852 14539 36908
rect 14607 36852 14663 36908
rect 14902 38174 14958 38176
rect 14902 38122 14904 38174
rect 14904 38122 14956 38174
rect 14956 38122 14958 38174
rect 14902 38066 14958 38122
rect 14902 38014 14904 38066
rect 14904 38014 14956 38066
rect 14956 38014 14958 38066
rect 14902 37958 14958 38014
rect 14902 37906 14904 37958
rect 14904 37906 14956 37958
rect 14956 37906 14958 37958
rect 14902 37850 14958 37906
rect 14902 37798 14904 37850
rect 14904 37798 14956 37850
rect 14956 37798 14958 37850
rect 14902 37742 14958 37798
rect 14902 37690 14904 37742
rect 14904 37690 14956 37742
rect 14956 37690 14958 37742
rect 14902 37634 14958 37690
rect 14902 37582 14904 37634
rect 14904 37582 14956 37634
rect 14956 37582 14958 37634
rect 14902 37526 14958 37582
rect 14902 37474 14904 37526
rect 14904 37474 14956 37526
rect 14956 37474 14958 37526
rect 14902 37418 14958 37474
rect 14902 37366 14904 37418
rect 14904 37366 14956 37418
rect 14956 37366 14958 37418
rect 14902 37310 14958 37366
rect 14902 37258 14904 37310
rect 14904 37258 14956 37310
rect 14956 37258 14958 37310
rect 14902 37202 14958 37258
rect 14902 37150 14904 37202
rect 14904 37150 14956 37202
rect 14956 37150 14958 37202
rect 14902 37094 14958 37150
rect 14902 37042 14904 37094
rect 14904 37042 14956 37094
rect 14956 37042 14958 37094
rect 14902 36986 14958 37042
rect 14902 36934 14904 36986
rect 14904 36934 14956 36986
rect 14956 36934 14958 36986
rect 14902 36878 14958 36934
rect 14902 36826 14904 36878
rect 14904 36826 14956 36878
rect 14956 36826 14958 36878
rect 14902 36824 14958 36826
<< metal3 >>
rect 305 56043 2117 57235
rect 2798 56043 4734 57235
rect 5168 56043 7104 57235
rect 7874 56043 9810 57235
rect 10244 56043 12180 57235
rect 12861 56043 14673 57235
rect 2481 54442 2681 55758
rect 4851 54442 5051 55758
rect 7265 54442 7713 55758
rect 9927 54442 10127 55758
rect 12297 54442 12497 55758
rect 149 52830 14839 54180
rect 10 52580 86 52586
rect 14892 52580 14968 52586
rect 10 52576 14968 52580
rect 10 51224 20 52576
rect 76 52548 14902 52576
rect 76 52492 315 52548
rect 371 52492 439 52548
rect 495 52492 563 52548
rect 619 52492 687 52548
rect 743 52492 811 52548
rect 867 52492 935 52548
rect 991 52492 1059 52548
rect 1115 52492 1183 52548
rect 1239 52492 1307 52548
rect 1363 52492 1431 52548
rect 1487 52492 1555 52548
rect 1611 52492 1679 52548
rect 1735 52492 1803 52548
rect 1859 52492 1927 52548
rect 1983 52492 2051 52548
rect 2107 52492 2808 52548
rect 2864 52492 2932 52548
rect 2988 52492 3056 52548
rect 3112 52492 3180 52548
rect 3236 52492 3304 52548
rect 3360 52492 3428 52548
rect 3484 52492 3552 52548
rect 3608 52492 3676 52548
rect 3732 52492 3800 52548
rect 3856 52492 3924 52548
rect 3980 52492 4048 52548
rect 4104 52492 4172 52548
rect 4228 52492 4296 52548
rect 4352 52492 4420 52548
rect 4476 52492 4544 52548
rect 4600 52492 4668 52548
rect 4724 52492 5178 52548
rect 5234 52492 5302 52548
rect 5358 52492 5426 52548
rect 5482 52492 5550 52548
rect 5606 52492 5674 52548
rect 5730 52492 5798 52548
rect 5854 52492 5922 52548
rect 5978 52492 6046 52548
rect 6102 52492 6170 52548
rect 6226 52492 6294 52548
rect 6350 52492 6418 52548
rect 6474 52492 6542 52548
rect 6598 52492 6666 52548
rect 6722 52492 6790 52548
rect 6846 52492 6914 52548
rect 6970 52492 7038 52548
rect 7094 52492 7884 52548
rect 7940 52492 8008 52548
rect 8064 52492 8132 52548
rect 8188 52492 8256 52548
rect 8312 52492 8380 52548
rect 8436 52492 8504 52548
rect 8560 52492 8628 52548
rect 8684 52492 8752 52548
rect 8808 52492 8876 52548
rect 8932 52492 9000 52548
rect 9056 52492 9124 52548
rect 9180 52492 9248 52548
rect 9304 52492 9372 52548
rect 9428 52492 9496 52548
rect 9552 52492 9620 52548
rect 9676 52492 9744 52548
rect 9800 52492 10254 52548
rect 10310 52492 10378 52548
rect 10434 52492 10502 52548
rect 10558 52492 10626 52548
rect 10682 52492 10750 52548
rect 10806 52492 10874 52548
rect 10930 52492 10998 52548
rect 11054 52492 11122 52548
rect 11178 52492 11246 52548
rect 11302 52492 11370 52548
rect 11426 52492 11494 52548
rect 11550 52492 11618 52548
rect 11674 52492 11742 52548
rect 11798 52492 11866 52548
rect 11922 52492 11990 52548
rect 12046 52492 12114 52548
rect 12170 52492 12871 52548
rect 12927 52492 12995 52548
rect 13051 52492 13119 52548
rect 13175 52492 13243 52548
rect 13299 52492 13367 52548
rect 13423 52492 13491 52548
rect 13547 52492 13615 52548
rect 13671 52492 13739 52548
rect 13795 52492 13863 52548
rect 13919 52492 13987 52548
rect 14043 52492 14111 52548
rect 14167 52492 14235 52548
rect 14291 52492 14359 52548
rect 14415 52492 14483 52548
rect 14539 52492 14607 52548
rect 14663 52492 14902 52548
rect 76 52424 14902 52492
rect 76 52368 315 52424
rect 371 52368 439 52424
rect 495 52368 563 52424
rect 619 52368 687 52424
rect 743 52368 811 52424
rect 867 52368 935 52424
rect 991 52368 1059 52424
rect 1115 52368 1183 52424
rect 1239 52368 1307 52424
rect 1363 52368 1431 52424
rect 1487 52368 1555 52424
rect 1611 52368 1679 52424
rect 1735 52368 1803 52424
rect 1859 52368 1927 52424
rect 1983 52368 2051 52424
rect 2107 52368 2808 52424
rect 2864 52368 2932 52424
rect 2988 52368 3056 52424
rect 3112 52368 3180 52424
rect 3236 52368 3304 52424
rect 3360 52368 3428 52424
rect 3484 52368 3552 52424
rect 3608 52368 3676 52424
rect 3732 52368 3800 52424
rect 3856 52368 3924 52424
rect 3980 52368 4048 52424
rect 4104 52368 4172 52424
rect 4228 52368 4296 52424
rect 4352 52368 4420 52424
rect 4476 52368 4544 52424
rect 4600 52368 4668 52424
rect 4724 52368 5178 52424
rect 5234 52368 5302 52424
rect 5358 52368 5426 52424
rect 5482 52368 5550 52424
rect 5606 52368 5674 52424
rect 5730 52368 5798 52424
rect 5854 52368 5922 52424
rect 5978 52368 6046 52424
rect 6102 52368 6170 52424
rect 6226 52368 6294 52424
rect 6350 52368 6418 52424
rect 6474 52368 6542 52424
rect 6598 52368 6666 52424
rect 6722 52368 6790 52424
rect 6846 52368 6914 52424
rect 6970 52368 7038 52424
rect 7094 52368 7884 52424
rect 7940 52368 8008 52424
rect 8064 52368 8132 52424
rect 8188 52368 8256 52424
rect 8312 52368 8380 52424
rect 8436 52368 8504 52424
rect 8560 52368 8628 52424
rect 8684 52368 8752 52424
rect 8808 52368 8876 52424
rect 8932 52368 9000 52424
rect 9056 52368 9124 52424
rect 9180 52368 9248 52424
rect 9304 52368 9372 52424
rect 9428 52368 9496 52424
rect 9552 52368 9620 52424
rect 9676 52368 9744 52424
rect 9800 52368 10254 52424
rect 10310 52368 10378 52424
rect 10434 52368 10502 52424
rect 10558 52368 10626 52424
rect 10682 52368 10750 52424
rect 10806 52368 10874 52424
rect 10930 52368 10998 52424
rect 11054 52368 11122 52424
rect 11178 52368 11246 52424
rect 11302 52368 11370 52424
rect 11426 52368 11494 52424
rect 11550 52368 11618 52424
rect 11674 52368 11742 52424
rect 11798 52368 11866 52424
rect 11922 52368 11990 52424
rect 12046 52368 12114 52424
rect 12170 52368 12871 52424
rect 12927 52368 12995 52424
rect 13051 52368 13119 52424
rect 13175 52368 13243 52424
rect 13299 52368 13367 52424
rect 13423 52368 13491 52424
rect 13547 52368 13615 52424
rect 13671 52368 13739 52424
rect 13795 52368 13863 52424
rect 13919 52368 13987 52424
rect 14043 52368 14111 52424
rect 14167 52368 14235 52424
rect 14291 52368 14359 52424
rect 14415 52368 14483 52424
rect 14539 52368 14607 52424
rect 14663 52368 14902 52424
rect 76 52300 14902 52368
rect 76 52244 315 52300
rect 371 52244 439 52300
rect 495 52244 563 52300
rect 619 52244 687 52300
rect 743 52244 811 52300
rect 867 52244 935 52300
rect 991 52244 1059 52300
rect 1115 52244 1183 52300
rect 1239 52244 1307 52300
rect 1363 52244 1431 52300
rect 1487 52244 1555 52300
rect 1611 52244 1679 52300
rect 1735 52244 1803 52300
rect 1859 52244 1927 52300
rect 1983 52244 2051 52300
rect 2107 52244 2808 52300
rect 2864 52244 2932 52300
rect 2988 52244 3056 52300
rect 3112 52244 3180 52300
rect 3236 52244 3304 52300
rect 3360 52244 3428 52300
rect 3484 52244 3552 52300
rect 3608 52244 3676 52300
rect 3732 52244 3800 52300
rect 3856 52244 3924 52300
rect 3980 52244 4048 52300
rect 4104 52244 4172 52300
rect 4228 52244 4296 52300
rect 4352 52244 4420 52300
rect 4476 52244 4544 52300
rect 4600 52244 4668 52300
rect 4724 52244 5178 52300
rect 5234 52244 5302 52300
rect 5358 52244 5426 52300
rect 5482 52244 5550 52300
rect 5606 52244 5674 52300
rect 5730 52244 5798 52300
rect 5854 52244 5922 52300
rect 5978 52244 6046 52300
rect 6102 52244 6170 52300
rect 6226 52244 6294 52300
rect 6350 52244 6418 52300
rect 6474 52244 6542 52300
rect 6598 52244 6666 52300
rect 6722 52244 6790 52300
rect 6846 52244 6914 52300
rect 6970 52244 7038 52300
rect 7094 52244 7884 52300
rect 7940 52244 8008 52300
rect 8064 52244 8132 52300
rect 8188 52244 8256 52300
rect 8312 52244 8380 52300
rect 8436 52244 8504 52300
rect 8560 52244 8628 52300
rect 8684 52244 8752 52300
rect 8808 52244 8876 52300
rect 8932 52244 9000 52300
rect 9056 52244 9124 52300
rect 9180 52244 9248 52300
rect 9304 52244 9372 52300
rect 9428 52244 9496 52300
rect 9552 52244 9620 52300
rect 9676 52244 9744 52300
rect 9800 52244 10254 52300
rect 10310 52244 10378 52300
rect 10434 52244 10502 52300
rect 10558 52244 10626 52300
rect 10682 52244 10750 52300
rect 10806 52244 10874 52300
rect 10930 52244 10998 52300
rect 11054 52244 11122 52300
rect 11178 52244 11246 52300
rect 11302 52244 11370 52300
rect 11426 52244 11494 52300
rect 11550 52244 11618 52300
rect 11674 52244 11742 52300
rect 11798 52244 11866 52300
rect 11922 52244 11990 52300
rect 12046 52244 12114 52300
rect 12170 52244 12871 52300
rect 12927 52244 12995 52300
rect 13051 52244 13119 52300
rect 13175 52244 13243 52300
rect 13299 52244 13367 52300
rect 13423 52244 13491 52300
rect 13547 52244 13615 52300
rect 13671 52244 13739 52300
rect 13795 52244 13863 52300
rect 13919 52244 13987 52300
rect 14043 52244 14111 52300
rect 14167 52244 14235 52300
rect 14291 52244 14359 52300
rect 14415 52244 14483 52300
rect 14539 52244 14607 52300
rect 14663 52244 14902 52300
rect 76 52176 14902 52244
rect 76 52120 315 52176
rect 371 52120 439 52176
rect 495 52120 563 52176
rect 619 52120 687 52176
rect 743 52120 811 52176
rect 867 52120 935 52176
rect 991 52120 1059 52176
rect 1115 52120 1183 52176
rect 1239 52120 1307 52176
rect 1363 52120 1431 52176
rect 1487 52120 1555 52176
rect 1611 52120 1679 52176
rect 1735 52120 1803 52176
rect 1859 52120 1927 52176
rect 1983 52120 2051 52176
rect 2107 52120 2808 52176
rect 2864 52120 2932 52176
rect 2988 52120 3056 52176
rect 3112 52120 3180 52176
rect 3236 52120 3304 52176
rect 3360 52120 3428 52176
rect 3484 52120 3552 52176
rect 3608 52120 3676 52176
rect 3732 52120 3800 52176
rect 3856 52120 3924 52176
rect 3980 52120 4048 52176
rect 4104 52120 4172 52176
rect 4228 52120 4296 52176
rect 4352 52120 4420 52176
rect 4476 52120 4544 52176
rect 4600 52120 4668 52176
rect 4724 52120 5178 52176
rect 5234 52120 5302 52176
rect 5358 52120 5426 52176
rect 5482 52120 5550 52176
rect 5606 52120 5674 52176
rect 5730 52120 5798 52176
rect 5854 52120 5922 52176
rect 5978 52120 6046 52176
rect 6102 52120 6170 52176
rect 6226 52120 6294 52176
rect 6350 52120 6418 52176
rect 6474 52120 6542 52176
rect 6598 52120 6666 52176
rect 6722 52120 6790 52176
rect 6846 52120 6914 52176
rect 6970 52120 7038 52176
rect 7094 52120 7884 52176
rect 7940 52120 8008 52176
rect 8064 52120 8132 52176
rect 8188 52120 8256 52176
rect 8312 52120 8380 52176
rect 8436 52120 8504 52176
rect 8560 52120 8628 52176
rect 8684 52120 8752 52176
rect 8808 52120 8876 52176
rect 8932 52120 9000 52176
rect 9056 52120 9124 52176
rect 9180 52120 9248 52176
rect 9304 52120 9372 52176
rect 9428 52120 9496 52176
rect 9552 52120 9620 52176
rect 9676 52120 9744 52176
rect 9800 52120 10254 52176
rect 10310 52120 10378 52176
rect 10434 52120 10502 52176
rect 10558 52120 10626 52176
rect 10682 52120 10750 52176
rect 10806 52120 10874 52176
rect 10930 52120 10998 52176
rect 11054 52120 11122 52176
rect 11178 52120 11246 52176
rect 11302 52120 11370 52176
rect 11426 52120 11494 52176
rect 11550 52120 11618 52176
rect 11674 52120 11742 52176
rect 11798 52120 11866 52176
rect 11922 52120 11990 52176
rect 12046 52120 12114 52176
rect 12170 52120 12871 52176
rect 12927 52120 12995 52176
rect 13051 52120 13119 52176
rect 13175 52120 13243 52176
rect 13299 52120 13367 52176
rect 13423 52120 13491 52176
rect 13547 52120 13615 52176
rect 13671 52120 13739 52176
rect 13795 52120 13863 52176
rect 13919 52120 13987 52176
rect 14043 52120 14111 52176
rect 14167 52120 14235 52176
rect 14291 52120 14359 52176
rect 14415 52120 14483 52176
rect 14539 52120 14607 52176
rect 14663 52120 14902 52176
rect 76 52052 14902 52120
rect 76 51996 315 52052
rect 371 51996 439 52052
rect 495 51996 563 52052
rect 619 51996 687 52052
rect 743 51996 811 52052
rect 867 51996 935 52052
rect 991 51996 1059 52052
rect 1115 51996 1183 52052
rect 1239 51996 1307 52052
rect 1363 51996 1431 52052
rect 1487 51996 1555 52052
rect 1611 51996 1679 52052
rect 1735 51996 1803 52052
rect 1859 51996 1927 52052
rect 1983 51996 2051 52052
rect 2107 51996 2808 52052
rect 2864 51996 2932 52052
rect 2988 51996 3056 52052
rect 3112 51996 3180 52052
rect 3236 51996 3304 52052
rect 3360 51996 3428 52052
rect 3484 51996 3552 52052
rect 3608 51996 3676 52052
rect 3732 51996 3800 52052
rect 3856 51996 3924 52052
rect 3980 51996 4048 52052
rect 4104 51996 4172 52052
rect 4228 51996 4296 52052
rect 4352 51996 4420 52052
rect 4476 51996 4544 52052
rect 4600 51996 4668 52052
rect 4724 51996 5178 52052
rect 5234 51996 5302 52052
rect 5358 51996 5426 52052
rect 5482 51996 5550 52052
rect 5606 51996 5674 52052
rect 5730 51996 5798 52052
rect 5854 51996 5922 52052
rect 5978 51996 6046 52052
rect 6102 51996 6170 52052
rect 6226 51996 6294 52052
rect 6350 51996 6418 52052
rect 6474 51996 6542 52052
rect 6598 51996 6666 52052
rect 6722 51996 6790 52052
rect 6846 51996 6914 52052
rect 6970 51996 7038 52052
rect 7094 51996 7884 52052
rect 7940 51996 8008 52052
rect 8064 51996 8132 52052
rect 8188 51996 8256 52052
rect 8312 51996 8380 52052
rect 8436 51996 8504 52052
rect 8560 51996 8628 52052
rect 8684 51996 8752 52052
rect 8808 51996 8876 52052
rect 8932 51996 9000 52052
rect 9056 51996 9124 52052
rect 9180 51996 9248 52052
rect 9304 51996 9372 52052
rect 9428 51996 9496 52052
rect 9552 51996 9620 52052
rect 9676 51996 9744 52052
rect 9800 51996 10254 52052
rect 10310 51996 10378 52052
rect 10434 51996 10502 52052
rect 10558 51996 10626 52052
rect 10682 51996 10750 52052
rect 10806 51996 10874 52052
rect 10930 51996 10998 52052
rect 11054 51996 11122 52052
rect 11178 51996 11246 52052
rect 11302 51996 11370 52052
rect 11426 51996 11494 52052
rect 11550 51996 11618 52052
rect 11674 51996 11742 52052
rect 11798 51996 11866 52052
rect 11922 51996 11990 52052
rect 12046 51996 12114 52052
rect 12170 51996 12871 52052
rect 12927 51996 12995 52052
rect 13051 51996 13119 52052
rect 13175 51996 13243 52052
rect 13299 51996 13367 52052
rect 13423 51996 13491 52052
rect 13547 51996 13615 52052
rect 13671 51996 13739 52052
rect 13795 51996 13863 52052
rect 13919 51996 13987 52052
rect 14043 51996 14111 52052
rect 14167 51996 14235 52052
rect 14291 51996 14359 52052
rect 14415 51996 14483 52052
rect 14539 51996 14607 52052
rect 14663 51996 14902 52052
rect 76 51928 14902 51996
rect 76 51872 315 51928
rect 371 51872 439 51928
rect 495 51872 563 51928
rect 619 51872 687 51928
rect 743 51872 811 51928
rect 867 51872 935 51928
rect 991 51872 1059 51928
rect 1115 51872 1183 51928
rect 1239 51872 1307 51928
rect 1363 51872 1431 51928
rect 1487 51872 1555 51928
rect 1611 51872 1679 51928
rect 1735 51872 1803 51928
rect 1859 51872 1927 51928
rect 1983 51872 2051 51928
rect 2107 51872 2808 51928
rect 2864 51872 2932 51928
rect 2988 51872 3056 51928
rect 3112 51872 3180 51928
rect 3236 51872 3304 51928
rect 3360 51872 3428 51928
rect 3484 51872 3552 51928
rect 3608 51872 3676 51928
rect 3732 51872 3800 51928
rect 3856 51872 3924 51928
rect 3980 51872 4048 51928
rect 4104 51872 4172 51928
rect 4228 51872 4296 51928
rect 4352 51872 4420 51928
rect 4476 51872 4544 51928
rect 4600 51872 4668 51928
rect 4724 51872 5178 51928
rect 5234 51872 5302 51928
rect 5358 51872 5426 51928
rect 5482 51872 5550 51928
rect 5606 51872 5674 51928
rect 5730 51872 5798 51928
rect 5854 51872 5922 51928
rect 5978 51872 6046 51928
rect 6102 51872 6170 51928
rect 6226 51872 6294 51928
rect 6350 51872 6418 51928
rect 6474 51872 6542 51928
rect 6598 51872 6666 51928
rect 6722 51872 6790 51928
rect 6846 51872 6914 51928
rect 6970 51872 7038 51928
rect 7094 51872 7884 51928
rect 7940 51872 8008 51928
rect 8064 51872 8132 51928
rect 8188 51872 8256 51928
rect 8312 51872 8380 51928
rect 8436 51872 8504 51928
rect 8560 51872 8628 51928
rect 8684 51872 8752 51928
rect 8808 51872 8876 51928
rect 8932 51872 9000 51928
rect 9056 51872 9124 51928
rect 9180 51872 9248 51928
rect 9304 51872 9372 51928
rect 9428 51872 9496 51928
rect 9552 51872 9620 51928
rect 9676 51872 9744 51928
rect 9800 51872 10254 51928
rect 10310 51872 10378 51928
rect 10434 51872 10502 51928
rect 10558 51872 10626 51928
rect 10682 51872 10750 51928
rect 10806 51872 10874 51928
rect 10930 51872 10998 51928
rect 11054 51872 11122 51928
rect 11178 51872 11246 51928
rect 11302 51872 11370 51928
rect 11426 51872 11494 51928
rect 11550 51872 11618 51928
rect 11674 51872 11742 51928
rect 11798 51872 11866 51928
rect 11922 51872 11990 51928
rect 12046 51872 12114 51928
rect 12170 51872 12871 51928
rect 12927 51872 12995 51928
rect 13051 51872 13119 51928
rect 13175 51872 13243 51928
rect 13299 51872 13367 51928
rect 13423 51872 13491 51928
rect 13547 51872 13615 51928
rect 13671 51872 13739 51928
rect 13795 51872 13863 51928
rect 13919 51872 13987 51928
rect 14043 51872 14111 51928
rect 14167 51872 14235 51928
rect 14291 51872 14359 51928
rect 14415 51872 14483 51928
rect 14539 51872 14607 51928
rect 14663 51872 14902 51928
rect 76 51804 14902 51872
rect 76 51748 315 51804
rect 371 51748 439 51804
rect 495 51748 563 51804
rect 619 51748 687 51804
rect 743 51748 811 51804
rect 867 51748 935 51804
rect 991 51748 1059 51804
rect 1115 51748 1183 51804
rect 1239 51748 1307 51804
rect 1363 51748 1431 51804
rect 1487 51748 1555 51804
rect 1611 51748 1679 51804
rect 1735 51748 1803 51804
rect 1859 51748 1927 51804
rect 1983 51748 2051 51804
rect 2107 51748 2808 51804
rect 2864 51748 2932 51804
rect 2988 51748 3056 51804
rect 3112 51748 3180 51804
rect 3236 51748 3304 51804
rect 3360 51748 3428 51804
rect 3484 51748 3552 51804
rect 3608 51748 3676 51804
rect 3732 51748 3800 51804
rect 3856 51748 3924 51804
rect 3980 51748 4048 51804
rect 4104 51748 4172 51804
rect 4228 51748 4296 51804
rect 4352 51748 4420 51804
rect 4476 51748 4544 51804
rect 4600 51748 4668 51804
rect 4724 51748 5178 51804
rect 5234 51748 5302 51804
rect 5358 51748 5426 51804
rect 5482 51748 5550 51804
rect 5606 51748 5674 51804
rect 5730 51748 5798 51804
rect 5854 51748 5922 51804
rect 5978 51748 6046 51804
rect 6102 51748 6170 51804
rect 6226 51748 6294 51804
rect 6350 51748 6418 51804
rect 6474 51748 6542 51804
rect 6598 51748 6666 51804
rect 6722 51748 6790 51804
rect 6846 51748 6914 51804
rect 6970 51748 7038 51804
rect 7094 51748 7884 51804
rect 7940 51748 8008 51804
rect 8064 51748 8132 51804
rect 8188 51748 8256 51804
rect 8312 51748 8380 51804
rect 8436 51748 8504 51804
rect 8560 51748 8628 51804
rect 8684 51748 8752 51804
rect 8808 51748 8876 51804
rect 8932 51748 9000 51804
rect 9056 51748 9124 51804
rect 9180 51748 9248 51804
rect 9304 51748 9372 51804
rect 9428 51748 9496 51804
rect 9552 51748 9620 51804
rect 9676 51748 9744 51804
rect 9800 51748 10254 51804
rect 10310 51748 10378 51804
rect 10434 51748 10502 51804
rect 10558 51748 10626 51804
rect 10682 51748 10750 51804
rect 10806 51748 10874 51804
rect 10930 51748 10998 51804
rect 11054 51748 11122 51804
rect 11178 51748 11246 51804
rect 11302 51748 11370 51804
rect 11426 51748 11494 51804
rect 11550 51748 11618 51804
rect 11674 51748 11742 51804
rect 11798 51748 11866 51804
rect 11922 51748 11990 51804
rect 12046 51748 12114 51804
rect 12170 51748 12871 51804
rect 12927 51748 12995 51804
rect 13051 51748 13119 51804
rect 13175 51748 13243 51804
rect 13299 51748 13367 51804
rect 13423 51748 13491 51804
rect 13547 51748 13615 51804
rect 13671 51748 13739 51804
rect 13795 51748 13863 51804
rect 13919 51748 13987 51804
rect 14043 51748 14111 51804
rect 14167 51748 14235 51804
rect 14291 51748 14359 51804
rect 14415 51748 14483 51804
rect 14539 51748 14607 51804
rect 14663 51748 14902 51804
rect 76 51680 14902 51748
rect 76 51624 315 51680
rect 371 51624 439 51680
rect 495 51624 563 51680
rect 619 51624 687 51680
rect 743 51624 811 51680
rect 867 51624 935 51680
rect 991 51624 1059 51680
rect 1115 51624 1183 51680
rect 1239 51624 1307 51680
rect 1363 51624 1431 51680
rect 1487 51624 1555 51680
rect 1611 51624 1679 51680
rect 1735 51624 1803 51680
rect 1859 51624 1927 51680
rect 1983 51624 2051 51680
rect 2107 51624 2808 51680
rect 2864 51624 2932 51680
rect 2988 51624 3056 51680
rect 3112 51624 3180 51680
rect 3236 51624 3304 51680
rect 3360 51624 3428 51680
rect 3484 51624 3552 51680
rect 3608 51624 3676 51680
rect 3732 51624 3800 51680
rect 3856 51624 3924 51680
rect 3980 51624 4048 51680
rect 4104 51624 4172 51680
rect 4228 51624 4296 51680
rect 4352 51624 4420 51680
rect 4476 51624 4544 51680
rect 4600 51624 4668 51680
rect 4724 51624 5178 51680
rect 5234 51624 5302 51680
rect 5358 51624 5426 51680
rect 5482 51624 5550 51680
rect 5606 51624 5674 51680
rect 5730 51624 5798 51680
rect 5854 51624 5922 51680
rect 5978 51624 6046 51680
rect 6102 51624 6170 51680
rect 6226 51624 6294 51680
rect 6350 51624 6418 51680
rect 6474 51624 6542 51680
rect 6598 51624 6666 51680
rect 6722 51624 6790 51680
rect 6846 51624 6914 51680
rect 6970 51624 7038 51680
rect 7094 51624 7884 51680
rect 7940 51624 8008 51680
rect 8064 51624 8132 51680
rect 8188 51624 8256 51680
rect 8312 51624 8380 51680
rect 8436 51624 8504 51680
rect 8560 51624 8628 51680
rect 8684 51624 8752 51680
rect 8808 51624 8876 51680
rect 8932 51624 9000 51680
rect 9056 51624 9124 51680
rect 9180 51624 9248 51680
rect 9304 51624 9372 51680
rect 9428 51624 9496 51680
rect 9552 51624 9620 51680
rect 9676 51624 9744 51680
rect 9800 51624 10254 51680
rect 10310 51624 10378 51680
rect 10434 51624 10502 51680
rect 10558 51624 10626 51680
rect 10682 51624 10750 51680
rect 10806 51624 10874 51680
rect 10930 51624 10998 51680
rect 11054 51624 11122 51680
rect 11178 51624 11246 51680
rect 11302 51624 11370 51680
rect 11426 51624 11494 51680
rect 11550 51624 11618 51680
rect 11674 51624 11742 51680
rect 11798 51624 11866 51680
rect 11922 51624 11990 51680
rect 12046 51624 12114 51680
rect 12170 51624 12871 51680
rect 12927 51624 12995 51680
rect 13051 51624 13119 51680
rect 13175 51624 13243 51680
rect 13299 51624 13367 51680
rect 13423 51624 13491 51680
rect 13547 51624 13615 51680
rect 13671 51624 13739 51680
rect 13795 51624 13863 51680
rect 13919 51624 13987 51680
rect 14043 51624 14111 51680
rect 14167 51624 14235 51680
rect 14291 51624 14359 51680
rect 14415 51624 14483 51680
rect 14539 51624 14607 51680
rect 14663 51624 14902 51680
rect 76 51556 14902 51624
rect 76 51500 315 51556
rect 371 51500 439 51556
rect 495 51500 563 51556
rect 619 51500 687 51556
rect 743 51500 811 51556
rect 867 51500 935 51556
rect 991 51500 1059 51556
rect 1115 51500 1183 51556
rect 1239 51500 1307 51556
rect 1363 51500 1431 51556
rect 1487 51500 1555 51556
rect 1611 51500 1679 51556
rect 1735 51500 1803 51556
rect 1859 51500 1927 51556
rect 1983 51500 2051 51556
rect 2107 51500 2808 51556
rect 2864 51500 2932 51556
rect 2988 51500 3056 51556
rect 3112 51500 3180 51556
rect 3236 51500 3304 51556
rect 3360 51500 3428 51556
rect 3484 51500 3552 51556
rect 3608 51500 3676 51556
rect 3732 51500 3800 51556
rect 3856 51500 3924 51556
rect 3980 51500 4048 51556
rect 4104 51500 4172 51556
rect 4228 51500 4296 51556
rect 4352 51500 4420 51556
rect 4476 51500 4544 51556
rect 4600 51500 4668 51556
rect 4724 51500 5178 51556
rect 5234 51500 5302 51556
rect 5358 51500 5426 51556
rect 5482 51500 5550 51556
rect 5606 51500 5674 51556
rect 5730 51500 5798 51556
rect 5854 51500 5922 51556
rect 5978 51500 6046 51556
rect 6102 51500 6170 51556
rect 6226 51500 6294 51556
rect 6350 51500 6418 51556
rect 6474 51500 6542 51556
rect 6598 51500 6666 51556
rect 6722 51500 6790 51556
rect 6846 51500 6914 51556
rect 6970 51500 7038 51556
rect 7094 51500 7884 51556
rect 7940 51500 8008 51556
rect 8064 51500 8132 51556
rect 8188 51500 8256 51556
rect 8312 51500 8380 51556
rect 8436 51500 8504 51556
rect 8560 51500 8628 51556
rect 8684 51500 8752 51556
rect 8808 51500 8876 51556
rect 8932 51500 9000 51556
rect 9056 51500 9124 51556
rect 9180 51500 9248 51556
rect 9304 51500 9372 51556
rect 9428 51500 9496 51556
rect 9552 51500 9620 51556
rect 9676 51500 9744 51556
rect 9800 51500 10254 51556
rect 10310 51500 10378 51556
rect 10434 51500 10502 51556
rect 10558 51500 10626 51556
rect 10682 51500 10750 51556
rect 10806 51500 10874 51556
rect 10930 51500 10998 51556
rect 11054 51500 11122 51556
rect 11178 51500 11246 51556
rect 11302 51500 11370 51556
rect 11426 51500 11494 51556
rect 11550 51500 11618 51556
rect 11674 51500 11742 51556
rect 11798 51500 11866 51556
rect 11922 51500 11990 51556
rect 12046 51500 12114 51556
rect 12170 51500 12871 51556
rect 12927 51500 12995 51556
rect 13051 51500 13119 51556
rect 13175 51500 13243 51556
rect 13299 51500 13367 51556
rect 13423 51500 13491 51556
rect 13547 51500 13615 51556
rect 13671 51500 13739 51556
rect 13795 51500 13863 51556
rect 13919 51500 13987 51556
rect 14043 51500 14111 51556
rect 14167 51500 14235 51556
rect 14291 51500 14359 51556
rect 14415 51500 14483 51556
rect 14539 51500 14607 51556
rect 14663 51500 14902 51556
rect 76 51432 14902 51500
rect 76 51376 315 51432
rect 371 51376 439 51432
rect 495 51376 563 51432
rect 619 51376 687 51432
rect 743 51376 811 51432
rect 867 51376 935 51432
rect 991 51376 1059 51432
rect 1115 51376 1183 51432
rect 1239 51376 1307 51432
rect 1363 51376 1431 51432
rect 1487 51376 1555 51432
rect 1611 51376 1679 51432
rect 1735 51376 1803 51432
rect 1859 51376 1927 51432
rect 1983 51376 2051 51432
rect 2107 51376 2808 51432
rect 2864 51376 2932 51432
rect 2988 51376 3056 51432
rect 3112 51376 3180 51432
rect 3236 51376 3304 51432
rect 3360 51376 3428 51432
rect 3484 51376 3552 51432
rect 3608 51376 3676 51432
rect 3732 51376 3800 51432
rect 3856 51376 3924 51432
rect 3980 51376 4048 51432
rect 4104 51376 4172 51432
rect 4228 51376 4296 51432
rect 4352 51376 4420 51432
rect 4476 51376 4544 51432
rect 4600 51376 4668 51432
rect 4724 51376 5178 51432
rect 5234 51376 5302 51432
rect 5358 51376 5426 51432
rect 5482 51376 5550 51432
rect 5606 51376 5674 51432
rect 5730 51376 5798 51432
rect 5854 51376 5922 51432
rect 5978 51376 6046 51432
rect 6102 51376 6170 51432
rect 6226 51376 6294 51432
rect 6350 51376 6418 51432
rect 6474 51376 6542 51432
rect 6598 51376 6666 51432
rect 6722 51376 6790 51432
rect 6846 51376 6914 51432
rect 6970 51376 7038 51432
rect 7094 51376 7884 51432
rect 7940 51376 8008 51432
rect 8064 51376 8132 51432
rect 8188 51376 8256 51432
rect 8312 51376 8380 51432
rect 8436 51376 8504 51432
rect 8560 51376 8628 51432
rect 8684 51376 8752 51432
rect 8808 51376 8876 51432
rect 8932 51376 9000 51432
rect 9056 51376 9124 51432
rect 9180 51376 9248 51432
rect 9304 51376 9372 51432
rect 9428 51376 9496 51432
rect 9552 51376 9620 51432
rect 9676 51376 9744 51432
rect 9800 51376 10254 51432
rect 10310 51376 10378 51432
rect 10434 51376 10502 51432
rect 10558 51376 10626 51432
rect 10682 51376 10750 51432
rect 10806 51376 10874 51432
rect 10930 51376 10998 51432
rect 11054 51376 11122 51432
rect 11178 51376 11246 51432
rect 11302 51376 11370 51432
rect 11426 51376 11494 51432
rect 11550 51376 11618 51432
rect 11674 51376 11742 51432
rect 11798 51376 11866 51432
rect 11922 51376 11990 51432
rect 12046 51376 12114 51432
rect 12170 51376 12871 51432
rect 12927 51376 12995 51432
rect 13051 51376 13119 51432
rect 13175 51376 13243 51432
rect 13299 51376 13367 51432
rect 13423 51376 13491 51432
rect 13547 51376 13615 51432
rect 13671 51376 13739 51432
rect 13795 51376 13863 51432
rect 13919 51376 13987 51432
rect 14043 51376 14111 51432
rect 14167 51376 14235 51432
rect 14291 51376 14359 51432
rect 14415 51376 14483 51432
rect 14539 51376 14607 51432
rect 14663 51376 14902 51432
rect 76 51308 14902 51376
rect 76 51252 315 51308
rect 371 51252 439 51308
rect 495 51252 563 51308
rect 619 51252 687 51308
rect 743 51252 811 51308
rect 867 51252 935 51308
rect 991 51252 1059 51308
rect 1115 51252 1183 51308
rect 1239 51252 1307 51308
rect 1363 51252 1431 51308
rect 1487 51252 1555 51308
rect 1611 51252 1679 51308
rect 1735 51252 1803 51308
rect 1859 51252 1927 51308
rect 1983 51252 2051 51308
rect 2107 51252 2808 51308
rect 2864 51252 2932 51308
rect 2988 51252 3056 51308
rect 3112 51252 3180 51308
rect 3236 51252 3304 51308
rect 3360 51252 3428 51308
rect 3484 51252 3552 51308
rect 3608 51252 3676 51308
rect 3732 51252 3800 51308
rect 3856 51252 3924 51308
rect 3980 51252 4048 51308
rect 4104 51252 4172 51308
rect 4228 51252 4296 51308
rect 4352 51252 4420 51308
rect 4476 51252 4544 51308
rect 4600 51252 4668 51308
rect 4724 51252 5178 51308
rect 5234 51252 5302 51308
rect 5358 51252 5426 51308
rect 5482 51252 5550 51308
rect 5606 51252 5674 51308
rect 5730 51252 5798 51308
rect 5854 51252 5922 51308
rect 5978 51252 6046 51308
rect 6102 51252 6170 51308
rect 6226 51252 6294 51308
rect 6350 51252 6418 51308
rect 6474 51252 6542 51308
rect 6598 51252 6666 51308
rect 6722 51252 6790 51308
rect 6846 51252 6914 51308
rect 6970 51252 7038 51308
rect 7094 51252 7884 51308
rect 7940 51252 8008 51308
rect 8064 51252 8132 51308
rect 8188 51252 8256 51308
rect 8312 51252 8380 51308
rect 8436 51252 8504 51308
rect 8560 51252 8628 51308
rect 8684 51252 8752 51308
rect 8808 51252 8876 51308
rect 8932 51252 9000 51308
rect 9056 51252 9124 51308
rect 9180 51252 9248 51308
rect 9304 51252 9372 51308
rect 9428 51252 9496 51308
rect 9552 51252 9620 51308
rect 9676 51252 9744 51308
rect 9800 51252 10254 51308
rect 10310 51252 10378 51308
rect 10434 51252 10502 51308
rect 10558 51252 10626 51308
rect 10682 51252 10750 51308
rect 10806 51252 10874 51308
rect 10930 51252 10998 51308
rect 11054 51252 11122 51308
rect 11178 51252 11246 51308
rect 11302 51252 11370 51308
rect 11426 51252 11494 51308
rect 11550 51252 11618 51308
rect 11674 51252 11742 51308
rect 11798 51252 11866 51308
rect 11922 51252 11990 51308
rect 12046 51252 12114 51308
rect 12170 51252 12871 51308
rect 12927 51252 12995 51308
rect 13051 51252 13119 51308
rect 13175 51252 13243 51308
rect 13299 51252 13367 51308
rect 13423 51252 13491 51308
rect 13547 51252 13615 51308
rect 13671 51252 13739 51308
rect 13795 51252 13863 51308
rect 13919 51252 13987 51308
rect 14043 51252 14111 51308
rect 14167 51252 14235 51308
rect 14291 51252 14359 51308
rect 14415 51252 14483 51308
rect 14539 51252 14607 51308
rect 14663 51252 14902 51308
rect 76 51230 14902 51252
rect 76 51224 86 51230
rect 10 51214 86 51224
rect 14892 51224 14902 51230
rect 14958 51224 14968 52576
rect 14892 51214 14968 51224
rect 2481 50948 2681 50958
rect 2292 50926 2368 50936
rect 2292 50870 2302 50926
rect 2358 50870 2368 50926
rect 2292 50794 2368 50870
rect 2292 50738 2302 50794
rect 2358 50738 2368 50794
rect 2292 50662 2368 50738
rect 2292 50606 2302 50662
rect 2358 50606 2368 50662
rect 2292 50530 2368 50606
rect 2292 50474 2302 50530
rect 2358 50474 2368 50530
rect 2292 50398 2368 50474
rect 2292 50342 2302 50398
rect 2358 50342 2368 50398
rect 2292 50266 2368 50342
rect 2292 50210 2302 50266
rect 2358 50210 2368 50266
rect 2292 50134 2368 50210
rect 2292 50078 2302 50134
rect 2358 50078 2368 50134
rect 2292 50002 2368 50078
rect 2292 49946 2302 50002
rect 2358 49946 2368 50002
rect 2292 49870 2368 49946
rect 2292 49814 2302 49870
rect 2358 49814 2368 49870
rect 2292 49738 2368 49814
rect 2292 49682 2302 49738
rect 2358 49682 2368 49738
rect 2292 49672 2368 49682
rect 2481 50892 2491 50948
rect 2547 50892 2615 50948
rect 2671 50892 2681 50948
rect 2481 50824 2681 50892
rect 2481 50768 2491 50824
rect 2547 50768 2615 50824
rect 2671 50768 2681 50824
rect 2481 50700 2681 50768
rect 2481 50644 2491 50700
rect 2547 50644 2615 50700
rect 2671 50644 2681 50700
rect 2481 50576 2681 50644
rect 2481 50520 2491 50576
rect 2547 50520 2615 50576
rect 2671 50520 2681 50576
rect 2481 50452 2681 50520
rect 2481 50396 2491 50452
rect 2547 50396 2615 50452
rect 2671 50396 2681 50452
rect 2481 50328 2681 50396
rect 2481 50272 2491 50328
rect 2547 50272 2615 50328
rect 2671 50272 2681 50328
rect 2481 50204 2681 50272
rect 2481 50148 2491 50204
rect 2547 50148 2615 50204
rect 2671 50148 2681 50204
rect 2481 50080 2681 50148
rect 2481 50024 2491 50080
rect 2547 50024 2615 50080
rect 2671 50024 2681 50080
rect 2481 49956 2681 50024
rect 2481 49900 2491 49956
rect 2547 49900 2615 49956
rect 2671 49900 2681 49956
rect 2481 49832 2681 49900
rect 2481 49776 2491 49832
rect 2547 49776 2615 49832
rect 2671 49776 2681 49832
rect 2481 49708 2681 49776
rect 2481 49652 2491 49708
rect 2547 49652 2615 49708
rect 2671 49652 2681 49708
rect 2481 49642 2681 49652
rect 4851 50948 5051 50958
rect 4851 50892 4861 50948
rect 4917 50892 4985 50948
rect 5041 50892 5051 50948
rect 4851 50824 5051 50892
rect 4851 50768 4861 50824
rect 4917 50768 4985 50824
rect 5041 50768 5051 50824
rect 4851 50700 5051 50768
rect 4851 50644 4861 50700
rect 4917 50644 4985 50700
rect 5041 50644 5051 50700
rect 4851 50576 5051 50644
rect 4851 50520 4861 50576
rect 4917 50520 4985 50576
rect 5041 50520 5051 50576
rect 4851 50452 5051 50520
rect 4851 50396 4861 50452
rect 4917 50396 4985 50452
rect 5041 50396 5051 50452
rect 4851 50328 5051 50396
rect 4851 50272 4861 50328
rect 4917 50272 4985 50328
rect 5041 50272 5051 50328
rect 4851 50204 5051 50272
rect 4851 50148 4861 50204
rect 4917 50148 4985 50204
rect 5041 50148 5051 50204
rect 4851 50080 5051 50148
rect 4851 50024 4861 50080
rect 4917 50024 4985 50080
rect 5041 50024 5051 50080
rect 4851 49956 5051 50024
rect 4851 49900 4861 49956
rect 4917 49900 4985 49956
rect 5041 49900 5051 49956
rect 4851 49832 5051 49900
rect 4851 49776 4861 49832
rect 4917 49776 4985 49832
rect 5041 49776 5051 49832
rect 4851 49708 5051 49776
rect 4851 49652 4861 49708
rect 4917 49652 4985 49708
rect 5041 49652 5051 49708
rect 4851 49642 5051 49652
rect 7265 50948 7713 50958
rect 7265 50892 7275 50948
rect 7331 50892 7399 50948
rect 7455 50892 7523 50948
rect 7579 50892 7647 50948
rect 7703 50892 7713 50948
rect 7265 50824 7713 50892
rect 7265 50768 7275 50824
rect 7331 50768 7399 50824
rect 7455 50768 7523 50824
rect 7579 50768 7647 50824
rect 7703 50768 7713 50824
rect 7265 50700 7713 50768
rect 7265 50644 7275 50700
rect 7331 50644 7399 50700
rect 7455 50644 7523 50700
rect 7579 50644 7647 50700
rect 7703 50644 7713 50700
rect 7265 50576 7713 50644
rect 7265 50520 7275 50576
rect 7331 50520 7399 50576
rect 7455 50520 7523 50576
rect 7579 50520 7647 50576
rect 7703 50520 7713 50576
rect 7265 50452 7713 50520
rect 7265 50396 7275 50452
rect 7331 50396 7399 50452
rect 7455 50396 7523 50452
rect 7579 50396 7647 50452
rect 7703 50396 7713 50452
rect 7265 50328 7713 50396
rect 7265 50272 7275 50328
rect 7331 50272 7399 50328
rect 7455 50272 7523 50328
rect 7579 50272 7647 50328
rect 7703 50272 7713 50328
rect 7265 50204 7713 50272
rect 7265 50148 7275 50204
rect 7331 50148 7399 50204
rect 7455 50148 7523 50204
rect 7579 50148 7647 50204
rect 7703 50148 7713 50204
rect 7265 50080 7713 50148
rect 7265 50024 7275 50080
rect 7331 50024 7399 50080
rect 7455 50024 7523 50080
rect 7579 50024 7647 50080
rect 7703 50024 7713 50080
rect 7265 49956 7713 50024
rect 7265 49900 7275 49956
rect 7331 49900 7399 49956
rect 7455 49900 7523 49956
rect 7579 49900 7647 49956
rect 7703 49900 7713 49956
rect 7265 49832 7713 49900
rect 7265 49776 7275 49832
rect 7331 49776 7399 49832
rect 7455 49776 7523 49832
rect 7579 49776 7647 49832
rect 7703 49776 7713 49832
rect 7265 49708 7713 49776
rect 7265 49652 7275 49708
rect 7331 49652 7399 49708
rect 7455 49652 7523 49708
rect 7579 49652 7647 49708
rect 7703 49652 7713 49708
rect 7265 49642 7713 49652
rect 9927 50948 10127 50958
rect 9927 50892 9937 50948
rect 9993 50892 10061 50948
rect 10117 50892 10127 50948
rect 9927 50824 10127 50892
rect 9927 50768 9937 50824
rect 9993 50768 10061 50824
rect 10117 50768 10127 50824
rect 9927 50700 10127 50768
rect 9927 50644 9937 50700
rect 9993 50644 10061 50700
rect 10117 50644 10127 50700
rect 9927 50576 10127 50644
rect 9927 50520 9937 50576
rect 9993 50520 10061 50576
rect 10117 50520 10127 50576
rect 9927 50452 10127 50520
rect 9927 50396 9937 50452
rect 9993 50396 10061 50452
rect 10117 50396 10127 50452
rect 9927 50328 10127 50396
rect 9927 50272 9937 50328
rect 9993 50272 10061 50328
rect 10117 50272 10127 50328
rect 9927 50204 10127 50272
rect 9927 50148 9937 50204
rect 9993 50148 10061 50204
rect 10117 50148 10127 50204
rect 9927 50080 10127 50148
rect 9927 50024 9937 50080
rect 9993 50024 10061 50080
rect 10117 50024 10127 50080
rect 9927 49956 10127 50024
rect 9927 49900 9937 49956
rect 9993 49900 10061 49956
rect 10117 49900 10127 49956
rect 9927 49832 10127 49900
rect 9927 49776 9937 49832
rect 9993 49776 10061 49832
rect 10117 49776 10127 49832
rect 9927 49708 10127 49776
rect 9927 49652 9937 49708
rect 9993 49652 10061 49708
rect 10117 49652 10127 49708
rect 9927 49642 10127 49652
rect 12297 50948 12497 50958
rect 12297 50892 12307 50948
rect 12363 50892 12431 50948
rect 12487 50892 12497 50948
rect 12297 50824 12497 50892
rect 12297 50768 12307 50824
rect 12363 50768 12431 50824
rect 12487 50768 12497 50824
rect 12297 50700 12497 50768
rect 12297 50644 12307 50700
rect 12363 50644 12431 50700
rect 12487 50644 12497 50700
rect 12297 50576 12497 50644
rect 12297 50520 12307 50576
rect 12363 50520 12431 50576
rect 12487 50520 12497 50576
rect 12297 50452 12497 50520
rect 12297 50396 12307 50452
rect 12363 50396 12431 50452
rect 12487 50396 12497 50452
rect 12297 50328 12497 50396
rect 12297 50272 12307 50328
rect 12363 50272 12431 50328
rect 12487 50272 12497 50328
rect 12297 50204 12497 50272
rect 12297 50148 12307 50204
rect 12363 50148 12431 50204
rect 12487 50148 12497 50204
rect 12297 50080 12497 50148
rect 12297 50024 12307 50080
rect 12363 50024 12431 50080
rect 12487 50024 12497 50080
rect 12297 49956 12497 50024
rect 12297 49900 12307 49956
rect 12363 49900 12431 49956
rect 12487 49900 12497 49956
rect 12297 49832 12497 49900
rect 12297 49776 12307 49832
rect 12363 49776 12431 49832
rect 12487 49776 12497 49832
rect 12297 49708 12497 49776
rect 12297 49652 12307 49708
rect 12363 49652 12431 49708
rect 12487 49652 12497 49708
rect 12297 49642 12497 49652
rect 305 48042 2117 49358
rect 2798 48042 4734 49358
rect 5168 48042 7104 49358
rect 7874 48042 9810 49358
rect 10244 48042 12180 49358
rect 12861 48042 14673 49358
rect 2481 46442 2681 47758
rect 4851 46442 5051 47758
rect 7265 46442 7713 47758
rect 9927 46442 10127 47758
rect 12297 46442 12497 47758
rect 305 44842 2117 46158
rect 2798 44842 4734 46158
rect 5168 44842 7104 46158
rect 7874 44842 9810 46158
rect 10244 44842 12180 46158
rect 12861 44842 14673 46158
rect 2481 43242 2681 44558
rect 4851 43242 5051 44558
rect 7265 43242 7713 44558
rect 9927 43242 10127 44558
rect 12297 43242 12497 44558
rect 2481 41642 2681 42958
rect 4851 41642 5051 42958
rect 7265 41642 7713 42958
rect 9927 41642 10127 42958
rect 12297 41642 12497 42958
rect 2481 40042 2681 41358
rect 4851 40042 5051 41358
rect 7265 40042 7713 41358
rect 9927 40042 10127 41358
rect 12297 40042 12497 41358
rect 2481 39748 2681 39758
rect 2292 39727 2368 39737
rect 2292 39671 2302 39727
rect 2358 39671 2368 39727
rect 2292 39595 2368 39671
rect 2292 39539 2302 39595
rect 2358 39539 2368 39595
rect 2292 39463 2368 39539
rect 2292 39407 2302 39463
rect 2358 39407 2368 39463
rect 2292 39331 2368 39407
rect 2292 39275 2302 39331
rect 2358 39275 2368 39331
rect 2292 39199 2368 39275
rect 2292 39143 2302 39199
rect 2358 39143 2368 39199
rect 2292 39067 2368 39143
rect 2292 39011 2302 39067
rect 2358 39011 2368 39067
rect 2292 38935 2368 39011
rect 2292 38879 2302 38935
rect 2358 38879 2368 38935
rect 2292 38803 2368 38879
rect 2292 38747 2302 38803
rect 2358 38747 2368 38803
rect 2292 38671 2368 38747
rect 2292 38615 2302 38671
rect 2358 38615 2368 38671
rect 2292 38539 2368 38615
rect 2292 38483 2302 38539
rect 2358 38483 2368 38539
rect 2292 38473 2368 38483
rect 2481 39692 2491 39748
rect 2547 39692 2615 39748
rect 2671 39692 2681 39748
rect 2481 39624 2681 39692
rect 2481 39568 2491 39624
rect 2547 39568 2615 39624
rect 2671 39568 2681 39624
rect 2481 39500 2681 39568
rect 2481 39444 2491 39500
rect 2547 39444 2615 39500
rect 2671 39444 2681 39500
rect 2481 39376 2681 39444
rect 2481 39320 2491 39376
rect 2547 39320 2615 39376
rect 2671 39320 2681 39376
rect 2481 39252 2681 39320
rect 2481 39196 2491 39252
rect 2547 39196 2615 39252
rect 2671 39196 2681 39252
rect 2481 39128 2681 39196
rect 2481 39072 2491 39128
rect 2547 39072 2615 39128
rect 2671 39072 2681 39128
rect 2481 39004 2681 39072
rect 2481 38948 2491 39004
rect 2547 38948 2615 39004
rect 2671 38948 2681 39004
rect 2481 38880 2681 38948
rect 2481 38824 2491 38880
rect 2547 38824 2615 38880
rect 2671 38824 2681 38880
rect 2481 38756 2681 38824
rect 2481 38700 2491 38756
rect 2547 38700 2615 38756
rect 2671 38700 2681 38756
rect 2481 38632 2681 38700
rect 2481 38576 2491 38632
rect 2547 38576 2615 38632
rect 2671 38576 2681 38632
rect 2481 38508 2681 38576
rect 2481 38452 2491 38508
rect 2547 38452 2615 38508
rect 2671 38452 2681 38508
rect 2481 38442 2681 38452
rect 4851 39748 5051 39758
rect 4851 39692 4861 39748
rect 4917 39692 4985 39748
rect 5041 39692 5051 39748
rect 4851 39624 5051 39692
rect 4851 39568 4861 39624
rect 4917 39568 4985 39624
rect 5041 39568 5051 39624
rect 4851 39500 5051 39568
rect 4851 39444 4861 39500
rect 4917 39444 4985 39500
rect 5041 39444 5051 39500
rect 4851 39376 5051 39444
rect 4851 39320 4861 39376
rect 4917 39320 4985 39376
rect 5041 39320 5051 39376
rect 4851 39252 5051 39320
rect 4851 39196 4861 39252
rect 4917 39196 4985 39252
rect 5041 39196 5051 39252
rect 4851 39128 5051 39196
rect 4851 39072 4861 39128
rect 4917 39072 4985 39128
rect 5041 39072 5051 39128
rect 4851 39004 5051 39072
rect 4851 38948 4861 39004
rect 4917 38948 4985 39004
rect 5041 38948 5051 39004
rect 4851 38880 5051 38948
rect 4851 38824 4861 38880
rect 4917 38824 4985 38880
rect 5041 38824 5051 38880
rect 4851 38756 5051 38824
rect 4851 38700 4861 38756
rect 4917 38700 4985 38756
rect 5041 38700 5051 38756
rect 4851 38632 5051 38700
rect 4851 38576 4861 38632
rect 4917 38576 4985 38632
rect 5041 38576 5051 38632
rect 4851 38508 5051 38576
rect 4851 38452 4861 38508
rect 4917 38452 4985 38508
rect 5041 38452 5051 38508
rect 4851 38442 5051 38452
rect 7265 39748 7713 39758
rect 7265 39692 7275 39748
rect 7331 39692 7399 39748
rect 7455 39692 7523 39748
rect 7579 39692 7647 39748
rect 7703 39692 7713 39748
rect 7265 39624 7713 39692
rect 7265 39568 7275 39624
rect 7331 39568 7399 39624
rect 7455 39568 7523 39624
rect 7579 39568 7647 39624
rect 7703 39568 7713 39624
rect 7265 39500 7713 39568
rect 7265 39444 7275 39500
rect 7331 39444 7399 39500
rect 7455 39444 7523 39500
rect 7579 39444 7647 39500
rect 7703 39444 7713 39500
rect 7265 39376 7713 39444
rect 7265 39320 7275 39376
rect 7331 39320 7399 39376
rect 7455 39320 7523 39376
rect 7579 39320 7647 39376
rect 7703 39320 7713 39376
rect 7265 39252 7713 39320
rect 7265 39196 7275 39252
rect 7331 39196 7399 39252
rect 7455 39196 7523 39252
rect 7579 39196 7647 39252
rect 7703 39196 7713 39252
rect 7265 39128 7713 39196
rect 7265 39072 7275 39128
rect 7331 39072 7399 39128
rect 7455 39072 7523 39128
rect 7579 39072 7647 39128
rect 7703 39072 7713 39128
rect 7265 39004 7713 39072
rect 7265 38948 7275 39004
rect 7331 38948 7399 39004
rect 7455 38948 7523 39004
rect 7579 38948 7647 39004
rect 7703 38948 7713 39004
rect 7265 38880 7713 38948
rect 7265 38824 7275 38880
rect 7331 38824 7399 38880
rect 7455 38824 7523 38880
rect 7579 38824 7647 38880
rect 7703 38824 7713 38880
rect 7265 38756 7713 38824
rect 7265 38700 7275 38756
rect 7331 38700 7399 38756
rect 7455 38700 7523 38756
rect 7579 38700 7647 38756
rect 7703 38700 7713 38756
rect 7265 38632 7713 38700
rect 7265 38576 7275 38632
rect 7331 38576 7399 38632
rect 7455 38576 7523 38632
rect 7579 38576 7647 38632
rect 7703 38576 7713 38632
rect 7265 38508 7713 38576
rect 7265 38452 7275 38508
rect 7331 38452 7399 38508
rect 7455 38452 7523 38508
rect 7579 38452 7647 38508
rect 7703 38452 7713 38508
rect 7265 38442 7713 38452
rect 9927 39748 10127 39758
rect 9927 39692 9937 39748
rect 9993 39692 10061 39748
rect 10117 39692 10127 39748
rect 9927 39624 10127 39692
rect 9927 39568 9937 39624
rect 9993 39568 10061 39624
rect 10117 39568 10127 39624
rect 9927 39500 10127 39568
rect 9927 39444 9937 39500
rect 9993 39444 10061 39500
rect 10117 39444 10127 39500
rect 9927 39376 10127 39444
rect 9927 39320 9937 39376
rect 9993 39320 10061 39376
rect 10117 39320 10127 39376
rect 9927 39252 10127 39320
rect 9927 39196 9937 39252
rect 9993 39196 10061 39252
rect 10117 39196 10127 39252
rect 9927 39128 10127 39196
rect 9927 39072 9937 39128
rect 9993 39072 10061 39128
rect 10117 39072 10127 39128
rect 9927 39004 10127 39072
rect 9927 38948 9937 39004
rect 9993 38948 10061 39004
rect 10117 38948 10127 39004
rect 9927 38880 10127 38948
rect 9927 38824 9937 38880
rect 9993 38824 10061 38880
rect 10117 38824 10127 38880
rect 9927 38756 10127 38824
rect 9927 38700 9937 38756
rect 9993 38700 10061 38756
rect 10117 38700 10127 38756
rect 9927 38632 10127 38700
rect 9927 38576 9937 38632
rect 9993 38576 10061 38632
rect 10117 38576 10127 38632
rect 9927 38508 10127 38576
rect 9927 38452 9937 38508
rect 9993 38452 10061 38508
rect 10117 38452 10127 38508
rect 9927 38442 10127 38452
rect 12297 39748 12497 39758
rect 12297 39692 12307 39748
rect 12363 39692 12431 39748
rect 12487 39692 12497 39748
rect 12297 39624 12497 39692
rect 12297 39568 12307 39624
rect 12363 39568 12431 39624
rect 12487 39568 12497 39624
rect 12297 39500 12497 39568
rect 12297 39444 12307 39500
rect 12363 39444 12431 39500
rect 12487 39444 12497 39500
rect 12297 39376 12497 39444
rect 12297 39320 12307 39376
rect 12363 39320 12431 39376
rect 12487 39320 12497 39376
rect 12297 39252 12497 39320
rect 12297 39196 12307 39252
rect 12363 39196 12431 39252
rect 12487 39196 12497 39252
rect 12297 39128 12497 39196
rect 12297 39072 12307 39128
rect 12363 39072 12431 39128
rect 12487 39072 12497 39128
rect 12297 39004 12497 39072
rect 12297 38948 12307 39004
rect 12363 38948 12431 39004
rect 12487 38948 12497 39004
rect 12297 38880 12497 38948
rect 12297 38824 12307 38880
rect 12363 38824 12431 38880
rect 12487 38824 12497 38880
rect 12297 38756 12497 38824
rect 12297 38700 12307 38756
rect 12363 38700 12431 38756
rect 12487 38700 12497 38756
rect 12297 38632 12497 38700
rect 12297 38576 12307 38632
rect 12363 38576 12431 38632
rect 12487 38576 12497 38632
rect 12297 38508 12497 38576
rect 12297 38452 12307 38508
rect 12363 38452 12431 38508
rect 12487 38452 12497 38508
rect 12297 38442 12497 38452
rect 10 38180 86 38186
rect 14892 38180 14968 38186
rect 10 38176 14968 38180
rect 10 36824 20 38176
rect 76 38148 14902 38176
rect 76 38092 315 38148
rect 371 38092 439 38148
rect 495 38092 563 38148
rect 619 38092 687 38148
rect 743 38092 811 38148
rect 867 38092 935 38148
rect 991 38092 1059 38148
rect 1115 38092 1183 38148
rect 1239 38092 1307 38148
rect 1363 38092 1431 38148
rect 1487 38092 1555 38148
rect 1611 38092 1679 38148
rect 1735 38092 1803 38148
rect 1859 38092 1927 38148
rect 1983 38092 2051 38148
rect 2107 38092 2808 38148
rect 2864 38092 2932 38148
rect 2988 38092 3056 38148
rect 3112 38092 3180 38148
rect 3236 38092 3304 38148
rect 3360 38092 3428 38148
rect 3484 38092 3552 38148
rect 3608 38092 3676 38148
rect 3732 38092 3800 38148
rect 3856 38092 3924 38148
rect 3980 38092 4048 38148
rect 4104 38092 4172 38148
rect 4228 38092 4296 38148
rect 4352 38092 4420 38148
rect 4476 38092 4544 38148
rect 4600 38092 4668 38148
rect 4724 38092 5178 38148
rect 5234 38092 5302 38148
rect 5358 38092 5426 38148
rect 5482 38092 5550 38148
rect 5606 38092 5674 38148
rect 5730 38092 5798 38148
rect 5854 38092 5922 38148
rect 5978 38092 6046 38148
rect 6102 38092 6170 38148
rect 6226 38092 6294 38148
rect 6350 38092 6418 38148
rect 6474 38092 6542 38148
rect 6598 38092 6666 38148
rect 6722 38092 6790 38148
rect 6846 38092 6914 38148
rect 6970 38092 7038 38148
rect 7094 38092 7884 38148
rect 7940 38092 8008 38148
rect 8064 38092 8132 38148
rect 8188 38092 8256 38148
rect 8312 38092 8380 38148
rect 8436 38092 8504 38148
rect 8560 38092 8628 38148
rect 8684 38092 8752 38148
rect 8808 38092 8876 38148
rect 8932 38092 9000 38148
rect 9056 38092 9124 38148
rect 9180 38092 9248 38148
rect 9304 38092 9372 38148
rect 9428 38092 9496 38148
rect 9552 38092 9620 38148
rect 9676 38092 9744 38148
rect 9800 38092 10254 38148
rect 10310 38092 10378 38148
rect 10434 38092 10502 38148
rect 10558 38092 10626 38148
rect 10682 38092 10750 38148
rect 10806 38092 10874 38148
rect 10930 38092 10998 38148
rect 11054 38092 11122 38148
rect 11178 38092 11246 38148
rect 11302 38092 11370 38148
rect 11426 38092 11494 38148
rect 11550 38092 11618 38148
rect 11674 38092 11742 38148
rect 11798 38092 11866 38148
rect 11922 38092 11990 38148
rect 12046 38092 12114 38148
rect 12170 38092 12871 38148
rect 12927 38092 12995 38148
rect 13051 38092 13119 38148
rect 13175 38092 13243 38148
rect 13299 38092 13367 38148
rect 13423 38092 13491 38148
rect 13547 38092 13615 38148
rect 13671 38092 13739 38148
rect 13795 38092 13863 38148
rect 13919 38092 13987 38148
rect 14043 38092 14111 38148
rect 14167 38092 14235 38148
rect 14291 38092 14359 38148
rect 14415 38092 14483 38148
rect 14539 38092 14607 38148
rect 14663 38092 14902 38148
rect 76 38024 14902 38092
rect 76 37968 315 38024
rect 371 37968 439 38024
rect 495 37968 563 38024
rect 619 37968 687 38024
rect 743 37968 811 38024
rect 867 37968 935 38024
rect 991 37968 1059 38024
rect 1115 37968 1183 38024
rect 1239 37968 1307 38024
rect 1363 37968 1431 38024
rect 1487 37968 1555 38024
rect 1611 37968 1679 38024
rect 1735 37968 1803 38024
rect 1859 37968 1927 38024
rect 1983 37968 2051 38024
rect 2107 37968 2808 38024
rect 2864 37968 2932 38024
rect 2988 37968 3056 38024
rect 3112 37968 3180 38024
rect 3236 37968 3304 38024
rect 3360 37968 3428 38024
rect 3484 37968 3552 38024
rect 3608 37968 3676 38024
rect 3732 37968 3800 38024
rect 3856 37968 3924 38024
rect 3980 37968 4048 38024
rect 4104 37968 4172 38024
rect 4228 37968 4296 38024
rect 4352 37968 4420 38024
rect 4476 37968 4544 38024
rect 4600 37968 4668 38024
rect 4724 37968 5178 38024
rect 5234 37968 5302 38024
rect 5358 37968 5426 38024
rect 5482 37968 5550 38024
rect 5606 37968 5674 38024
rect 5730 37968 5798 38024
rect 5854 37968 5922 38024
rect 5978 37968 6046 38024
rect 6102 37968 6170 38024
rect 6226 37968 6294 38024
rect 6350 37968 6418 38024
rect 6474 37968 6542 38024
rect 6598 37968 6666 38024
rect 6722 37968 6790 38024
rect 6846 37968 6914 38024
rect 6970 37968 7038 38024
rect 7094 37968 7884 38024
rect 7940 37968 8008 38024
rect 8064 37968 8132 38024
rect 8188 37968 8256 38024
rect 8312 37968 8380 38024
rect 8436 37968 8504 38024
rect 8560 37968 8628 38024
rect 8684 37968 8752 38024
rect 8808 37968 8876 38024
rect 8932 37968 9000 38024
rect 9056 37968 9124 38024
rect 9180 37968 9248 38024
rect 9304 37968 9372 38024
rect 9428 37968 9496 38024
rect 9552 37968 9620 38024
rect 9676 37968 9744 38024
rect 9800 37968 10254 38024
rect 10310 37968 10378 38024
rect 10434 37968 10502 38024
rect 10558 37968 10626 38024
rect 10682 37968 10750 38024
rect 10806 37968 10874 38024
rect 10930 37968 10998 38024
rect 11054 37968 11122 38024
rect 11178 37968 11246 38024
rect 11302 37968 11370 38024
rect 11426 37968 11494 38024
rect 11550 37968 11618 38024
rect 11674 37968 11742 38024
rect 11798 37968 11866 38024
rect 11922 37968 11990 38024
rect 12046 37968 12114 38024
rect 12170 37968 12871 38024
rect 12927 37968 12995 38024
rect 13051 37968 13119 38024
rect 13175 37968 13243 38024
rect 13299 37968 13367 38024
rect 13423 37968 13491 38024
rect 13547 37968 13615 38024
rect 13671 37968 13739 38024
rect 13795 37968 13863 38024
rect 13919 37968 13987 38024
rect 14043 37968 14111 38024
rect 14167 37968 14235 38024
rect 14291 37968 14359 38024
rect 14415 37968 14483 38024
rect 14539 37968 14607 38024
rect 14663 37968 14902 38024
rect 76 37900 14902 37968
rect 76 37844 315 37900
rect 371 37844 439 37900
rect 495 37844 563 37900
rect 619 37844 687 37900
rect 743 37844 811 37900
rect 867 37844 935 37900
rect 991 37844 1059 37900
rect 1115 37844 1183 37900
rect 1239 37844 1307 37900
rect 1363 37844 1431 37900
rect 1487 37844 1555 37900
rect 1611 37844 1679 37900
rect 1735 37844 1803 37900
rect 1859 37844 1927 37900
rect 1983 37844 2051 37900
rect 2107 37844 2808 37900
rect 2864 37844 2932 37900
rect 2988 37844 3056 37900
rect 3112 37844 3180 37900
rect 3236 37844 3304 37900
rect 3360 37844 3428 37900
rect 3484 37844 3552 37900
rect 3608 37844 3676 37900
rect 3732 37844 3800 37900
rect 3856 37844 3924 37900
rect 3980 37844 4048 37900
rect 4104 37844 4172 37900
rect 4228 37844 4296 37900
rect 4352 37844 4420 37900
rect 4476 37844 4544 37900
rect 4600 37844 4668 37900
rect 4724 37844 5178 37900
rect 5234 37844 5302 37900
rect 5358 37844 5426 37900
rect 5482 37844 5550 37900
rect 5606 37844 5674 37900
rect 5730 37844 5798 37900
rect 5854 37844 5922 37900
rect 5978 37844 6046 37900
rect 6102 37844 6170 37900
rect 6226 37844 6294 37900
rect 6350 37844 6418 37900
rect 6474 37844 6542 37900
rect 6598 37844 6666 37900
rect 6722 37844 6790 37900
rect 6846 37844 6914 37900
rect 6970 37844 7038 37900
rect 7094 37844 7884 37900
rect 7940 37844 8008 37900
rect 8064 37844 8132 37900
rect 8188 37844 8256 37900
rect 8312 37844 8380 37900
rect 8436 37844 8504 37900
rect 8560 37844 8628 37900
rect 8684 37844 8752 37900
rect 8808 37844 8876 37900
rect 8932 37844 9000 37900
rect 9056 37844 9124 37900
rect 9180 37844 9248 37900
rect 9304 37844 9372 37900
rect 9428 37844 9496 37900
rect 9552 37844 9620 37900
rect 9676 37844 9744 37900
rect 9800 37844 10254 37900
rect 10310 37844 10378 37900
rect 10434 37844 10502 37900
rect 10558 37844 10626 37900
rect 10682 37844 10750 37900
rect 10806 37844 10874 37900
rect 10930 37844 10998 37900
rect 11054 37844 11122 37900
rect 11178 37844 11246 37900
rect 11302 37844 11370 37900
rect 11426 37844 11494 37900
rect 11550 37844 11618 37900
rect 11674 37844 11742 37900
rect 11798 37844 11866 37900
rect 11922 37844 11990 37900
rect 12046 37844 12114 37900
rect 12170 37844 12871 37900
rect 12927 37844 12995 37900
rect 13051 37844 13119 37900
rect 13175 37844 13243 37900
rect 13299 37844 13367 37900
rect 13423 37844 13491 37900
rect 13547 37844 13615 37900
rect 13671 37844 13739 37900
rect 13795 37844 13863 37900
rect 13919 37844 13987 37900
rect 14043 37844 14111 37900
rect 14167 37844 14235 37900
rect 14291 37844 14359 37900
rect 14415 37844 14483 37900
rect 14539 37844 14607 37900
rect 14663 37844 14902 37900
rect 76 37776 14902 37844
rect 76 37720 315 37776
rect 371 37720 439 37776
rect 495 37720 563 37776
rect 619 37720 687 37776
rect 743 37720 811 37776
rect 867 37720 935 37776
rect 991 37720 1059 37776
rect 1115 37720 1183 37776
rect 1239 37720 1307 37776
rect 1363 37720 1431 37776
rect 1487 37720 1555 37776
rect 1611 37720 1679 37776
rect 1735 37720 1803 37776
rect 1859 37720 1927 37776
rect 1983 37720 2051 37776
rect 2107 37720 2808 37776
rect 2864 37720 2932 37776
rect 2988 37720 3056 37776
rect 3112 37720 3180 37776
rect 3236 37720 3304 37776
rect 3360 37720 3428 37776
rect 3484 37720 3552 37776
rect 3608 37720 3676 37776
rect 3732 37720 3800 37776
rect 3856 37720 3924 37776
rect 3980 37720 4048 37776
rect 4104 37720 4172 37776
rect 4228 37720 4296 37776
rect 4352 37720 4420 37776
rect 4476 37720 4544 37776
rect 4600 37720 4668 37776
rect 4724 37720 5178 37776
rect 5234 37720 5302 37776
rect 5358 37720 5426 37776
rect 5482 37720 5550 37776
rect 5606 37720 5674 37776
rect 5730 37720 5798 37776
rect 5854 37720 5922 37776
rect 5978 37720 6046 37776
rect 6102 37720 6170 37776
rect 6226 37720 6294 37776
rect 6350 37720 6418 37776
rect 6474 37720 6542 37776
rect 6598 37720 6666 37776
rect 6722 37720 6790 37776
rect 6846 37720 6914 37776
rect 6970 37720 7038 37776
rect 7094 37720 7884 37776
rect 7940 37720 8008 37776
rect 8064 37720 8132 37776
rect 8188 37720 8256 37776
rect 8312 37720 8380 37776
rect 8436 37720 8504 37776
rect 8560 37720 8628 37776
rect 8684 37720 8752 37776
rect 8808 37720 8876 37776
rect 8932 37720 9000 37776
rect 9056 37720 9124 37776
rect 9180 37720 9248 37776
rect 9304 37720 9372 37776
rect 9428 37720 9496 37776
rect 9552 37720 9620 37776
rect 9676 37720 9744 37776
rect 9800 37720 10254 37776
rect 10310 37720 10378 37776
rect 10434 37720 10502 37776
rect 10558 37720 10626 37776
rect 10682 37720 10750 37776
rect 10806 37720 10874 37776
rect 10930 37720 10998 37776
rect 11054 37720 11122 37776
rect 11178 37720 11246 37776
rect 11302 37720 11370 37776
rect 11426 37720 11494 37776
rect 11550 37720 11618 37776
rect 11674 37720 11742 37776
rect 11798 37720 11866 37776
rect 11922 37720 11990 37776
rect 12046 37720 12114 37776
rect 12170 37720 12871 37776
rect 12927 37720 12995 37776
rect 13051 37720 13119 37776
rect 13175 37720 13243 37776
rect 13299 37720 13367 37776
rect 13423 37720 13491 37776
rect 13547 37720 13615 37776
rect 13671 37720 13739 37776
rect 13795 37720 13863 37776
rect 13919 37720 13987 37776
rect 14043 37720 14111 37776
rect 14167 37720 14235 37776
rect 14291 37720 14359 37776
rect 14415 37720 14483 37776
rect 14539 37720 14607 37776
rect 14663 37720 14902 37776
rect 76 37652 14902 37720
rect 76 37596 315 37652
rect 371 37596 439 37652
rect 495 37596 563 37652
rect 619 37596 687 37652
rect 743 37596 811 37652
rect 867 37596 935 37652
rect 991 37596 1059 37652
rect 1115 37596 1183 37652
rect 1239 37596 1307 37652
rect 1363 37596 1431 37652
rect 1487 37596 1555 37652
rect 1611 37596 1679 37652
rect 1735 37596 1803 37652
rect 1859 37596 1927 37652
rect 1983 37596 2051 37652
rect 2107 37596 2808 37652
rect 2864 37596 2932 37652
rect 2988 37596 3056 37652
rect 3112 37596 3180 37652
rect 3236 37596 3304 37652
rect 3360 37596 3428 37652
rect 3484 37596 3552 37652
rect 3608 37596 3676 37652
rect 3732 37596 3800 37652
rect 3856 37596 3924 37652
rect 3980 37596 4048 37652
rect 4104 37596 4172 37652
rect 4228 37596 4296 37652
rect 4352 37596 4420 37652
rect 4476 37596 4544 37652
rect 4600 37596 4668 37652
rect 4724 37596 5178 37652
rect 5234 37596 5302 37652
rect 5358 37596 5426 37652
rect 5482 37596 5550 37652
rect 5606 37596 5674 37652
rect 5730 37596 5798 37652
rect 5854 37596 5922 37652
rect 5978 37596 6046 37652
rect 6102 37596 6170 37652
rect 6226 37596 6294 37652
rect 6350 37596 6418 37652
rect 6474 37596 6542 37652
rect 6598 37596 6666 37652
rect 6722 37596 6790 37652
rect 6846 37596 6914 37652
rect 6970 37596 7038 37652
rect 7094 37596 7884 37652
rect 7940 37596 8008 37652
rect 8064 37596 8132 37652
rect 8188 37596 8256 37652
rect 8312 37596 8380 37652
rect 8436 37596 8504 37652
rect 8560 37596 8628 37652
rect 8684 37596 8752 37652
rect 8808 37596 8876 37652
rect 8932 37596 9000 37652
rect 9056 37596 9124 37652
rect 9180 37596 9248 37652
rect 9304 37596 9372 37652
rect 9428 37596 9496 37652
rect 9552 37596 9620 37652
rect 9676 37596 9744 37652
rect 9800 37596 10254 37652
rect 10310 37596 10378 37652
rect 10434 37596 10502 37652
rect 10558 37596 10626 37652
rect 10682 37596 10750 37652
rect 10806 37596 10874 37652
rect 10930 37596 10998 37652
rect 11054 37596 11122 37652
rect 11178 37596 11246 37652
rect 11302 37596 11370 37652
rect 11426 37596 11494 37652
rect 11550 37596 11618 37652
rect 11674 37596 11742 37652
rect 11798 37596 11866 37652
rect 11922 37596 11990 37652
rect 12046 37596 12114 37652
rect 12170 37596 12871 37652
rect 12927 37596 12995 37652
rect 13051 37596 13119 37652
rect 13175 37596 13243 37652
rect 13299 37596 13367 37652
rect 13423 37596 13491 37652
rect 13547 37596 13615 37652
rect 13671 37596 13739 37652
rect 13795 37596 13863 37652
rect 13919 37596 13987 37652
rect 14043 37596 14111 37652
rect 14167 37596 14235 37652
rect 14291 37596 14359 37652
rect 14415 37596 14483 37652
rect 14539 37596 14607 37652
rect 14663 37596 14902 37652
rect 76 37528 14902 37596
rect 76 37472 315 37528
rect 371 37472 439 37528
rect 495 37472 563 37528
rect 619 37472 687 37528
rect 743 37472 811 37528
rect 867 37472 935 37528
rect 991 37472 1059 37528
rect 1115 37472 1183 37528
rect 1239 37472 1307 37528
rect 1363 37472 1431 37528
rect 1487 37472 1555 37528
rect 1611 37472 1679 37528
rect 1735 37472 1803 37528
rect 1859 37472 1927 37528
rect 1983 37472 2051 37528
rect 2107 37472 2808 37528
rect 2864 37472 2932 37528
rect 2988 37472 3056 37528
rect 3112 37472 3180 37528
rect 3236 37472 3304 37528
rect 3360 37472 3428 37528
rect 3484 37472 3552 37528
rect 3608 37472 3676 37528
rect 3732 37472 3800 37528
rect 3856 37472 3924 37528
rect 3980 37472 4048 37528
rect 4104 37472 4172 37528
rect 4228 37472 4296 37528
rect 4352 37472 4420 37528
rect 4476 37472 4544 37528
rect 4600 37472 4668 37528
rect 4724 37472 5178 37528
rect 5234 37472 5302 37528
rect 5358 37472 5426 37528
rect 5482 37472 5550 37528
rect 5606 37472 5674 37528
rect 5730 37472 5798 37528
rect 5854 37472 5922 37528
rect 5978 37472 6046 37528
rect 6102 37472 6170 37528
rect 6226 37472 6294 37528
rect 6350 37472 6418 37528
rect 6474 37472 6542 37528
rect 6598 37472 6666 37528
rect 6722 37472 6790 37528
rect 6846 37472 6914 37528
rect 6970 37472 7038 37528
rect 7094 37472 7884 37528
rect 7940 37472 8008 37528
rect 8064 37472 8132 37528
rect 8188 37472 8256 37528
rect 8312 37472 8380 37528
rect 8436 37472 8504 37528
rect 8560 37472 8628 37528
rect 8684 37472 8752 37528
rect 8808 37472 8876 37528
rect 8932 37472 9000 37528
rect 9056 37472 9124 37528
rect 9180 37472 9248 37528
rect 9304 37472 9372 37528
rect 9428 37472 9496 37528
rect 9552 37472 9620 37528
rect 9676 37472 9744 37528
rect 9800 37472 10254 37528
rect 10310 37472 10378 37528
rect 10434 37472 10502 37528
rect 10558 37472 10626 37528
rect 10682 37472 10750 37528
rect 10806 37472 10874 37528
rect 10930 37472 10998 37528
rect 11054 37472 11122 37528
rect 11178 37472 11246 37528
rect 11302 37472 11370 37528
rect 11426 37472 11494 37528
rect 11550 37472 11618 37528
rect 11674 37472 11742 37528
rect 11798 37472 11866 37528
rect 11922 37472 11990 37528
rect 12046 37472 12114 37528
rect 12170 37472 12871 37528
rect 12927 37472 12995 37528
rect 13051 37472 13119 37528
rect 13175 37472 13243 37528
rect 13299 37472 13367 37528
rect 13423 37472 13491 37528
rect 13547 37472 13615 37528
rect 13671 37472 13739 37528
rect 13795 37472 13863 37528
rect 13919 37472 13987 37528
rect 14043 37472 14111 37528
rect 14167 37472 14235 37528
rect 14291 37472 14359 37528
rect 14415 37472 14483 37528
rect 14539 37472 14607 37528
rect 14663 37472 14902 37528
rect 76 37404 14902 37472
rect 76 37348 315 37404
rect 371 37348 439 37404
rect 495 37348 563 37404
rect 619 37348 687 37404
rect 743 37348 811 37404
rect 867 37348 935 37404
rect 991 37348 1059 37404
rect 1115 37348 1183 37404
rect 1239 37348 1307 37404
rect 1363 37348 1431 37404
rect 1487 37348 1555 37404
rect 1611 37348 1679 37404
rect 1735 37348 1803 37404
rect 1859 37348 1927 37404
rect 1983 37348 2051 37404
rect 2107 37348 2808 37404
rect 2864 37348 2932 37404
rect 2988 37348 3056 37404
rect 3112 37348 3180 37404
rect 3236 37348 3304 37404
rect 3360 37348 3428 37404
rect 3484 37348 3552 37404
rect 3608 37348 3676 37404
rect 3732 37348 3800 37404
rect 3856 37348 3924 37404
rect 3980 37348 4048 37404
rect 4104 37348 4172 37404
rect 4228 37348 4296 37404
rect 4352 37348 4420 37404
rect 4476 37348 4544 37404
rect 4600 37348 4668 37404
rect 4724 37348 5178 37404
rect 5234 37348 5302 37404
rect 5358 37348 5426 37404
rect 5482 37348 5550 37404
rect 5606 37348 5674 37404
rect 5730 37348 5798 37404
rect 5854 37348 5922 37404
rect 5978 37348 6046 37404
rect 6102 37348 6170 37404
rect 6226 37348 6294 37404
rect 6350 37348 6418 37404
rect 6474 37348 6542 37404
rect 6598 37348 6666 37404
rect 6722 37348 6790 37404
rect 6846 37348 6914 37404
rect 6970 37348 7038 37404
rect 7094 37348 7884 37404
rect 7940 37348 8008 37404
rect 8064 37348 8132 37404
rect 8188 37348 8256 37404
rect 8312 37348 8380 37404
rect 8436 37348 8504 37404
rect 8560 37348 8628 37404
rect 8684 37348 8752 37404
rect 8808 37348 8876 37404
rect 8932 37348 9000 37404
rect 9056 37348 9124 37404
rect 9180 37348 9248 37404
rect 9304 37348 9372 37404
rect 9428 37348 9496 37404
rect 9552 37348 9620 37404
rect 9676 37348 9744 37404
rect 9800 37348 10254 37404
rect 10310 37348 10378 37404
rect 10434 37348 10502 37404
rect 10558 37348 10626 37404
rect 10682 37348 10750 37404
rect 10806 37348 10874 37404
rect 10930 37348 10998 37404
rect 11054 37348 11122 37404
rect 11178 37348 11246 37404
rect 11302 37348 11370 37404
rect 11426 37348 11494 37404
rect 11550 37348 11618 37404
rect 11674 37348 11742 37404
rect 11798 37348 11866 37404
rect 11922 37348 11990 37404
rect 12046 37348 12114 37404
rect 12170 37348 12871 37404
rect 12927 37348 12995 37404
rect 13051 37348 13119 37404
rect 13175 37348 13243 37404
rect 13299 37348 13367 37404
rect 13423 37348 13491 37404
rect 13547 37348 13615 37404
rect 13671 37348 13739 37404
rect 13795 37348 13863 37404
rect 13919 37348 13987 37404
rect 14043 37348 14111 37404
rect 14167 37348 14235 37404
rect 14291 37348 14359 37404
rect 14415 37348 14483 37404
rect 14539 37348 14607 37404
rect 14663 37348 14902 37404
rect 76 37280 14902 37348
rect 76 37224 315 37280
rect 371 37224 439 37280
rect 495 37224 563 37280
rect 619 37224 687 37280
rect 743 37224 811 37280
rect 867 37224 935 37280
rect 991 37224 1059 37280
rect 1115 37224 1183 37280
rect 1239 37224 1307 37280
rect 1363 37224 1431 37280
rect 1487 37224 1555 37280
rect 1611 37224 1679 37280
rect 1735 37224 1803 37280
rect 1859 37224 1927 37280
rect 1983 37224 2051 37280
rect 2107 37224 2808 37280
rect 2864 37224 2932 37280
rect 2988 37224 3056 37280
rect 3112 37224 3180 37280
rect 3236 37224 3304 37280
rect 3360 37224 3428 37280
rect 3484 37224 3552 37280
rect 3608 37224 3676 37280
rect 3732 37224 3800 37280
rect 3856 37224 3924 37280
rect 3980 37224 4048 37280
rect 4104 37224 4172 37280
rect 4228 37224 4296 37280
rect 4352 37224 4420 37280
rect 4476 37224 4544 37280
rect 4600 37224 4668 37280
rect 4724 37224 5178 37280
rect 5234 37224 5302 37280
rect 5358 37224 5426 37280
rect 5482 37224 5550 37280
rect 5606 37224 5674 37280
rect 5730 37224 5798 37280
rect 5854 37224 5922 37280
rect 5978 37224 6046 37280
rect 6102 37224 6170 37280
rect 6226 37224 6294 37280
rect 6350 37224 6418 37280
rect 6474 37224 6542 37280
rect 6598 37224 6666 37280
rect 6722 37224 6790 37280
rect 6846 37224 6914 37280
rect 6970 37224 7038 37280
rect 7094 37224 7884 37280
rect 7940 37224 8008 37280
rect 8064 37224 8132 37280
rect 8188 37224 8256 37280
rect 8312 37224 8380 37280
rect 8436 37224 8504 37280
rect 8560 37224 8628 37280
rect 8684 37224 8752 37280
rect 8808 37224 8876 37280
rect 8932 37224 9000 37280
rect 9056 37224 9124 37280
rect 9180 37224 9248 37280
rect 9304 37224 9372 37280
rect 9428 37224 9496 37280
rect 9552 37224 9620 37280
rect 9676 37224 9744 37280
rect 9800 37224 10254 37280
rect 10310 37224 10378 37280
rect 10434 37224 10502 37280
rect 10558 37224 10626 37280
rect 10682 37224 10750 37280
rect 10806 37224 10874 37280
rect 10930 37224 10998 37280
rect 11054 37224 11122 37280
rect 11178 37224 11246 37280
rect 11302 37224 11370 37280
rect 11426 37224 11494 37280
rect 11550 37224 11618 37280
rect 11674 37224 11742 37280
rect 11798 37224 11866 37280
rect 11922 37224 11990 37280
rect 12046 37224 12114 37280
rect 12170 37224 12871 37280
rect 12927 37224 12995 37280
rect 13051 37224 13119 37280
rect 13175 37224 13243 37280
rect 13299 37224 13367 37280
rect 13423 37224 13491 37280
rect 13547 37224 13615 37280
rect 13671 37224 13739 37280
rect 13795 37224 13863 37280
rect 13919 37224 13987 37280
rect 14043 37224 14111 37280
rect 14167 37224 14235 37280
rect 14291 37224 14359 37280
rect 14415 37224 14483 37280
rect 14539 37224 14607 37280
rect 14663 37224 14902 37280
rect 76 37156 14902 37224
rect 76 37100 315 37156
rect 371 37100 439 37156
rect 495 37100 563 37156
rect 619 37100 687 37156
rect 743 37100 811 37156
rect 867 37100 935 37156
rect 991 37100 1059 37156
rect 1115 37100 1183 37156
rect 1239 37100 1307 37156
rect 1363 37100 1431 37156
rect 1487 37100 1555 37156
rect 1611 37100 1679 37156
rect 1735 37100 1803 37156
rect 1859 37100 1927 37156
rect 1983 37100 2051 37156
rect 2107 37100 2808 37156
rect 2864 37100 2932 37156
rect 2988 37100 3056 37156
rect 3112 37100 3180 37156
rect 3236 37100 3304 37156
rect 3360 37100 3428 37156
rect 3484 37100 3552 37156
rect 3608 37100 3676 37156
rect 3732 37100 3800 37156
rect 3856 37100 3924 37156
rect 3980 37100 4048 37156
rect 4104 37100 4172 37156
rect 4228 37100 4296 37156
rect 4352 37100 4420 37156
rect 4476 37100 4544 37156
rect 4600 37100 4668 37156
rect 4724 37100 5178 37156
rect 5234 37100 5302 37156
rect 5358 37100 5426 37156
rect 5482 37100 5550 37156
rect 5606 37100 5674 37156
rect 5730 37100 5798 37156
rect 5854 37100 5922 37156
rect 5978 37100 6046 37156
rect 6102 37100 6170 37156
rect 6226 37100 6294 37156
rect 6350 37100 6418 37156
rect 6474 37100 6542 37156
rect 6598 37100 6666 37156
rect 6722 37100 6790 37156
rect 6846 37100 6914 37156
rect 6970 37100 7038 37156
rect 7094 37100 7884 37156
rect 7940 37100 8008 37156
rect 8064 37100 8132 37156
rect 8188 37100 8256 37156
rect 8312 37100 8380 37156
rect 8436 37100 8504 37156
rect 8560 37100 8628 37156
rect 8684 37100 8752 37156
rect 8808 37100 8876 37156
rect 8932 37100 9000 37156
rect 9056 37100 9124 37156
rect 9180 37100 9248 37156
rect 9304 37100 9372 37156
rect 9428 37100 9496 37156
rect 9552 37100 9620 37156
rect 9676 37100 9744 37156
rect 9800 37100 10254 37156
rect 10310 37100 10378 37156
rect 10434 37100 10502 37156
rect 10558 37100 10626 37156
rect 10682 37100 10750 37156
rect 10806 37100 10874 37156
rect 10930 37100 10998 37156
rect 11054 37100 11122 37156
rect 11178 37100 11246 37156
rect 11302 37100 11370 37156
rect 11426 37100 11494 37156
rect 11550 37100 11618 37156
rect 11674 37100 11742 37156
rect 11798 37100 11866 37156
rect 11922 37100 11990 37156
rect 12046 37100 12114 37156
rect 12170 37100 12871 37156
rect 12927 37100 12995 37156
rect 13051 37100 13119 37156
rect 13175 37100 13243 37156
rect 13299 37100 13367 37156
rect 13423 37100 13491 37156
rect 13547 37100 13615 37156
rect 13671 37100 13739 37156
rect 13795 37100 13863 37156
rect 13919 37100 13987 37156
rect 14043 37100 14111 37156
rect 14167 37100 14235 37156
rect 14291 37100 14359 37156
rect 14415 37100 14483 37156
rect 14539 37100 14607 37156
rect 14663 37100 14902 37156
rect 76 37032 14902 37100
rect 76 36976 315 37032
rect 371 36976 439 37032
rect 495 36976 563 37032
rect 619 36976 687 37032
rect 743 36976 811 37032
rect 867 36976 935 37032
rect 991 36976 1059 37032
rect 1115 36976 1183 37032
rect 1239 36976 1307 37032
rect 1363 36976 1431 37032
rect 1487 36976 1555 37032
rect 1611 36976 1679 37032
rect 1735 36976 1803 37032
rect 1859 36976 1927 37032
rect 1983 36976 2051 37032
rect 2107 36976 2808 37032
rect 2864 36976 2932 37032
rect 2988 36976 3056 37032
rect 3112 36976 3180 37032
rect 3236 36976 3304 37032
rect 3360 36976 3428 37032
rect 3484 36976 3552 37032
rect 3608 36976 3676 37032
rect 3732 36976 3800 37032
rect 3856 36976 3924 37032
rect 3980 36976 4048 37032
rect 4104 36976 4172 37032
rect 4228 36976 4296 37032
rect 4352 36976 4420 37032
rect 4476 36976 4544 37032
rect 4600 36976 4668 37032
rect 4724 36976 5178 37032
rect 5234 36976 5302 37032
rect 5358 36976 5426 37032
rect 5482 36976 5550 37032
rect 5606 36976 5674 37032
rect 5730 36976 5798 37032
rect 5854 36976 5922 37032
rect 5978 36976 6046 37032
rect 6102 36976 6170 37032
rect 6226 36976 6294 37032
rect 6350 36976 6418 37032
rect 6474 36976 6542 37032
rect 6598 36976 6666 37032
rect 6722 36976 6790 37032
rect 6846 36976 6914 37032
rect 6970 36976 7038 37032
rect 7094 36976 7884 37032
rect 7940 36976 8008 37032
rect 8064 36976 8132 37032
rect 8188 36976 8256 37032
rect 8312 36976 8380 37032
rect 8436 36976 8504 37032
rect 8560 36976 8628 37032
rect 8684 36976 8752 37032
rect 8808 36976 8876 37032
rect 8932 36976 9000 37032
rect 9056 36976 9124 37032
rect 9180 36976 9248 37032
rect 9304 36976 9372 37032
rect 9428 36976 9496 37032
rect 9552 36976 9620 37032
rect 9676 36976 9744 37032
rect 9800 36976 10254 37032
rect 10310 36976 10378 37032
rect 10434 36976 10502 37032
rect 10558 36976 10626 37032
rect 10682 36976 10750 37032
rect 10806 36976 10874 37032
rect 10930 36976 10998 37032
rect 11054 36976 11122 37032
rect 11178 36976 11246 37032
rect 11302 36976 11370 37032
rect 11426 36976 11494 37032
rect 11550 36976 11618 37032
rect 11674 36976 11742 37032
rect 11798 36976 11866 37032
rect 11922 36976 11990 37032
rect 12046 36976 12114 37032
rect 12170 36976 12871 37032
rect 12927 36976 12995 37032
rect 13051 36976 13119 37032
rect 13175 36976 13243 37032
rect 13299 36976 13367 37032
rect 13423 36976 13491 37032
rect 13547 36976 13615 37032
rect 13671 36976 13739 37032
rect 13795 36976 13863 37032
rect 13919 36976 13987 37032
rect 14043 36976 14111 37032
rect 14167 36976 14235 37032
rect 14291 36976 14359 37032
rect 14415 36976 14483 37032
rect 14539 36976 14607 37032
rect 14663 36976 14902 37032
rect 76 36908 14902 36976
rect 76 36852 315 36908
rect 371 36852 439 36908
rect 495 36852 563 36908
rect 619 36852 687 36908
rect 743 36852 811 36908
rect 867 36852 935 36908
rect 991 36852 1059 36908
rect 1115 36852 1183 36908
rect 1239 36852 1307 36908
rect 1363 36852 1431 36908
rect 1487 36852 1555 36908
rect 1611 36852 1679 36908
rect 1735 36852 1803 36908
rect 1859 36852 1927 36908
rect 1983 36852 2051 36908
rect 2107 36852 2808 36908
rect 2864 36852 2932 36908
rect 2988 36852 3056 36908
rect 3112 36852 3180 36908
rect 3236 36852 3304 36908
rect 3360 36852 3428 36908
rect 3484 36852 3552 36908
rect 3608 36852 3676 36908
rect 3732 36852 3800 36908
rect 3856 36852 3924 36908
rect 3980 36852 4048 36908
rect 4104 36852 4172 36908
rect 4228 36852 4296 36908
rect 4352 36852 4420 36908
rect 4476 36852 4544 36908
rect 4600 36852 4668 36908
rect 4724 36852 5178 36908
rect 5234 36852 5302 36908
rect 5358 36852 5426 36908
rect 5482 36852 5550 36908
rect 5606 36852 5674 36908
rect 5730 36852 5798 36908
rect 5854 36852 5922 36908
rect 5978 36852 6046 36908
rect 6102 36852 6170 36908
rect 6226 36852 6294 36908
rect 6350 36852 6418 36908
rect 6474 36852 6542 36908
rect 6598 36852 6666 36908
rect 6722 36852 6790 36908
rect 6846 36852 6914 36908
rect 6970 36852 7038 36908
rect 7094 36852 7884 36908
rect 7940 36852 8008 36908
rect 8064 36852 8132 36908
rect 8188 36852 8256 36908
rect 8312 36852 8380 36908
rect 8436 36852 8504 36908
rect 8560 36852 8628 36908
rect 8684 36852 8752 36908
rect 8808 36852 8876 36908
rect 8932 36852 9000 36908
rect 9056 36852 9124 36908
rect 9180 36852 9248 36908
rect 9304 36852 9372 36908
rect 9428 36852 9496 36908
rect 9552 36852 9620 36908
rect 9676 36852 9744 36908
rect 9800 36852 10254 36908
rect 10310 36852 10378 36908
rect 10434 36852 10502 36908
rect 10558 36852 10626 36908
rect 10682 36852 10750 36908
rect 10806 36852 10874 36908
rect 10930 36852 10998 36908
rect 11054 36852 11122 36908
rect 11178 36852 11246 36908
rect 11302 36852 11370 36908
rect 11426 36852 11494 36908
rect 11550 36852 11618 36908
rect 11674 36852 11742 36908
rect 11798 36852 11866 36908
rect 11922 36852 11990 36908
rect 12046 36852 12114 36908
rect 12170 36852 12871 36908
rect 12927 36852 12995 36908
rect 13051 36852 13119 36908
rect 13175 36852 13243 36908
rect 13299 36852 13367 36908
rect 13423 36852 13491 36908
rect 13547 36852 13615 36908
rect 13671 36852 13739 36908
rect 13795 36852 13863 36908
rect 13919 36852 13987 36908
rect 14043 36852 14111 36908
rect 14167 36852 14235 36908
rect 14291 36852 14359 36908
rect 14415 36852 14483 36908
rect 14539 36852 14607 36908
rect 14663 36852 14902 36908
rect 76 36830 14902 36852
rect 76 36824 86 36830
rect 10 36814 86 36824
rect 14892 36824 14902 36830
rect 14958 36824 14968 38176
rect 14892 36814 14968 36824
rect 305 33636 2117 36564
rect 2798 33636 4734 36564
rect 5168 33636 7104 36564
rect 7874 33636 9810 36564
rect 10244 33636 12180 36564
rect 12861 33636 14673 36564
rect 2481 30436 2681 33364
rect 4851 30436 5051 33364
rect 7265 30436 7713 33364
rect 9927 30436 10127 33364
rect 12297 30436 12497 33364
rect 2481 28842 2681 30158
rect 4851 28842 5051 30158
rect 7265 28842 7713 30158
rect 9927 28842 10127 30158
rect 12297 28842 12497 30158
rect 305 27242 2117 28558
rect 2798 27242 4734 28558
rect 5168 27242 7104 28558
rect 7874 27242 9810 28558
rect 10244 27242 12180 28558
rect 12861 27242 14673 28558
rect 2481 24036 2681 26964
rect 4851 24036 5051 26964
rect 7265 24036 7713 26964
rect 9927 24036 10127 26964
rect 12297 24036 12497 26964
rect 2481 20836 2681 23764
rect 4851 20836 5051 23764
rect 7265 20836 7713 23764
rect 9927 20836 10127 23764
rect 12297 20836 12497 23764
rect 2481 17636 2681 20564
rect 4851 17636 5051 20564
rect 7265 17636 7713 20564
rect 9927 17636 10127 20564
rect 12297 17636 12497 20564
rect 2481 14436 2681 17364
rect 4851 14436 5051 17364
rect 7265 14436 7713 17364
rect 9927 14436 10127 17364
rect 12297 14436 12497 17364
rect 305 12842 2117 14158
rect 2798 12842 4734 14158
rect 5168 12842 7104 14158
rect 7874 12842 9810 14158
rect 10244 12842 12180 14158
rect 12861 12842 14673 14158
rect 2481 11242 2681 12558
rect 4851 11242 5051 12558
rect 7265 11242 7713 12558
rect 9927 11242 10127 12558
rect 12297 11242 12497 12558
rect 305 8036 2117 10964
rect 2798 8036 4734 10964
rect 5168 8036 7104 10964
rect 7874 8036 9810 10964
rect 10244 8036 12180 10964
rect 12861 8036 14673 10964
rect 305 4836 2117 7764
rect 2798 4836 4734 7764
rect 5168 4836 7104 7764
rect 7874 4836 9810 7764
rect 10244 4836 12180 7764
rect 12861 4836 14673 7764
rect 305 1636 2117 4564
rect 2798 1636 4734 4564
rect 5168 1636 7104 4564
rect 7874 1636 9810 4564
rect 10244 1636 12180 4564
rect 12861 1636 14673 4564
use comp018green_esd_clamp_v5p0_DVSS  comp018green_esd_clamp_v5p0_DVSS_0
timestamp 1764349902
transform 1 0 1008 0 1 1090
box -747 -51 13709 46134
<< labels >>
rlabel metal3 s 705 6432 705 6432 4 DVSS
port 1 nsew
rlabel metal3 s 752 3261 752 3261 4 DVSS
port 1 nsew
rlabel metal3 s 774 9418 774 9418 4 DVSS
port 1 nsew
rlabel metal3 s 774 13611 774 13611 4 DVSS
port 1 nsew
rlabel metal3 s 774 11795 774 11795 4 DVDD
port 2 nsew
rlabel metal3 s 774 22234 774 22234 4 DVDD
port 2 nsew
rlabel metal3 s 774 19120 774 19120 4 DVDD
port 2 nsew
rlabel metal3 s 774 15905 774 15905 4 DVDD
port 2 nsew
rlabel metal3 s 774 27853 774 27853 4 DVSS
port 1 nsew
rlabel metal3 s 774 29488 774 29488 4 DVDD
port 2 nsew
rlabel metal3 s 774 25470 774 25470 4 DVDD
port 2 nsew
rlabel metal3 s 774 35106 774 35106 4 DVSS
port 1 nsew
rlabel metal3 s 774 31879 774 31879 4 DVDD
port 2 nsew
rlabel metal3 s 774 38969 774 38969 4 VDD
port 3 nsew
rlabel metal3 s 774 45369 774 45369 4 DVSS
port 1 nsew
rlabel metal3 s 774 43934 774 43934 4 DVDD
port 2 nsew
rlabel metal3 s 774 42169 774 42169 4 DVDD
port 2 nsew
rlabel metal3 s 774 40734 774 40734 4 DVDD
port 2 nsew
rlabel metal3 s 774 50334 774 50334 4 VDD
port 3 nsew
rlabel metal3 s 774 48569 774 48569 4 DVSS
port 1 nsew
rlabel metal3 s 774 53534 774 53534 4 DVSS
port 1 nsew
rlabel metal3 s 774 56560 774 56560 4 DVSS
port 1 nsew
rlabel metal3 s 774 54969 774 54969 4 DVDD
port 2 nsew
rlabel metal3 s 774 47134 774 47134 4 DVDD
port 2 nsew
rlabel metal3 s 774 51934 774 51934 4 VSS
port 4 nsew
rlabel metal3 s 774 37534 774 37534 4 VSS
port 4 nsew
<< end >>
