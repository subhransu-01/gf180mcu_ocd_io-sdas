** sch_path: /home/subhransu/gitRepo/gf180mcu_ocd_io-sdas/runs/RUN_2026-01-12_06-34-59/parameters/transient_response/run_3/io_inv_1_tran.sch
**.subckt io_inv_1_tran
x1 VDD Vout Vin VSS io_inv_1
V1 VSS GND 0
V2 VDD GND cace{vdd}
V3 Vin GND 0 PULSE(0 1.8 0 1n 1n 10n 20n)
C1 Vout GND 1p m=1
**** begin user architecture code

.include /home/subhransu/share/pdk/gf180mcuD/libs.tech/ngspice/design.ngspice
.lib /home/subhransu/share/pdk/gf180mcuD/libs.tech/ngspice/sm141064.ngspice typical




*.lib /home/subhransu/share/pdk/gf180mcuD/libs.tech/ngspice/sm141064.ngspice ss
.include /home/subhransu/gitRepo/gf180mcu_ocd_io-sdas/netlist/schematic/io_inv_1.spice
.temp 27
.option SEED=12345
.option warn=1






.control
tran 0.1n 5.0000000000000004e-08
set wr_singlescale
wrdata /home/subhransu/gitRepo/gf180mcu_ocd_io-sdas/runs/RUN_2026-01-12_06-34-59/parameters/transient_response/run_3/io_inv_1_tran_3.data V(Vout) V(Vin)
.endc


**** end user architecture code
**.ends
.GLOBAL GND
.end
