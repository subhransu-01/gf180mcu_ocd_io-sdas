** sch_path: /home/subhransu/gitRepo/gf180mcu_ocd_io-sdas/runs/RUN_2026-01-12_06-25-34/parameters/dc_response/run_1/io_inv_1_dc.sch
**.subckt io_inv_1_dc
V1 VSS GND 0
V2 VDD GND cace{vdd}
V3 Vin GND 1.8
C1 Vout GND 1e-15 m=1
x1 VDD Vout Vin VSS io_inv_1
**** begin user architecture code

.include /home/subhransu/share/pdk/gf180mcuD/libs.tech/ngspice/design.ngspice
.lib /home/subhransu/share/pdk/gf180mcuD/libs.tech/ngspice/sm141064.ngspice typical




*.lib /home/subhransu/share/pdk/gf180mcuD/libs.tech/ngspice/sm141064.ngspice tt
.include /home/subhransu/gitRepo/gf180mcu_ocd_io-sdas/netlist/schematic/io_inv_1.spice
.temp -40
.option SEED=12345
.option warn=1






.control
dc V3 0 1.8 0.01
set wr_singlescale
wrdata /home/subhransu/gitRepo/gf180mcu_ocd_io-sdas/runs/RUN_2026-01-12_06-25-34/parameters/dc_response/run_1/io_inv_1_dc_1.data V(Vin) V(Vout)
.endc


**** end user architecture code
**.ends
.GLOBAL GND
.end
