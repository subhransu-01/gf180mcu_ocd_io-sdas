magic
tech gf180mcuD
magscale 1 10
timestamp 1764347740
<< isosubstrate >>
rect 392 -83 2701 2911
<< nwell >>
rect 1382 2911 2704 2914
rect 392 2575 2704 2911
rect 1382 1242 2704 2575
rect 1385 1213 2701 1242
<< hvnmos >>
rect 1913 270 2053 870
rect 2157 270 2297 870
<< hvpmos >>
rect 1913 1358 2053 2558
rect 2157 1358 2297 2558
<< mvndiff >>
rect 1825 857 1913 870
rect 1825 811 1838 857
rect 1884 811 1913 857
rect 1825 752 1913 811
rect 1825 706 1838 752
rect 1884 706 1913 752
rect 1825 647 1913 706
rect 1825 601 1838 647
rect 1884 601 1913 647
rect 1825 541 1913 601
rect 1825 495 1838 541
rect 1884 495 1913 541
rect 1825 435 1913 495
rect 1825 389 1838 435
rect 1884 389 1913 435
rect 1825 329 1913 389
rect 1825 283 1838 329
rect 1884 283 1913 329
rect 1825 270 1913 283
rect 2053 857 2157 870
rect 2053 811 2082 857
rect 2128 811 2157 857
rect 2053 752 2157 811
rect 2053 706 2082 752
rect 2128 706 2157 752
rect 2053 647 2157 706
rect 2053 601 2082 647
rect 2128 601 2157 647
rect 2053 541 2157 601
rect 2053 495 2082 541
rect 2128 495 2157 541
rect 2053 435 2157 495
rect 2053 389 2082 435
rect 2128 389 2157 435
rect 2053 329 2157 389
rect 2053 283 2082 329
rect 2128 283 2157 329
rect 2053 270 2157 283
rect 2297 857 2385 870
rect 2297 811 2326 857
rect 2372 811 2385 857
rect 2297 752 2385 811
rect 2297 706 2326 752
rect 2372 706 2385 752
rect 2297 647 2385 706
rect 2297 601 2326 647
rect 2372 601 2385 647
rect 2297 541 2385 601
rect 2297 495 2326 541
rect 2372 495 2385 541
rect 2297 435 2385 495
rect 2297 389 2326 435
rect 2372 389 2385 435
rect 2297 329 2385 389
rect 2297 283 2326 329
rect 2372 283 2385 329
rect 2297 270 2385 283
<< mvpdiff >>
rect 1825 2545 1913 2558
rect 1825 1989 1838 2545
rect 1884 1989 1913 2545
rect 1825 1932 1913 1989
rect 1825 1886 1838 1932
rect 1884 1886 1913 1932
rect 1825 1829 1913 1886
rect 1825 1783 1838 1829
rect 1884 1783 1913 1829
rect 1825 1726 1913 1783
rect 1825 1680 1838 1726
rect 1884 1680 1913 1726
rect 1825 1623 1913 1680
rect 1825 1577 1838 1623
rect 1884 1577 1913 1623
rect 1825 1520 1913 1577
rect 1825 1474 1838 1520
rect 1884 1474 1913 1520
rect 1825 1417 1913 1474
rect 1825 1371 1838 1417
rect 1884 1371 1913 1417
rect 1825 1358 1913 1371
rect 2053 2545 2157 2558
rect 2053 1989 2082 2545
rect 2128 1989 2157 2545
rect 2053 1932 2157 1989
rect 2053 1886 2082 1932
rect 2128 1886 2157 1932
rect 2053 1829 2157 1886
rect 2053 1783 2082 1829
rect 2128 1783 2157 1829
rect 2053 1726 2157 1783
rect 2053 1680 2082 1726
rect 2128 1680 2157 1726
rect 2053 1623 2157 1680
rect 2053 1577 2082 1623
rect 2128 1577 2157 1623
rect 2053 1520 2157 1577
rect 2053 1474 2082 1520
rect 2128 1474 2157 1520
rect 2053 1417 2157 1474
rect 2053 1371 2082 1417
rect 2128 1371 2157 1417
rect 2053 1358 2157 1371
rect 2297 2545 2385 2558
rect 2297 1989 2326 2545
rect 2372 1989 2385 2545
rect 2297 1932 2385 1989
rect 2297 1886 2326 1932
rect 2372 1886 2385 1932
rect 2297 1829 2385 1886
rect 2297 1783 2326 1829
rect 2372 1783 2385 1829
rect 2297 1726 2385 1783
rect 2297 1680 2326 1726
rect 2372 1680 2385 1726
rect 2297 1623 2385 1680
rect 2297 1577 2326 1623
rect 2372 1577 2385 1623
rect 2297 1520 2385 1577
rect 2297 1474 2326 1520
rect 2372 1474 2385 1520
rect 2297 1417 2385 1474
rect 2297 1371 2326 1417
rect 2372 1371 2385 1417
rect 2297 1358 2385 1371
<< mvndiffc >>
rect 1838 811 1884 857
rect 1838 706 1884 752
rect 1838 601 1884 647
rect 1838 495 1884 541
rect 1838 389 1884 435
rect 1838 283 1884 329
rect 2082 811 2128 857
rect 2082 706 2128 752
rect 2082 601 2128 647
rect 2082 495 2128 541
rect 2082 389 2128 435
rect 2082 283 2128 329
rect 2326 811 2372 857
rect 2326 706 2372 752
rect 2326 601 2372 647
rect 2326 495 2372 541
rect 2326 389 2372 435
rect 2326 283 2372 329
<< mvpdiffc >>
rect 1838 1989 1884 2545
rect 1838 1886 1884 1932
rect 1838 1783 1884 1829
rect 1838 1680 1884 1726
rect 1838 1577 1884 1623
rect 1838 1474 1884 1520
rect 1838 1371 1884 1417
rect 2082 1989 2128 2545
rect 2082 1886 2128 1932
rect 2082 1783 2128 1829
rect 2082 1680 2128 1726
rect 2082 1577 2128 1623
rect 2082 1474 2128 1520
rect 2082 1371 2128 1417
rect 2326 1989 2372 2545
rect 2326 1886 2372 1932
rect 2326 1783 2372 1829
rect 2326 1680 2372 1726
rect 2326 1577 2372 1623
rect 2326 1474 2372 1520
rect 2326 1371 2372 1417
<< psubdiff >>
rect 1468 914 1558 936
rect 1468 22 1490 914
rect 1536 90 1558 914
rect 2528 1008 2618 1030
rect 2528 90 2550 1008
rect 1536 68 2550 90
rect 1536 22 1644 68
rect 2442 22 2550 68
rect 2596 22 2618 1008
rect 1468 0 2618 22
<< nsubdiff >>
rect 1468 2806 2618 2828
rect 1468 1350 1490 2806
rect 1536 2760 1644 2806
rect 2442 2760 2550 2806
rect 1536 2738 2550 2760
rect 1536 1350 1558 2738
rect 1468 1328 1558 1350
rect 2528 1350 2550 2738
rect 2596 1350 2618 2806
rect 2528 1328 2618 1350
<< psubdiffcont >>
rect 1490 22 1536 914
rect 1644 22 2442 68
rect 2550 22 2596 1008
<< nsubdiffcont >>
rect 1490 1350 1536 2806
rect 1644 2760 2442 2806
rect 2550 1350 2596 2806
<< polysilicon >>
rect 1913 2558 2053 2602
rect 2157 2558 2297 2602
rect 1913 1283 2053 1358
rect 1697 1248 2053 1283
rect 1697 1108 1716 1248
rect 1762 1108 2053 1248
rect 1697 1072 2053 1108
rect 1913 870 2053 1072
rect 2157 1248 2297 1358
rect 2157 1108 2196 1248
rect 2242 1108 2297 1248
rect 2157 870 2297 1108
rect 1913 226 2053 270
rect 2157 226 2297 270
<< polycontact >>
rect 1716 1108 1762 1248
rect 2196 1108 2242 1248
<< metal1 >>
rect 1479 2806 2607 2817
rect 1479 1350 1490 2806
rect 1536 2760 1644 2806
rect 2442 2760 2550 2806
rect 1536 2749 2550 2760
rect 1536 1350 1547 2749
rect 1479 1339 1547 1350
rect 1823 2545 1899 2558
rect 1823 1989 1838 2545
rect 1884 1989 1899 2545
rect 1823 1932 1899 1989
rect 1823 1886 1838 1932
rect 1884 1886 1899 1932
rect 1823 1829 1899 1886
rect 1823 1783 1838 1829
rect 1884 1783 1899 1829
rect 1823 1726 1899 1783
rect 1823 1680 1838 1726
rect 1884 1680 1899 1726
rect 1823 1623 1899 1680
rect 1823 1577 1838 1623
rect 1884 1577 1899 1623
rect 1823 1520 1899 1577
rect 1823 1474 1838 1520
rect 1884 1474 1899 1520
rect 1823 1417 1899 1474
rect 1823 1371 1838 1417
rect 1884 1371 1899 1417
rect 1823 1267 1899 1371
rect 2067 2545 2143 2749
rect 2067 1989 2082 2545
rect 2128 1989 2143 2545
rect 2067 1932 2143 1989
rect 2067 1886 2082 1932
rect 2128 1886 2143 1932
rect 2067 1829 2143 1886
rect 2067 1783 2082 1829
rect 2128 1783 2143 1829
rect 2067 1726 2143 1783
rect 2067 1680 2082 1726
rect 2128 1680 2143 1726
rect 2067 1623 2143 1680
rect 2067 1577 2082 1623
rect 2128 1577 2143 1623
rect 2067 1520 2143 1577
rect 2067 1474 2082 1520
rect 2128 1474 2143 1520
rect 2067 1417 2143 1474
rect 2067 1371 2082 1417
rect 2128 1371 2143 1417
rect 2067 1358 2143 1371
rect 2311 2545 2387 2558
rect 2311 1989 2326 2545
rect 2372 1989 2387 2545
rect 2311 1932 2387 1989
rect 2311 1886 2326 1932
rect 2372 1886 2387 1932
rect 2311 1829 2387 1886
rect 2311 1783 2326 1829
rect 2372 1783 2387 1829
rect 2311 1726 2387 1783
rect 2311 1680 2326 1726
rect 2372 1680 2387 1726
rect 2311 1623 2387 1680
rect 2311 1577 2326 1623
rect 2372 1577 2387 1623
rect 2311 1520 2387 1577
rect 2311 1474 2326 1520
rect 2372 1474 2387 1520
rect 2311 1417 2387 1474
rect 2311 1371 2326 1417
rect 2372 1371 2387 1417
rect 1140 1248 1773 1267
rect 1140 1108 1716 1248
rect 1762 1108 1773 1248
rect 1140 1089 1773 1108
rect 1823 1248 2261 1267
rect 1823 1108 2196 1248
rect 2242 1108 2261 1248
rect 1823 1089 2261 1108
rect 1479 914 1547 925
rect 1479 22 1490 914
rect 1536 79 1547 914
rect 1823 857 1899 1089
rect 1823 811 1838 857
rect 1884 811 1899 857
rect 1823 752 1899 811
rect 1823 706 1838 752
rect 1884 706 1899 752
rect 1823 647 1899 706
rect 1823 601 1838 647
rect 1884 601 1899 647
rect 1823 541 1899 601
rect 1823 495 1838 541
rect 1884 495 1899 541
rect 1823 435 1899 495
rect 1823 389 1838 435
rect 1884 389 1899 435
rect 1823 329 1899 389
rect 1823 283 1838 329
rect 1884 283 1899 329
rect 1823 270 1899 283
rect 2067 857 2143 870
rect 2067 811 2082 857
rect 2128 811 2143 857
rect 2067 752 2143 811
rect 2067 706 2082 752
rect 2128 706 2143 752
rect 2067 647 2143 706
rect 2067 601 2082 647
rect 2128 601 2143 647
rect 2067 541 2143 601
rect 2067 495 2082 541
rect 2128 495 2143 541
rect 2067 435 2143 495
rect 2067 389 2082 435
rect 2128 389 2143 435
rect 2067 329 2143 389
rect 2067 283 2082 329
rect 2128 283 2143 329
rect 2067 79 2143 283
rect 2311 857 2387 1371
rect 2539 1350 2550 2749
rect 2596 1350 2607 2806
rect 2539 1339 2607 1350
rect 2311 811 2326 857
rect 2372 811 2387 857
rect 2311 752 2387 811
rect 2311 706 2326 752
rect 2372 706 2387 752
rect 2311 647 2387 706
rect 2311 601 2326 647
rect 2372 601 2387 647
rect 2311 541 2387 601
rect 2311 495 2326 541
rect 2372 495 2387 541
rect 2311 435 2387 495
rect 2311 389 2326 435
rect 2372 389 2387 435
rect 2311 329 2387 389
rect 2311 283 2326 329
rect 2372 283 2387 329
rect 2311 270 2387 283
rect 2539 1008 2607 1019
rect 2539 79 2550 1008
rect 1536 68 2550 79
rect 1536 22 1644 68
rect 2442 22 2550 68
rect 2596 22 2607 1008
rect 1479 11 2607 22
use lvlshift_up  lvlshift_up_0
timestamp 1764347740
transform 1 0 -17795 0 1 -53410
box 18130 53410 19237 55988
<< labels >>
rlabel metal1 s 2349 1100 2349 1100 4 AB
port 2 nsew
rlabel metal1 s 2245 45 2245 45 4 DVSS
port 4 nsew
rlabel metal1 s 2254 2788 2254 2788 4 DVDD
port 5 nsew
<< end >>
