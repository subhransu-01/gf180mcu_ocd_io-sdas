magic
tech gf180mcuD
magscale 1 10
timestamp 1764281188
<< polysilicon >>
rect 794 8377 972 8396
rect 794 8331 813 8377
rect 953 8331 972 8377
rect 794 8312 972 8331
rect 2598 8377 2776 8396
rect 2598 8331 2617 8377
rect 2757 8331 2776 8377
rect 2598 8312 2776 8331
rect 3002 8377 3180 8396
rect 3002 8331 3021 8377
rect 3161 8331 3180 8377
rect 3002 8312 3180 8331
rect 4806 8377 4984 8396
rect 4806 8331 4825 8377
rect 4965 8331 4984 8377
rect 4806 8312 4984 8331
rect 5210 8377 5388 8396
rect 5210 8331 5229 8377
rect 5369 8331 5388 8377
rect 5210 8312 5388 8331
rect 7014 8377 7192 8396
rect 7014 8331 7033 8377
rect 7173 8331 7192 8377
rect 7014 8312 7192 8331
rect 7418 8377 7596 8396
rect 7418 8331 7437 8377
rect 7577 8331 7596 8377
rect 7418 8312 7596 8331
rect 9222 8377 9400 8396
rect 9222 8331 9241 8377
rect 9381 8331 9400 8377
rect 9222 8312 9400 8331
rect 803 8300 963 8312
rect 2607 8300 2767 8312
rect 3011 8300 3171 8312
rect 4815 8300 4975 8312
rect 5219 8300 5379 8312
rect 7023 8300 7183 8312
rect 7427 8300 7587 8312
rect 9231 8300 9391 8312
rect 794 703 972 722
rect 794 657 813 703
rect 953 657 972 703
rect 794 638 972 657
rect 2598 703 2776 722
rect 2598 657 2617 703
rect 2757 657 2776 703
rect 2598 638 2776 657
rect 3002 703 3180 722
rect 3002 657 3021 703
rect 3161 657 3180 703
rect 3002 638 3180 657
rect 4806 703 4984 722
rect 4806 657 4825 703
rect 4965 657 4984 703
rect 4806 638 4984 657
rect 5211 703 5389 722
rect 5211 657 5230 703
rect 5370 657 5389 703
rect 5211 638 5389 657
rect 7014 703 7192 722
rect 7014 657 7033 703
rect 7173 657 7192 703
rect 7014 638 7192 657
rect 7417 703 7595 722
rect 7417 657 7436 703
rect 7576 657 7595 703
rect 7417 638 7595 657
rect 9222 703 9400 722
rect 9222 657 9241 703
rect 9381 657 9400 703
rect 9222 638 9400 657
<< polycontact >>
rect 813 8331 953 8377
rect 2617 8331 2757 8377
rect 3021 8331 3161 8377
rect 4825 8331 4965 8377
rect 5229 8331 5369 8377
rect 7033 8331 7173 8377
rect 7437 8331 7577 8377
rect 9241 8331 9381 8377
rect 813 657 953 703
rect 2617 657 2757 703
rect 3021 657 3161 703
rect 4825 657 4965 703
rect 5230 657 5370 703
rect 7033 657 7173 703
rect 7436 657 7576 703
rect 9241 657 9381 703
<< metal1 >>
rect -251 9400 4976 9508
rect -251 9240 3172 9340
rect -251 9080 2768 9180
rect -251 8920 964 9020
rect 802 8377 964 8920
rect 802 8331 813 8377
rect 953 8331 964 8377
rect 802 8320 964 8331
rect 2606 8377 2768 9080
rect 2606 8331 2617 8377
rect 2757 8331 2768 8377
rect 2606 8320 2768 8331
rect 3010 8377 3172 9240
rect 3010 8331 3021 8377
rect 3161 8331 3172 8377
rect 3010 8320 3172 8331
rect 4814 8377 4976 9400
rect 4814 8331 4825 8377
rect 4965 8331 4976 8377
rect 4814 8320 4976 8331
rect 5218 9400 10510 9508
rect 5218 8377 5380 9400
rect 5218 8331 5229 8377
rect 5369 8331 5380 8377
rect 5218 8320 5380 8331
rect 7022 9240 10510 9340
rect 7022 8377 7184 9240
rect 7022 8331 7033 8377
rect 7173 8331 7184 8377
rect 7022 8320 7184 8331
rect 7426 9080 10510 9180
rect 7426 8377 7588 9080
rect 7426 8331 7437 8377
rect 7577 8331 7588 8377
rect 7426 8320 7588 8331
rect 9230 8920 10510 9020
rect 9230 8377 9392 8920
rect 9230 8331 9241 8377
rect 9381 8331 9392 8377
rect 9230 8320 9392 8331
rect 302 363 559 8212
rect 849 714 895 8320
rect 2675 714 2721 8320
rect 3057 714 3103 8320
rect 4883 714 4929 8320
rect 5265 714 5311 8320
rect 7091 714 7137 8320
rect 7473 714 7519 8320
rect 9299 714 9345 8320
rect 9391 812 9967 8212
rect 802 703 964 714
rect 802 657 813 703
rect 953 657 964 703
rect 802 646 964 657
rect 2606 703 2768 714
rect 2606 657 2617 703
rect 2757 657 2768 703
rect 2606 646 2768 657
rect 3010 703 3172 714
rect 3010 657 3021 703
rect 3161 657 3172 703
rect 3010 646 3172 657
rect 4814 703 4976 714
rect 4814 657 4825 703
rect 4965 657 4976 703
rect 4814 646 4976 657
rect 5219 703 5381 714
rect 5219 657 5230 703
rect 5370 657 5381 703
rect 5219 646 5381 657
rect 7022 703 7184 714
rect 7022 657 7033 703
rect 7173 657 7184 703
rect 7022 646 7184 657
rect 7425 703 7587 714
rect 7425 657 7436 703
rect 7576 657 7587 703
rect 7425 646 7587 657
rect 9230 703 9392 714
rect 9230 657 9241 703
rect 9381 657 9392 703
rect 9230 646 9392 657
rect 9730 363 9967 812
use comp018green_out_drv_nleg_6T  comp018green_out_drv_nleg_6T_0
timestamp 1764281188
transform 1 0 7221 0 1 680
box 48 42 2328 7632
use comp018green_out_drv_nleg_6T  comp018green_out_drv_nleg_6T_1
timestamp 1764281188
transform 1 0 5013 0 1 680
box 48 42 2328 7632
use comp018green_out_drv_nleg_6T  comp018green_out_drv_nleg_6T_2
timestamp 1764281188
transform 1 0 2805 0 1 680
box 48 42 2328 7632
use comp018green_out_drv_nleg_6T  comp018green_out_drv_nleg_6T_3
timestamp 1764281188
transform 1 0 597 0 1 680
box 48 42 2328 7632
use GR_NMOS  GR_NMOS_0
timestamp 1764270562
transform 1 0 363 0 1 436
box -1789 -834 11222 10481
use nmos_metal_stack  nmos_metal_stack_0
timestamp 1758724778
transform -1 0 9591 0 1 812
box -44 0 2004 7400
use nmos_metal_stack  nmos_metal_stack_1
timestamp 1758724778
transform 1 0 7227 0 1 812
box -44 0 2004 7400
use nmos_metal_stack  nmos_metal_stack_2
timestamp 1758724778
transform 1 0 5019 0 1 812
box -44 0 2004 7400
use nmos_metal_stack  nmos_metal_stack_3
timestamp 1758724778
transform 1 0 2811 0 1 812
box -44 0 2004 7400
use nmos_metal_stack  nmos_metal_stack_4
timestamp 1758724778
transform 1 0 603 0 1 812
box -44 0 2004 7400
<< end >>
