** sch_path: /home/subhransu/gitRepo/gf180mcu_ocd_io-sdas/runs/RUN_2026-01-13_06-45-48/parameters/dc_response/run_1/io_inv_1_dc.sch
**.subckt io_inv_1_dc
x1 Vin Vout VDD VSS io_inv_1
V1 VSS GND 0
V2 VDD GND 1.8
V3 Vin GND 1.8
C1 Vout GND 1e-15 m=1
**** begin user architecture code





*.include {PDK_ROOT}/{PDK}/libs.tech/ngspice/design.ngspice
*.lib {PDK_ROOT}/{PDK}/libs.tech/ngspice/sm141064.ngspice {corner}
.include /home/subhransu/gitRepo/gf180mcu_ocd_io-sdas/netlist/schematic/io_inv_1.spice
.temp 27
.option SEED=12345
.option warn=1





.control
dc V3 0 1.8 0.01
set wr_singlescale
wrdata /home/subhransu/gitRepo/gf180mcu_ocd_io-sdas/runs/RUN_2026-01-13_06-45-48/parameters/dc_response/run_1/io_inv_1_dc_1.data V(Vin) V(Vout)
.endc



.include /home/subhransu/share/pdk/gf180mcuD/libs.tech/ngspice/design.ngspice
.lib /home/subhransu/share/pdk/gf180mcuD/libs.tech/ngspice/sm141064.ngspice tt

**** end user architecture code
**.ends
.GLOBAL GND
.end
