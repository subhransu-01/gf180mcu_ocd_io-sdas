VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO gf180mcu_ocd_io__bi_a
  CLASS PAD INOUT ;
  FOREIGN gf180mcu_ocd_io__bi_a ;
  ORIGIN 0.000 0.000 ;
  SIZE 75.000 BY 350.000 ;
  SYMMETRY X Y R90 ;
  SITE GF_IO_Site ;
  PIN A
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.504000 ;
    ANTENNADIFFAREA 1.000000 ;
    PORT
      LAYER Metal2 ;
        RECT 69.400 267.070 69.780 350.000 ;
    END
  END A
  PIN ANA
    ANTENNAGATEAREA 21.490000 ;
    ANTENNADIFFAREA 80.000000 ;
    PORT
      LAYER Metal2 ;
        RECT 8.530 321.790 8.910 350.005 ;
    END
  END ANA
  PIN CS
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.504000 ;
    ANTENNADIFFAREA 1.000000 ;
    PORT
      LAYER Metal2 ;
        RECT 3.360 328.545 3.740 350.000 ;
    END
  END CS
  PIN DVDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 182.000 8.810 197.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0.000 214.000 5.000 229.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0.000 334.000 5.000 341.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0.000 294.000 17.930 301.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0.000 278.000 17.930 285.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0.000 270.000 17.930 277.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0.000 262.000 9.070 269.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0.000 206.000 9.815 213.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0.000 118.000 5.000 125.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0.000 134.000 8.810 149.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0.000 150.000 8.905 165.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0.000 166.000 8.905 181.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 70.000 182.000 75.000 197.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 70.000 214.000 75.000 229.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 70.000 334.000 75.000 341.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 70.000 294.000 75.000 301.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 49.445 278.000 75.000 285.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 67.195 270.000 75.000 277.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 70.000 262.000 75.000 269.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 70.000 206.000 75.000 213.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 70.000 118.000 75.000 125.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 70.000 134.000 75.000 149.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 70.000 150.000 75.000 165.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 70.000 166.000 75.000 181.000 ;
    END
  END DVDD
  PIN DVSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 86.000 5.000 101.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0.000 70.000 5.000 85.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0.000 230.000 5.000 245.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0.000 198.000 5.000 205.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0.000 102.000 5.000 117.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0.000 126.000 5.000 133.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0.000 286.000 22.880 293.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0.000 302.000 25.555 309.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0.000 326.000 9.320 333.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0.000 342.000 9.320 348.390 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 62.215 86.000 75.000 101.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 62.215 70.000 75.000 85.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 59.650 230.000 75.000 245.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 66.125 198.000 75.000 205.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 62.215 102.000 75.000 117.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 70.000 126.000 75.000 133.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 55.255 286.000 75.000 293.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 54.080 302.000 75.000 309.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 63.580 326.000 75.000 333.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 68.000 342.000 75.000 348.390 ;
    END
  END DVSS
  PIN IE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.504000 ;
    ANTENNADIFFAREA 1.000000 ;
    PORT
      LAYER Metal2 ;
        RECT 11.385 334.920 11.765 350.000 ;
    END
  END IE
  PIN OE
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 2.016000 ;
    ANTENNADIFFAREA 7.776000 ;
    PORT
      LAYER Metal2 ;
        RECT 70.130 283.445 70.510 350.000 ;
    END
  END OE
  PIN PAD
    DIRECTION INOUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 258.720001 ;
    PORT
      LAYER Metal3 ;
        RECT 7.500 2.000 67.500 62.000 ;
    END
  END PAD
  PIN PD
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.512000 ;
    ANTENNADIFFAREA 1.000000 ;
    PORT
      LAYER Metal2 ;
        RECT 10.330 330.100 10.710 350.000 ;
    END
  END PD
  PIN PDRV0
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.504000 ;
    ANTENNADIFFAREA 2.592000 ;
    PORT
      LAYER Metal2 ;
        RECT 7.110 326.870 7.490 350.000 ;
    END
  END PDRV0
  PIN PDRV1
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.504000 ;
    ANTENNADIFFAREA 2.592000 ;
    PORT
      LAYER Metal2 ;
        RECT 7.820 326.280 8.200 350.005 ;
    END
  END PDRV1
  PIN PU
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 1.008000 ;
    ANTENNADIFFAREA 1.795000 ;
    PORT
      LAYER Metal2 ;
        RECT 5.965 330.420 6.345 350.000 ;
    END
  END PU
  PIN SL
    DIRECTION INPUT ;
    USE SIGNAL ;
    ANTENNAGATEAREA 0.504000 ;
    ANTENNADIFFAREA 1.000000 ;
    PORT
      LAYER Metal2 ;
        RECT 68.670 266.340 69.050 350.000 ;
    END
  END SL
  PIN VDD
    DIRECTION INOUT ;
    USE POWER ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 254.000 5.000 261.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0.000 310.000 5.000 317.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 67.385 254.000 75.000 261.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 70.000 310.000 75.000 317.000 ;
    END
  END VDD
  PIN VSS
    DIRECTION INOUT ;
    USE GROUND ;
    PORT
      LAYER Metal3 ;
        RECT 0.000 318.000 5.000 325.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 0.000 246.000 5.000 253.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 70.000 318.000 75.000 325.000 ;
    END
    PORT
      LAYER Metal3 ;
        RECT 70.000 246.000 75.000 253.000 ;
    END
  END VSS
  PIN Y
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    ANTENNADIFFAREA 3.240000 ;
    PORT
      LAYER Metal2 ;
        RECT 70.860 319.900 71.240 350.000 ;
    END
  END Y
  OBS
      LAYER Nwell ;
        RECT 1.820 68.895 73.180 346.535 ;
      LAYER Metal1 ;
        RECT -0.160 65.540 75.160 349.785 ;
      LAYER Metal2 ;
        RECT 0.000 328.245 3.060 348.375 ;
        RECT 4.040 330.120 5.665 348.375 ;
        RECT 6.645 330.120 6.810 348.375 ;
        RECT 4.040 328.245 6.810 330.120 ;
        RECT 0.000 326.570 6.810 328.245 ;
        RECT 9.210 329.800 10.030 348.375 ;
        RECT 11.010 334.620 11.085 348.375 ;
        RECT 12.065 334.620 68.370 348.375 ;
        RECT 11.010 329.800 68.370 334.620 ;
        RECT 0.000 325.980 7.520 326.570 ;
        RECT 0.000 321.490 8.230 325.980 ;
        RECT 9.210 321.490 68.370 329.800 ;
        RECT 0.000 266.040 68.370 321.490 ;
        RECT 71.540 319.600 75.000 348.375 ;
        RECT 70.810 283.145 75.000 319.600 ;
        RECT 70.080 266.770 75.000 283.145 ;
        RECT 69.350 266.040 75.000 266.770 ;
        RECT 0.000 0.000 75.000 266.040 ;
      LAYER Metal3 ;
        RECT 11.120 340.200 66.200 348.390 ;
        RECT 6.800 334.800 68.200 340.200 ;
        RECT 11.120 324.200 61.780 334.800 ;
        RECT 6.800 310.800 68.200 324.200 ;
        RECT 27.355 300.200 52.280 310.800 ;
        RECT 19.730 294.800 68.200 300.200 ;
        RECT 24.680 286.800 53.455 294.800 ;
        RECT 24.680 284.200 47.645 286.800 ;
        RECT 19.730 276.200 47.645 284.200 ;
        RECT 19.730 268.200 65.395 276.200 ;
        RECT 10.870 262.800 68.200 268.200 ;
        RECT 10.870 260.200 65.585 262.800 ;
        RECT 6.800 252.200 65.585 260.200 ;
        RECT 6.800 246.800 68.200 252.200 ;
        RECT 6.800 228.200 57.850 246.800 ;
        RECT 6.800 214.800 68.200 228.200 ;
        RECT 11.615 206.800 68.200 214.800 ;
        RECT 11.615 204.200 64.325 206.800 ;
        RECT 6.800 198.800 64.325 204.200 ;
        RECT 10.610 196.200 64.325 198.800 ;
        RECT 10.610 182.800 68.200 196.200 ;
        RECT 10.705 148.200 68.200 182.800 ;
        RECT 10.610 132.200 68.200 148.200 ;
        RECT 6.800 118.800 68.200 132.200 ;
        RECT 6.800 68.200 60.415 118.800 ;
        RECT 0.665 63.800 73.640 68.200 ;
        RECT 0.665 0.200 5.700 63.800 ;
        RECT 69.300 0.200 73.640 63.800 ;
        RECT 0.665 0.000 73.640 0.200 ;
  END
END gf180mcu_ocd_io__bi_a
END LIBRARY

