magic
tech gf180mcuD
magscale 1 10
timestamp 1764277317
<< error_s >>
rect 29440 44570 32000 44578
rect 27739 44542 29055 44550
rect 29564 44446 32000 44454
rect 27741 44418 29057 44426
rect 29688 44322 32000 44330
rect 27731 44294 29171 44302
rect 29812 44198 32000 44206
rect 27762 44170 29326 44178
rect 29936 44074 32000 44082
rect 27752 44046 29440 44054
rect 30060 43950 32000 43958
rect 27833 43922 29577 43930
rect 30184 43826 32000 43834
rect 27957 43798 29701 43806
use comp018green_esd_clamp_v5p0_1  comp018green_esd_clamp_v5p0_1_0
timestamp 1764277317
transform 1 0 43564 0 1 51
box -4188 -51 13013 56967
use comp018green_esd_clamp_v5p0_2  comp018green_esd_clamp_v5p0_2_0
timestamp 1764277317
transform 0 1 51 1 0 43565
box -407 -51 13369 47415
use power_via_cor_3  power_via_cor_3_0
timestamp 1758726819
transform 1 0 42556 0 1 508
box 1094 35210 14833 56443
use power_via_cor_5  power_via_cor_5_0
timestamp 1758726819
transform 0 1 508 1 0 42557
box 1068 32 14833 50982
<< end >>
